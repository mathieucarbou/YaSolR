PK
     mdZ��9�h �h    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":[],"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":[],"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"],"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"],"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4":["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5":["pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"],"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6":["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7":["pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"],"pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10"],"pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_4":[],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6":["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7":["pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8":["pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9":["pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1"],"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10":["pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0"],"pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8"],"pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7"],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":[],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6"],"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":[],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6"],"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"],"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"],"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4"],"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5":["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0"],"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7":["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"],"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6":["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1":["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3":["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6":["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],"pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0":["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"],"pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1":["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7"],"pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5"],"pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]},"pin_to_color":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"#005F39","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"#9E008E","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"#FF6E41","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"#00FFC6","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"#774D00","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"#FFA6FE","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"#005F39","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"#9E008E","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"#B500FF","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"#FFB167","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"#001544","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"#91D0CB","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"#007DB5","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"#000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"#000000","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0":"#005F39","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1":"#FFB167","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2":"#B500FF","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3":"#9E008E","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4":"#FF6E41","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5":"#C28C9F","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6":"#00FFC6","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7":"#008F9C","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0":"#FFDB66","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1":"#90FB92","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0":"#9E008E","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1":"#005F39","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2":"#774D00","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3":"#FFA6FE","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_4":"#000000","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5":"#FF6E41","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6":"#00FFC6","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7":"#95003A","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8":"#FF937E","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9":"#90FB92","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10":"#FFDB66","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0":"#FF937E","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1":"#95003A","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"#000000","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"#FFE502","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"#E85EBE","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"#000000","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"#005F39","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"#010067","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"#0076FF","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"#85A900","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0":"#005F39","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1":"#FFB167","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2":"#B500FF","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3":"#9E008E","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4":"#FF6E41","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5":"#6A826C","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6":"#00FFC6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7":"#00AE7E","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"#0076FF","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"#85A900","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"#9E008E","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"#E85EBE","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"#0076FF","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"#85A900","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"#0E4CA1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"#010067","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0":"#005F39","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1":"#9E008E","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2":"#007DB5","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3":"#001544","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4":"#0E4CA1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5":"#010067","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6":"#005F39","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0":"#005F39","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1":"#9E008E","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2":"#007DB5","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3":"#91D0CB","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4":"#9E008E","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5":"#E85EBE","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6":"#FFE502","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0":"#6A826C","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1":"#00AE7E","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0":"#C28C9F","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1":"#008F9C","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"#0076FF","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"#85A900","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"#00FFC6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"#FF6E41"},"pin_to_state":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"neutral","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"neutral","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"neutral","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0":"neutral","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1":"neutral","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2":"neutral","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3":"neutral","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4":"neutral","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5":"neutral","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6":"neutral","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7":"neutral","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0":"neutral","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_4":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9":"neutral","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10":"neutral","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0":"neutral","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"neutral","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"neutral","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"neutral","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"neutral","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"neutral","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0":"neutral","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1":"neutral","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2":"neutral","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3":"neutral","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4":"neutral","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5":"neutral","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6":"neutral","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"neutral","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"neutral","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5":"neutral","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5":"neutral","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6":"neutral","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0":"neutral","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1":"neutral","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0":"neutral","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"neutral","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"neutral"},"next_color_idx":14,"wires_placed_in_order":[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28"],["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"],["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"],["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"],["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"],["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"],["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5"],["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"],["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"],["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1"],["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"],["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1"],["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],["pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"],["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"],["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"],["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"],["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0"],["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0"],["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28"]]],[[],[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"]]],[[],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15"]]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29"]]],[[],[]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_15","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0"]],[]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1"],["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_28","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]]],[[["pin-type-component_7596dca9-ef35-4a25-9667-71a309c38942_29","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"]]],[[],[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"]]],[[],[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"]]],[[],[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"]]],[[],[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"]]],[[],[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0","pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5"]]],[[],[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"]]],[[],[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"]]],[[],[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1"]]],[[],[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[["pin-type-component_a8221eb9-381c-43f6-a63c-1fa17c525231_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"]]],[[],[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"]]],[[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36"]],[]],[[["pin-type-component_87584d7b-427c-4128-9f1d-c39754565c83_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2"]],[]],[[["pin-type-component_a710ae78-12af-4c40-8eab-c282b0818a9f_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15"]],[]],[[["pin-type-component_3de1381f-af91-4dcf-856b-586dd46839d7_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_0","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_0"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_1","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_2"]],[]],[[["pin-type-component_72c2b56f-df5d-4021-9811-2825ccb29077_2","pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_1"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_0","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_0"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_2","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_1"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_1","pin-type-component_28a290ea-5e4c-4306-af0e-9b019cace231_2"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_164aeb04-09d1-4d57-afc3-356f83e7dfc8_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_9fb701f6-bd34-49c7-aee5-a09df94bb16b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_0","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_0"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_1","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_2"]],[]],[[["pin-type-component_61d88a57-e2bc-4d7f-ad52-bfcec31c3d76_2","pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_1"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_6bdfaf63-c660-411b-b5de-7e67c510171d_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23"]],[]],[[["pin-type-component_cff1c91e-23de-4c4e-aa78-b4dc7a6518dd_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25"]],[]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]]],[[],[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1"]]],[[],[["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[],[["pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]]],[[],[["pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"]]],[[["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"],["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_9774de9e-22ea-4833-97c5-561329cd52b5_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"],["pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_0"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_f4c5cbef-1786-408a-ad96-c821116a8865_1"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"],["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_0"]],[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_4505265e-df0a-43f9-9110-8440d5f596f6_1"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]],[]],[[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3"]],[]],[[["pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]],[]],[[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"]]],[[],[["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"]]],[[],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1"]]],[[],[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"]]],[[],[["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"]]],[[],[["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32"]]],[[],[["pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0"]]],[[],[["pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0"]]],[[],[["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"]]],[[],[["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"]]],[[],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"]]],[[],[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]],[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_1a407f64-89bd-4888-9631-f96c6341551c_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3"],["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5"],["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]],[]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"]]],[[["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]],[]],[[],[["pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"]]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]],[]],[[["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]],[]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"]]],[[],[["pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0":"0000000000000000","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1":"0000000000000001","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2":"0000000000000011","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3":"0000000000000010","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_0":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_1":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_2":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_3":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_4":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_5":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_6":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_7":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_8":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_9":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10":"0000000000000003","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11":"0000000000000002","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_12":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_13":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_14":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_15":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_16":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_17":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_18":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19":"0000000000000000","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_20":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_21":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_22":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_23":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24":"0000000000000001","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_25":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26":"0000000000000006","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27":"0000000000000007","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28":"0000000000000020","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29":"0000000000000021","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_30":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_31":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32":"0000000000000022","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_33":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_34":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_35":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_36":"_","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_37":"_","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0":"0000000000000000","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1":"0000000000000007","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2":"0000000000000006","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3":"0000000000000001","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4":"0000000000000011","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5":"0000000000000025","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6":"0000000000000010","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7":"0000000000000026","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0":"0000000000000008","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1":"0000000000000009","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0":"0000000000000001","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1":"0000000000000000","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2":"0000000000000003","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3":"0000000000000002","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_4":"_","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5":"0000000000000011","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6":"0000000000000010","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7":"0000000000000018","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8":"0000000000000019","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9":"0000000000000009","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10":"0000000000000008","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0":"0000000000000019","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1":"0000000000000018","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_0":"_","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1":"0000000000000016","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2":"0000000000000012","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_0":"_","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1":"0000000000000017","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2":"0000000000000013","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0":"0000000000000004","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1":"0000000000000005","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0":"0000000000000000","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1":"0000000000000007","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2":"0000000000000006","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3":"0000000000000001","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4":"0000000000000011","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5":"0000000000000023","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6":"0000000000000010","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7":"0000000000000024","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0":"0000000000000004","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1":"0000000000000005","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2":"0000000000000014","pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3":"0000000000000012","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0":"0000000000000004","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1":"0000000000000005","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2":"0000000000000015","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3":"0000000000000013","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0":"0000000000000000","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1":"0000000000000001","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2":"0000000000000022","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3":"0000000000000020","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4":"0000000000000015","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5":"0000000000000013","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6":"0000000000000017","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0":"0000000000000000","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1":"0000000000000001","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2":"0000000000000022","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3":"0000000000000021","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4":"0000000000000014","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5":"0000000000000012","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6":"0000000000000016","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0":"0000000000000023","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1":"0000000000000024","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0":"0000000000000025","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1":"0000000000000026","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0":"0000000000000004","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1":"0000000000000005","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2":"0000000000000010","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3":"0000000000000011"},"component_id_to_pins":{"d53bc8d1-adbf-42c3-9bdc-27d4d2b68588":["0","1","2","3"],"f7d25e04-bb51-41df-ba72-c452c270d3fb":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31","32","33","34","35","36","37"],"32608709-bcb5-4c22-82f1-0b5ac1739be0":[],"915b317b-63a4-4c37-8362-9a35870cbe7c":[],"22500cd3-352c-4d79-9f9c-f48cf0a80685":["0","1","2","3","4","5","6","7"],"7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a":["0","1"],"ae19664f-1584-4f12-9c79-f0e8930ce70b":["0","1","2","3","4","5","6","7","8","9","10"],"1a4c0ab2-15d7-4f55-82c5-02526f5965a4":["0","1"],"b8cf9931-5e29-4c19-b0ce-f047cf1b7a61":[],"9e0cc72b-cce0-4555-8c60-9928baea3faa":[],"41689d80-6f1a-478b-ad5a-826ce578b4af":[],"ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8":["0","1","2"],"00e3d6c2-f801-4d91-ad4d-237bada773bb":["0","1","2"],"1c19cc90-e27a-4c31-a566-dce6d12cc7bd":["0","1"],"8b4859a0-119b-4d24-8c3e-f008f1af2f35":[],"eb1dbc1c-94ee-4954-b264-2ba5f2bb6c04":[],"99cae55d-e9c7-468a-acc3-dcac762056db":["0","1","2","3","4","5","6","7"],"e5530feb-ce19-40b3-8da6-a6ca8e4b619a":[],"060f78c2-f7c5-4b91-a54e-26722a6a6eb1":["0","1","2","3"],"c483e859-dbe3-40ab-ad85-fdb0e9726a1e":["0","1","2","3"],"d7e83964-79f2-4e6f-ab07-dee67fd9dff8":["0","1","2","3","4","5","6"],"6bde5401-8877-4618-b129-167654a129ea":["0","1","2","3","4","5","6"],"786922c4-3cc4-4e2e-a1af-6f582a726cc5":[],"c6b89f01-cd33-4f53-a410-bd8ce0a19726":[],"028c5ed6-a9ce-4916-bd5a-20a0af91ff53":[],"d8ee4efe-302f-41eb-a87d-4235620299ce":[],"8c415f8f-024b-42a7-9906-fa5d9103b190":[],"f0886e27-8ec0-43da-a659-1cbab4912d9c":[],"265be517-7dce-4507-b222-49efa0b79d44":[],"4d6635ca-f74e-4111-b736-96f73dea815d":[],"34d49454-fe1f-4693-a2f3-2121a541126c":[],"320ab8ff-f5d3-4096-b4aa-da43287dff93":["0","1"],"d008a2f8-2853-4c0d-8d67-a8220f145d26":["0","1"],"cabc8f6d-4e36-40d8-b46e-f81e3606417d":[],"0532153d-ec59-4dd7-ad03-6d0401cd55c5":[],"9b271475-bebe-41b8-aded-20e21ef4734b":["0","1","2","3"]},"uid_to_net":{"_":[],"0000000000000001":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1"],"0000000000000000":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0"],"0000000000000002":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11"],"0000000000000003":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10"],"0000000000000006":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2"],"0000000000000007":["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27","pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1"],"0000000000000008":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0"],"0000000000000009":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9","pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1"],"0000000000000004":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0"],"0000000000000005":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1","pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1","pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1"],"0000000000000010":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3"],"0000000000000011":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4","pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3","pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5","pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2"],"0000000000000012":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2"],"0000000000000013":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2"],"0000000000000014":["pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4"],"0000000000000015":["pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2","pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4"],"0000000000000016":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6","pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1"],"0000000000000017":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6","pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1"],"0000000000000018":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1"],"0000000000000019":["pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8","pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0"],"0000000000000020":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28"],"0000000000000021":["pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29"],"0000000000000022":["pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2","pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32","pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2"],"0000000000000023":["pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0","pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5"],"0000000000000024":["pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7","pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1"],"0000000000000025":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0"],"0000000000000026":["pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7","pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1"]},"uid_to_text_label":{"0000000000000001":"Net 1","0000000000000000":"Net 0","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000006":"Net 6","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000009":"Net 9","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16","0000000000000017":"Net 17","0000000000000018":"Net 18","0000000000000019":"Net 19","0000000000000020":"Net 20","0000000000000021":"Net 21","0000000000000022":"Net 22","0000000000000023":"Net 23","0000000000000024":"Net 24","0000000000000025":"Net 25","0000000000000026":"Net 26"},"all_breadboard_info_list":[],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[202.3552975,529.8953134999997],"typeId":"c2a09f2b-df40-42a6-8e0c-c519ba38e9d5","componentVersion":1,"instanceId":"d53bc8d1-adbf-42c3-9bdc-27d4d2b68588","orientation":"up","circleData":[[197.5,395],[213.0759055000001,396.3743885],[213.99214600000005,649.2539554999994],[200.70681100000002,650.6282869999995]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"GND","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[259.59212209496786,426.2251000087314],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"32608709-bcb5-4c22-82f1-0b5ac1739be0","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"VCC +5V","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[126.11683130463507,423.8059167969202],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"915b317b-63a4-4c37-8362-9a35870cbe7c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-165.78929000000034,-252.08162800000107],"typeId":"25d95763-f48b-4a99-bdb2-8bb3b7ccff88","componentVersion":1,"instanceId":"22500cd3-352c-4d79-9f9c-f48cf0a80685","orientation":"down","circleData":[[-12.500000000000426,-235.00000000000085],[-12.500000000000426,-250.00000000000085],[-12.500000000000426,-265.000000000001],[-12.500000000000426,-280.0000000000008],[-350.00000000000017,-235.00000000000085],[-350.00000000000017,-265.000000000001],[-350.00000000000017,-212.50000000000074],[-350.00000000000017,-295.00000000000114]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3397.3552479999994,1286.995553000001],"typeId":"2ce95dbd-bb8b-430f-8511-f580783f914c","componentVersion":1,"instanceId":"7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a","orientation":"left","circleData":[[3407.5,1190],[3422.5,1182.5]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[2142.5005030000007,435.00049550000006],"typeId":"840a331c-2aef-4dd8-892c-7ae81d6bcea5","componentVersion":2,"instanceId":"ae19664f-1584-4f12-9c79-f0e8930ce70b","orientation":"up","circleData":[[1967.5,395],[1967.9580910000004,425],[1967.5,455],[1967.5,492.50000000000006],[2110,567.5],[2305.000000000001,410],[2305.000000000001,462.49999999999983],[2054.1325,309.50149999999974],[2079.5350000000003,308.6104999999998],[2206.8475000000008,310.3924999999998],[2230.6180000000004,310.8394999999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[2214.4955529999997,2010.1447519999992],"typeId":"2ce95dbd-bb8b-430f-8511-f580783f914c","componentVersion":1,"instanceId":"1a4c0ab2-15d7-4f55-82c5-02526f5965a4","orientation":"down","circleData":[[2117.5,2000],[2110,1984.9999999999995]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[816.5526985000006,-114.18805750000007],"typeId":"b975acdd-73e3-4b18-a5a5-9b66f369afa0","componentVersion":2,"instanceId":"f7d25e04-bb51-41df-ba72-c452c270d3fb","orientation":"up","circleData":[[947.5,-340.00000000000006],[948.1030000000001,-312.73920549999985],[948.1231135000003,-286.7030244999998],[947.5,-258.2146149999999],[948.7261135000003,-232.17843399999987],[947.5,-206.1221394999999],[948.7261135000003,-178.25684499999983],[948.7261135000003,-152.22066399999994],[948.7261135000003,-124.95986949999983],[948.1030000000001,-99.55068849999985],[949.3291135000004,-71.68539399999995],[949.3291135000004,-44.42309949999995],[949.3291135000004,-16.561691499999938],[949.9306135000002,9.472989500000153],[949.3291135000004,35.48905700000002],[950.5552270000003,64.60058],[949.9306135000002,90.63676099999971],[949.9306135000002,118.52216899999956],[951.7813405000002,146.98896349999978],[678.5382805000002,148.19346349999984],[677.312167,120.32966899999968],[678.5382805000002,94.29348799999975],[677.9352805000001,66.42969349999983],[677.9352805000001,39.16739899999983],[679.1613940000002,12.528216500000212],[678.5382805000002,-14.131078000000002],[679.1613940000002,-43.24259950000001],[677.9352805000001,-70.48328049999995],[677.9352805000001,-95.9164614999999],[677.3322805000003,-121.95264249999988],[677.3322805000003,-149.81793699999986],[677.312167,-176.45323149999984],[678.5583940000001,-203.71402599999982],[677.3322805000003,-229.73009349999984],[675.4824745000001,-258.842026],[677.3322805000003,-284.294911],[677.9349745000002,-310.9130259999999],[677.3322805000003,-338.77388650000006]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 1 AC Circuit\n(behind a breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2521.1223679499117,1492.667604045154],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"9e0cc72b-cce0-4555-8c60-9928baea3faa","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 2 AC Circuit\n(behind a breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2767.5835720784066,1691.9991453659359],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"41689d80-6f1a-478b-ad5a-826ce578b4af","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"AC Circuit for components\n(behind 2A breaker)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3037.3754870576977,1907.3736162088799],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"b8cf9931-5e29-4c19-b0ce-f047cf1b7a61","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[544.7008329999994,1699.1917940000021],"typeId":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"instanceId":"ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8","orientation":"up","circleData":[[4067.500000000001,3905],[812.4999999999995,1715.0000000000018],[812.4999999999995,1745.0000000000018]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[754.7008330000026,1909.1917939999958],"typeId":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"instanceId":"00e3d6c2-f801-4d91-ad4d-237bada773bb","orientation":"up","circleData":[[4277.5,4115],[1022.5000000000039,1924.9999999999943],[1022.5000000000039,1954.9999999999939]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3123.2036904999995,1157.474882],"typeId":"5ac8a9e5-bb24-45ef-9b03-1161364522fb","componentVersion":1,"instanceId":"1c19cc90-e27a-4c31-a566-dce6d12cc7bd","orientation":"up","circleData":[[2987.5,1145],[3259.5265,1145]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Main line\n(phase) - L\n(Enedis in France)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3292.519774875356,1084.5794073453549],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"8b4859a0-119b-4d24-8c3e-f008f1af2f35","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Main neutral - N\n(Enedis in France)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2953.4352836968415,1091.5820712351226],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"eb1dbc1c-94ee-4954-b264-2ba5f2bb6c04","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[-165.78929000000016,-12.081628000000478],"typeId":"25d95763-f48b-4a99-bdb2-8bb3b7ccff88","componentVersion":1,"instanceId":"99cae55d-e9c7-468a-acc3-dcac762056db","orientation":"down","circleData":[[-12.500000000000007,5.00000000000002],[-12.500000000000007,-9.999999999999979],[-12.500000000000004,-25.0000000000002],[-12.500000000000014,-39.99999999999994],[-350,5.000000000000049],[-350,-25.00000000000017],[-350,27.50000000000002],[-350,-55.00000000000037]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"CT Clamp for\nGrid Power (in/out)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[3407.007981255236,1407.136824464781],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"e5530feb-ce19-40b3-8da6-a6ca8e4b619a","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[2528.8436755,1583.142836],"typeId":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"instanceId":"060f78c2-f7c5-4b91-a54e-26722a6a6eb1","orientation":"up","circleData":[[2507.5,1430],[2544.3571255,1429.1428745],[2545.6428145,1755.2857490000001],[2509.6428145,1753.1428744999998]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[2768.8436755000002,1778.142836],"typeId":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"instanceId":"c483e859-dbe3-40ab-ad85-fdb0e9726a1e","orientation":"up","circleData":[[2747.5,1625],[2784.3571255000006,1624.1428745],[2785.6428145,1950.2857490000008],[2749.6428145,1948.1428745000005]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1217.8757440000002,806.7131704999999],"typeId":"21a0a3b7-bfd8-4958-92f9-fb21adb71ce0","componentVersion":1,"instanceId":"d7e83964-79f2-4e6f-ab07-dee67fd9dff8","orientation":"right","circleData":[[1247.5,650],[1228.2216325000002,649.5517129999998],[1207.5982270000002,649.5517129999998],[1187.4231685,648.6550204999999],[1292.7818110000003,925.7259259999998],[1216.5649210000001,924.3808864999999],[1141.2446650000002,923.0359054999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1667.8757440000002,806.7131704999999],"typeId":"21a0a3b7-bfd8-4958-92f9-fb21adb71ce0","componentVersion":1,"instanceId":"6bde5401-8877-4618-b129-167654a129ea","orientation":"right","circleData":[[1697.5,650],[1678.2216325000002,649.5517129999998],[1657.5982270000002,649.5517129999998],[1637.4231685,648.6550204999999],[1742.7818110000003,925.7259259999998],[1666.5649210000001,924.3808864999999],[1591.2446650000002,923.0359055000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"N","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[153.35924144430763,655.2637795986317],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"786922c4-3cc4-4e2e-a1af-6f582a726cc5","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"L","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[257.0687211747471,655.9967802938984],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"c6b89f01-cd33-4f53-a410-bd8ce0a19726","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[468.922115048887,1657.2346746943958],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"028c5ed6-a9ce-4916-bd5a-20a0af91ff53","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"LOAD 2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[685.3637402494104,1881.2640404554054],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"d8ee4efe-302f-41eb-a87d-4235620299ce","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Dimmer\nOutput 2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1023.8439203020007,795.1529920546972],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"8c415f8f-024b-42a7-9906-fa5d9103b190","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Dimmer\nOutput 1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[1483.0932434380895,794.8020298127515],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"f0886e27-8ec0-43da-a659-1cbab4912d9c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Channel 2\nGrid Power","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2235.7808942171437,256.4715337095425],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"265be517-7dce-4507-b222-49efa0b79d44","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Channel 1:\nAll Output Power","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2046.6998402833278,257.233205403509],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"4d6635ca-f74e-4111-b736-96f73dea815d","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"Channel 1 clamp\naround all input \nphase wires (L)","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[2346.984033092402,1941.0591972016282],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"34d49454-fe1f-4693-a2f3-2121a541126c","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1047.6447520000002,1153.0044469999993],"typeId":"2ce95dbd-bb8b-430f-8511-f580783f914c","componentVersion":1,"instanceId":"320ab8ff-f5d3-4096-b4aa-da43287dff93","orientation":"right","circleData":[[1037.5,1250],[1022.5,1257.5]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1512.6447520000006,1378.004446999999],"typeId":"2ce95dbd-bb8b-430f-8511-f580783f914c","componentVersion":1,"instanceId":"d008a2f8-2853-4c0d-8d67-a8220f145d26","orientation":"right","circleData":[[1502.5,1475],[1487.5,1482.5]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"PZEM Output 1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[-162.67117562189352,-360.85974684688705],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"cabc8f6d-4e36-40d8-b46e-f81e3606417d","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Comment":{"version":2,"id":"Comment","label":"Comment","description":"","units":"","type":"string","value":"PZEM Output 2","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"Comment","unit":"","required":true},"backgroundColor":{"version":2,"id":"backgroundColor","label":"backgroundColor","description":"","units":"","type":"string","value":"#FFFFFF","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundColor","unit":"","required":true},"backgroundOpacity":{"version":2,"id":"backgroundOpacity","label":"backgroundOpacity","description":"","units":"","type":"decimal","value":"1","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"backgroundOpacity","unit":"","required":true},"textColor":{"version":2,"id":"textColor","label":"textColor","description":"","units":"","type":"string","value":"#000000","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"textColor","unit":"","required":true},"fontSize":{"version":2,"id":"fontSize","label":"fontSize","description":"","units":"","type":"integer","value":"16","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"fontSize","unit":"","required":true},"font":{"version":2,"id":"font","label":"font","description":"","units":"","type":"string","value":"Courier New","displayFormat":"input","showOnComp":false,"isVisibleToUser":true,"name":"font","unit":"","required":true}},"position":[-172.22891391829182,-119.31184204440922],"typeId":"458264b2-a399-d1b4-4e83-61faa437620f","componentVersion":1,"instanceId":"0532153d-ec59-4dd7-ad03-6d0401cd55c5","orientation":"up","circleData":[],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[3006.71431,2014.5000244999999],"typeId":"5ce5e9a0-0484-4e7a-b171-46d0c4edfd48","componentVersion":2,"instanceId":"9b271475-bebe-41b8-aded-20e21ef4734b","orientation":"up","circleData":[[2987.5,1850],[3029.499982,1850.8571344999998],[2986.6428895,2182.999983499998],[3030.7857474999996,2183.8571599999987]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-484.25286","left":"-372.27002","width":"4663.77002","height":"4613.25286","x":"-372.27002","y":"-484.25286"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_24\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"213.0759055000_396.3743885000\\\",\\\"212.5000000000_396.3743885000\\\",\\\"212.5000000000_12.5282165000\\\",\\\"679.1613940000_12.5282165000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawStartPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_0\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1967.5000000000_395.0000000000\\\",\\\"212.5000000000_395.0000000000\\\",\\\"212.5000000000_350.0000000000\\\",\\\"213.0759055000_350.0000000000\\\",\\\"213.0759055000_396.3743885000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawStartPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_3\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-12.5000000000_-40.0000000000\\\",\\\"212.5000000000_-40.0000000000\\\",\\\"212.5000000000_396.3743885000\\\",\\\"213.0759055000_396.3743885000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_3\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-12.5000000000_-280.0000000000\\\",\\\"212.5000000000_-280.0000000000\\\",\\\"212.5000000000_396.3743885000\\\",\\\"213.0759055000_396.3743885000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"213.0759055000_396.3743885000\\\",\\\"213.0759055000_395.0000000000\\\",\\\"1228.2216325000_395.0000000000\\\",\\\"1228.2216325000_649.5517130000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_1\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1678.2216325000_649.5517130000\\\",\\\"1678.2216325000_395.0000000000\\\",\\\"213.0759055000_395.0000000000\\\",\\\"213.0759055000_396.3743885000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_19\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"197.5000000000_395.0000000000\\\",\\\"197.5000000000_335.0000000000\\\",\\\"678.5382805000_335.0000000000\\\",\\\"678.5382805000_148.1934635000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawStartPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_1\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1967.9580910000_425.0000000000\\\",\\\"1907.5000000000_425.0000000000\\\",\\\"1907.5000000000_335.0000000000\\\",\\\"197.5000000000_335.0000000000\\\",\\\"197.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawStartPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_0\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-12.5000000000_5.0000000000\\\",\\\"182.5000000000_5.0000000000\\\",\\\"182.5000000000_335.0000000000\\\",\\\"197.5000000000_335.0000000000\\\",\\\"197.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_0\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-12.5000000000_-235.0000000000\\\",\\\"197.5000000000_-235.0000000000\\\",\\\"197.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0\",\"rawStartPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"197.5000000000_395.0000000000\\\",\\\"197.5000000000_335.0000000000\\\",\\\"1247.5000000000_335.0000000000\\\",\\\"1247.5000000000_650.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_0\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1697.5000000000_650.0000000000\\\",\\\"1697.5000000000_335.0000000000\\\",\\\"197.5000000000_335.0000000000\\\",\\\"197.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#FFA6FE\",\"startPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11\",\"rawStartPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_3\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_11\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1967.5000000000_492.5000000000\\\",\\\"1847.5000000000_492.5000000000\\\",\\\"1847.5000000000_-44.4230995000\\\",\\\"949.3291135000_-44.4230995000\\\"]}\"}","{\"color\":\"#774D00\",\"startPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10\",\"rawStartPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_2\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1967.5000000000_455.0000000000\\\",\\\"1877.5000000000_455.0000000000\\\",\\\"1877.5000000000_-71.6853940000\\\",\\\"949.3291135000_-71.6853940000\\\"]}\"}","{\"color\":\"#B500FF\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_2\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-12.5000000000_-265.0000000000\\\",\\\"347.5000000000_-265.0000000000\\\",\\\"347.5000000000_-43.2425995000\\\",\\\"679.1613940000_-43.2425995000\\\"]}\"}","{\"color\":\"#B500FF\",\"startPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26\",\"rawStartPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_2\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_26\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-12.5000000000_-25.0000000000\\\",\\\"347.5000000000_-25.0000000000\\\",\\\"347.5000000000_-43.2425995000\\\",\\\"679.1613940000_-43.2425995000\\\"]}\"}","{\"color\":\"#FFB167\",\"startPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27\",\"rawStartPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_1\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-12.5000000000_-10.0000000000\\\",\\\"370.0000000000_-10.0000000000\\\",\\\"370.0000000000_-70.4832805000\\\",\\\"677.9352805000_-70.4832805000\\\"]}\"}","{\"color\":\"#FFB167\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_1\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_27\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-12.5000000000_-250.0000000000\\\",\\\"370.0000000000_-250.0000000000\\\",\\\"370.0000000000_-70.4832805000\\\",\\\"677.9352805000_-70.4832805000\\\"]}\"}","{\"color\":\"#FFDB66\",\"startPinId\":\"pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0\",\"endPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10\",\"rawStartPinId\":\"pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_0\",\"rawEndPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_10\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3407.5000000000_1190.0000000000\\\",\\\"3407.5000000000_972.5000000000\\\",\\\"2230.6180000000_972.5000000000\\\",\\\"2230.6180000000_310.8395000000\\\"]}\"}","{\"color\":\"#90FB92\",\"startPinId\":\"pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1\",\"endPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9\",\"rawStartPinId\":\"pin-type-component_7cf7ad7f-dee5-4409-b6bd-1e28c1d7dc2a_1\",\"rawEndPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_9\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3422.5000000000_1182.5000000000\\\",\\\"3422.5000000000_995.0000000000\\\",\\\"2206.8475000000_995.0000000000\\\",\\\"2206.8475000000_310.3925000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2987.5000000000_1145.0000000000\\\",\\\"2747.5000000000_1145.0000000000\\\",\\\"2747.5000000000_1625.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0\",\"endPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_0\",\"rawEndPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2507.5000000000_1430.0000000000\\\",\\\"2507.5000000000_1145.0000000000\\\",\\\"2987.5000000000_1145.0000000000\\\"]}\"}","{\"color\":\"#0076FF\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"endPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_0\",\"rawEndPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2987.5000000000_1145.0000000000\\\",\\\"2987.5000000000_1850.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1\",\"endPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_1\",\"rawEndPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2544.3571255000_1429.1428745000\\\",\\\"2544.3571255000_1310.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3259.5265000000_1145.0000000000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3259.5265000000_1145.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"2784.3571255000_1310.0000000000\\\",\\\"2784.3571255000_1624.1428745000\\\"]}\"}","{\"color\":\"#85A900\",\"startPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"endPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1\",\"rawStartPinId\":\"pin-type-component_1c19cc90-e27a-4c31-a566-dce6d12cc7bd_1\",\"rawEndPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3259.5265000000_1145.0000000000\\\",\\\"3317.5000000000_1145.0000000000\\\",\\\"3317.5000000000_1310.0000000000\\\",\\\"3032.5000000000_1310.0000000000\\\",\\\"3032.5000000000_1850.8571345000\\\",\\\"3029.4999820000_1850.8571345000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6\",\"endPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6\",\"rawEndPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-350.0000000000_-212.5000000000\\\",\\\"-560.0000000000_-212.5000000000\\\",\\\"-560.0000000000_27.5000000000\\\",\\\"-350.0000000000_27.5000000000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6\",\"endPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_6\",\"rawEndPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-350.0000000000_-212.5000000000\\\",\\\"-560.0000000000_-212.5000000000\\\",\\\"-560.0000000000_2247.5000000000\\\",\\\"2986.6428895000_2247.5000000000\\\",\\\"2986.6428895000_2182.9999835000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"endPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6\",\"rawStartPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"rawEndPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2986.6428895000_2182.9999835000\\\",\\\"2986.6428895000_2247.5000000000\\\",\\\"3625.0000000000_2247.5000000000\\\",\\\"3625.0000000000_462.5000000000\\\",\\\"2305.0000000000_462.5000000000\\\"]}\"}","{\"color\":\"#00FFC6\",\"startPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3\",\"rawStartPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_2\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2986.6428895000_2182.9999835000\\\",\\\"2986.6428895000_2247.5000000000\\\",\\\"197.5000000000_2247.5000000000\\\",\\\"197.5000000000_650.6282870000\\\",\\\"200.7068110000_650.6282870000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4\",\"endPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4\",\"rawEndPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-350.0000000000_-235.0000000000\\\",\\\"-590.0000000000_-235.0000000000\\\",\\\"-590.0000000000_5.0000000000\\\",\\\"-350.0000000000_5.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4\",\"endPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_4\",\"rawEndPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-350.0000000000_-235.0000000000\\\",\\\"-590.0000000000_-235.0000000000\\\",\\\"-590.0000000000_2277.5000000000\\\",\\\"3032.5000000000_2277.5000000000\\\",\\\"3032.5000000000_2183.8571600000\\\",\\\"3030.7857475000_2183.8571600000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"endPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5\",\"rawStartPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"rawEndPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3030.7857475000_2183.8571600000\\\",\\\"3030.7857475000_2277.5000000000\\\",\\\"3662.5000000000_2277.5000000000\\\",\\\"3662.5000000000_410.0000000000\\\",\\\"2305.0000000000_410.0000000000\\\"]}\"}","{\"color\":\"#FF6E41\",\"startPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"endPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2\",\"rawStartPinId\":\"pin-type-component_9b271475-bebe-41b8-aded-20e21ef4734b_3\",\"rawEndPinId\":\"pin-type-component_d53bc8d1-adbf-42c3-9bdc-27d4d2b68588_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"3030.7857475000_2183.8571600000\\\",\\\"3032.5000000000_2183.8571600000\\\",\\\"3032.5000000000_2277.5000000000\\\",\\\"213.9921460000_2277.5000000000\\\",\\\"213.9921460000_649.2539555000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"endPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"rawEndPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2509.6428145000_1753.1428745000\\\",\\\"2509.6428145000_1820.0000000000\\\",\\\"1666.5649210000_1820.0000000000\\\",\\\"1666.5649210000_924.3808865000\\\"]}\"}","{\"color\":\"#E85EBE\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"endPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_3\",\"rawEndPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2509.6428145000_1753.1428745000\\\",\\\"2509.6428145000_1820.0000000000\\\",\\\"812.5000000000_1820.0000000000\\\",\\\"812.5000000000_1745.0000000000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5\",\"rawStartPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2749.6428145000_1948.1428745000\\\",\\\"2749.6428145000_2172.5000000000\\\",\\\"1216.5649210000_2172.5000000000\\\",\\\"1216.5649210000_924.3808865000\\\"]}\"}","{\"color\":\"#010067\",\"startPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2\",\"endPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"rawStartPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_2\",\"rawEndPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_1955.0000000000\\\",\\\"1022.5000000000_2172.5000000000\\\",\\\"2749.6428145000_2172.5000000000\\\",\\\"2749.6428145000_1948.1428745000\\\"]}\"}","{\"color\":\"#9E008E\",\"startPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2\",\"endPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4\",\"rawStartPinId\":\"pin-type-component_060f78c2-f7c5-4b91-a54e-26722a6a6eb1_2\",\"rawEndPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2545.6428145000_1755.2857490000\\\",\\\"2545.6428145000_2082.5000000000\\\",\\\"1742.5000000000_2082.5000000000\\\",\\\"1742.5000000000_925.7259260000\\\",\\\"1742.7818110000_925.7259260000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4\",\"rawStartPinId\":\"pin-type-component_c483e859-dbe3-40ab-ad85-fdb0e9726a1e_2\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2785.6428145000_1950.2857490000\\\",\\\"2785.0000000000_1950.2857490000\\\",\\\"2785.0000000000_2097.5000000000\\\",\\\"1292.7818110000_2097.5000000000\\\",\\\"1292.7818110000_925.7259260000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6\",\"endPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_6\",\"rawEndPinId\":\"pin-type-component_ee3599dd-7cc8-4121-aeb8-3fd6e229f0c8_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1591.2446650000_923.0359055000\\\",\\\"1591.2446650000_1715.0000000000\\\",\\\"812.5000000000_1715.0000000000\\\"]}\"}","{\"color\":\"#005F39\",\"startPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1\",\"endPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6\",\"rawStartPinId\":\"pin-type-component_00e3d6c2-f801-4d91-ad4d-237bada773bb_1\",\"rawEndPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_6\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_1925.0000000000\\\",\\\"1141.2446650000_1925.0000000000\\\",\\\"1141.2446650000_923.0359055000\\\"]}\"}","{\"color\":\"#95003A\",\"startPinId\":\"pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1\",\"endPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7\",\"rawStartPinId\":\"pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_1\",\"rawEndPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2110.0000000000_1985.0000000000\\\",\\\"2054.1325000000_1985.0000000000\\\",\\\"2054.1325000000_309.5015000000\\\"]}\"}","{\"color\":\"#FF937E\",\"startPinId\":\"pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0\",\"endPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8\",\"rawStartPinId\":\"pin-type-component_1a4c0ab2-15d7-4f55-82c5-02526f5965a4_0\",\"rawEndPinId\":\"pin-type-component_ae19664f-1584-4f12-9c79-f0e8930ce70b_8\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"2117.5000000000_2000.0000000000\\\",\\\"2080.0000000000_2000.0000000000\\\",\\\"2080.0000000000_552.5000000000\\\",\\\"2079.5350000000_552.5000000000\\\",\\\"2079.5350000000_308.6105000000\\\"]}\"}","{\"color\":\"#001544\",\"startPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28\",\"rawStartPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_3\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_28\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1187.4231685000_648.6550205000\\\",\\\"1187.4231685000_-467.5000000000\\\",\\\"550.0000000000_-467.5000000000\\\",\\\"550.0000000000_-95.9164615000\\\",\\\"677.9352805000_-95.9164615000\\\"]}\"}","{\"color\":\"#91D0CB\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_3\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_29\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1637.4231685000_648.6550205000\\\",\\\"1637.4231685000_-497.5000000000\\\",\\\"587.5000000000_-497.5000000000\\\",\\\"587.5000000000_-121.9526425000\\\",\\\"677.3322805000_-121.9526425000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32\",\"rawStartPinId\":\"pin-type-component_d7e83964-79f2-4e6f-ab07-dee67fd9dff8_2\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1207.5982270000_649.5517130000\\\",\\\"1207.5982270000_-527.5000000000\\\",\\\"617.5000000000_-527.5000000000\\\",\\\"617.5000000000_-203.7140260000\\\",\\\"678.5583940000_-203.7140260000\\\"]}\"}","{\"color\":\"#007DB5\",\"startPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2\",\"endPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32\",\"rawStartPinId\":\"pin-type-component_6bde5401-8877-4618-b129-167654a129ea_2\",\"rawEndPinId\":\"pin-type-component_f7d25e04-bb51-41df-ba72-c452c270d3fb_32\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1657.5982270000_649.5517130000\\\",\\\"1657.5982270000_-527.5000000000\\\",\\\"617.5000000000_-527.5000000000\\\",\\\"617.5000000000_-203.7140260000\\\",\\\"678.5583940000_-203.7140260000\\\"]}\"}","{\"color\":\"#6A826C\",\"startPinId\":\"pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0\",\"endPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5\",\"rawStartPinId\":\"pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_0\",\"rawEndPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1037.5000000000_1250.0000000000\\\",\\\"1037.5000000000_1325.0000000000\\\",\\\"-410.0000000000_1325.0000000000\\\",\\\"-410.0000000000_-25.0000000000\\\",\\\"-350.0000000000_-25.0000000000\\\"]}\"}","{\"color\":\"#00AE7E\",\"startPinId\":\"pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1\",\"endPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7\",\"rawStartPinId\":\"pin-type-component_320ab8ff-f5d3-4096-b4aa-da43287dff93_1\",\"rawEndPinId\":\"pin-type-component_99cae55d-e9c7-468a-acc3-dcac762056db_7\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1022.5000000000_1257.5000000000\\\",\\\"1022.5000000000_1302.5000000000\\\",\\\"-387.5000000000_1302.5000000000\\\",\\\"-387.5000000000_-55.0000000000\\\",\\\"-350.0000000000_-55.0000000000\\\"]}\"}","{\"color\":\"#C28C9F\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5\",\"endPinId\":\"pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_5\",\"rawEndPinId\":\"pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-350.0000000000_-265.0000000000\\\",\\\"-485.0000000000_-265.0000000000\\\",\\\"-485.0000000000_1535.0000000000\\\",\\\"1502.5000000000_1535.0000000000\\\",\\\"1502.5000000000_1475.0000000000\\\"]}\"}","{\"color\":\"#008F9C\",\"startPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7\",\"endPinId\":\"pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1\",\"rawStartPinId\":\"pin-type-component_22500cd3-352c-4d79-9f9c-f48cf0a80685_7\",\"rawEndPinId\":\"pin-type-component_d008a2f8-2853-4c0d-8d67-a8220f145d26_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"-350.0000000000_-295.0000000000\\\",\\\"-462.5000000000_-295.0000000000\\\",\\\"-462.5000000000_1512.5000000000\\\",\\\"1487.5000000000_1512.5000000000\\\",\\\"1487.5000000000_1482.5000000000\\\"]}\"}"],"projectDescription":""}PK
     mdZ               jsons/PK
     mdZ�E\��  ��     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"HDR-15-5 5V 2.4A","category":["User Defined"],"id":"c2a09f2b-df40-42a6-8e0c-c519ba38e9d5","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.png","iconPic":"7b19d218-2217-455d-9a43-b73a208c2c5c.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"3.54331","numDisplayRows":"21.25984","pins":[{"uniquePinIdString":"0","positionMil":"144.79685,1962.29409","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"248.63622,1953.13150","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"254.74449,267.26772","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"166.17559,258.10551","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"PZEM-004T V3","category":["User Defined"],"id":"25d95763-f48b-4a99-bdb2-8bb3b7ccff88","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"7139d0cb-a6f6-4338-81e1-1177b1f79563.png","iconPic":"e77f5de3-b891-4dea-bd4b-a791874bc34b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"26.19743","numDisplayRows":"11.64330","pins":[{"uniquePinIdString":"0","positionMil":"287.94290,696.04252","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"287.94290,596.04252","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"2","positionMil":"287.94290,496.04252","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"3","positionMil":"287.94290,396.04252","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"2537.94290,696.04252","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"5","positionMil":"2537.94290,496.04252","isAnchorPin":false,"label":"CT-"},{"uniquePinIdString":"6","positionMil":"2537.94290,846.04252","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"7","positionMil":"2537.94290,296.04252","isAnchorPin":false,"label":"CT+"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Current Tranformer","category":["User Defined"],"id":"2ce95dbd-bb8b-430f-8511-f580783f914c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e975526f-cfd2-4a7e-88b6-747cffbdf2da.png","iconPic":"2fc28fee-789f-4880-bf44-0d05ccb6f4b5.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"20.31772","numDisplayRows":"20.31772","pins":[{"uniquePinIdString":"0","positionMil":"1662.52302,948.25432","isAnchorPin":true,"label":"Negative"},{"uniquePinIdString":"1","positionMil":"1712.52302,848.25432","isAnchorPin":false,"label":"Positive"}],"pinType":"wired"},"properties":[]},{"subtypeName":"JSY-MK-194G","category":["User Defined"],"id":"840a331c-2aef-4dd8-892c-7ae81d6bcea5","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"9bf2961f-aa36-488c-987a-2819190a8ab9.png","iconPic":"446f47db-f7ac-4e06-8ce0-bf970f803875.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"25.59055","numDisplayRows":"18.89764","pins":[{"uniquePinIdString":"0","positionMil":"112.85748,1211.55197","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"115.91142,1011.55197","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"2","positionMil":"112.85748,811.55197","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"3","positionMil":"112.85748,561.55197","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"4","positionMil":"1062.85748,61.55197","isAnchorPin":false,"label":""},{"uniquePinIdString":"5","positionMil":"2362.85748,1111.55197","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"6","positionMil":"2362.85748,761.55197","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"7","positionMil":"690.40748,1781.54197","isAnchorPin":false,"label":"CT1+"},{"uniquePinIdString":"8","positionMil":"859.75748,1787.48197","isAnchorPin":false,"label":"CT1-"},{"uniquePinIdString":"9","positionMil":"1708.50748,1775.60197","isAnchorPin":false,"label":"CT2+"},{"uniquePinIdString":"10","positionMil":"1866.97748,1772.62197","isAnchorPin":false,"label":"CT2-"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Current Tranformer","category":["User Defined"],"id":"2ce95dbd-bb8b-430f-8511-f580783f914c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e975526f-cfd2-4a7e-88b6-747cffbdf2da.png","iconPic":"2fc28fee-789f-4880-bf44-0d05ccb6f4b5.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"20.31772","numDisplayRows":"20.31772","pins":[{"uniquePinIdString":"0","positionMil":"1662.52302,948.25432","isAnchorPin":true,"label":"Negative"},{"uniquePinIdString":"1","positionMil":"1712.52302,848.25432","isAnchorPin":false,"label":"Positive"}],"pinType":"wired"},"properties":[]},{"subtypeName":"ESP32 Devkit V4","category":["User Defined"],"id":"b975acdd-73e3-4b18-a5a5-9b66f369afa0","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.png","iconPic":"cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"48.00864","numDisplayRows":"48.00864","pins":[{"uniquePinIdString":"0","positionMil":"3273.41401,3905.84495","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"3277.43401,3724.10632","isAnchorPin":false,"label":"23"},{"uniquePinIdString":"2","positionMil":"3277.56810,3550.53178","isAnchorPin":false,"label":"22"},{"uniquePinIdString":"3","positionMil":"3273.41401,3360.60905","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"4","positionMil":"3281.58810,3187.03451","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"5","positionMil":"3273.41401,3013.32588","isAnchorPin":false,"label":"21"},{"uniquePinIdString":"6","positionMil":"3281.58810,2827.55725","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"3281.58810,2653.98271","isAnchorPin":false,"label":"19"},{"uniquePinIdString":"8","positionMil":"3281.58810,2472.24408","isAnchorPin":false,"label":"18"},{"uniquePinIdString":"9","positionMil":"3277.43401,2302.84954","isAnchorPin":false,"label":"5"},{"uniquePinIdString":"10","positionMil":"3285.60810,2117.08091","isAnchorPin":false,"label":"17"},{"uniquePinIdString":"11","positionMil":"3285.60810,1935.33228","isAnchorPin":false,"label":"16"},{"uniquePinIdString":"12","positionMil":"3285.60810,1749.58956","isAnchorPin":false,"label":"4"},{"uniquePinIdString":"13","positionMil":"3289.61810,1576.02502","isAnchorPin":false,"label":"0"},{"uniquePinIdString":"14","positionMil":"3285.60810,1402.58457","isAnchorPin":false,"label":"2"},{"uniquePinIdString":"15","positionMil":"3293.78219,1208.50775","isAnchorPin":false,"label":"15"},{"uniquePinIdString":"16","positionMil":"3289.61810,1034.93321","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"17","positionMil":"3289.61810,849.03049","isAnchorPin":false,"label":"D0"},{"uniquePinIdString":"18","positionMil":"3301.95628,659.25186","isAnchorPin":false,"label":"CLK"},{"uniquePinIdString":"19","positionMil":"1480.33588,651.22186","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"20","positionMil":"1472.16179,836.98049","isAnchorPin":false,"label":"CMD"},{"uniquePinIdString":"21","positionMil":"1480.33588,1010.55503","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"22","positionMil":"1476.31588,1196.31366","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"23","positionMil":"1476.31588,1378.06229","isAnchorPin":false,"label":"13"},{"uniquePinIdString":"24","positionMil":"1484.48997,1555.65684","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"25","positionMil":"1480.33588,1733.38547","isAnchorPin":false,"label":"12"},{"uniquePinIdString":"26","positionMil":"1484.48997,1927.46228","isAnchorPin":false,"label":"14"},{"uniquePinIdString":"27","positionMil":"1476.31588,2109.06682","isAnchorPin":false,"label":"27"},{"uniquePinIdString":"28","positionMil":"1476.31588,2278.62136","isAnchorPin":false,"label":"26"},{"uniquePinIdString":"29","positionMil":"1472.29588,2452.19590","isAnchorPin":false,"label":"25"},{"uniquePinIdString":"30","positionMil":"1472.29588,2637.96453","isAnchorPin":false,"label":"33"},{"uniquePinIdString":"31","positionMil":"1472.16179,2815.53316","isAnchorPin":false,"label":"32"},{"uniquePinIdString":"32","positionMil":"1480.46997,2997.27179","isAnchorPin":false,"label":"35"},{"uniquePinIdString":"33","positionMil":"1472.29588,3170.71224","isAnchorPin":false,"label":"34"},{"uniquePinIdString":"34","positionMil":"1459.96384,3364.79179","isAnchorPin":false,"label":"VIN"},{"uniquePinIdString":"35","positionMil":"1472.29588,3534.47769","isAnchorPin":false,"label":"VP"},{"uniquePinIdString":"36","positionMil":"1476.31384,3711.93179","isAnchorPin":false,"label":"EN"},{"uniquePinIdString":"37","positionMil":"1472.29588,3897.67086","isAnchorPin":false,"label":"3V3"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Water Heater","category":["User Defined"],"id":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"85e66502-362d-4a26-afcd-97fbc4859675.png","iconPic":"b13518ba-21c5-4f60-a735-1d8041d11d7b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"39.37008","numDisplayRows":"39.37008","pins":[{"uniquePinIdString":"0","positionMil":"25453.83178,-12736.88404","isAnchorPin":true,"label":""},{"uniquePinIdString":"1","positionMil":"3753.83178,1863.11596","isAnchorPin":false,"label":"V+"},{"uniquePinIdString":"2","positionMil":"3753.83178,1663.11596","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Water Heater","category":["User Defined"],"id":"fa95e5d1-b92a-410f-a873-a71d0089e7ad","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"85e66502-362d-4a26-afcd-97fbc4859675.png","iconPic":"b13518ba-21c5-4f60-a735-1d8041d11d7b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"39.37008","numDisplayRows":"39.37008","pins":[{"uniquePinIdString":"0","positionMil":"25453.83178,-12736.88404","isAnchorPin":true,"label":""},{"uniquePinIdString":"1","positionMil":"3753.83178,1863.11596","isAnchorPin":false,"label":"V+"},{"uniquePinIdString":"2","positionMil":"3753.83178,1663.11596","isAnchorPin":false,"label":"V-"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Alternative Current (AC) - Large","category":["User Defined"],"id":"5ac8a9e5-bb24-45ef-9b03-1161364522fb","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"8a1d81a5-79d4-450c-9f72-108cd2673013.png","iconPic":"aacc0029-e57d-4614-a443-d9bee65b5175.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.63677","numDisplayRows":"22.90067","pins":[{"uniquePinIdString":"0","positionMil":"277.14723,1228.19938","isAnchorPin":true,"label":"Neutral"},{"uniquePinIdString":"1","positionMil":"2090.65723,1228.19938","isAnchorPin":false,"label":"Line"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"PZEM-004T V3","category":["User Defined"],"id":"25d95763-f48b-4a99-bdb2-8bb3b7ccff88","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"7139d0cb-a6f6-4338-81e1-1177b1f79563.png","iconPic":"e77f5de3-b891-4dea-bd4b-a791874bc34b.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"26.19743","numDisplayRows":"11.64330","pins":[{"uniquePinIdString":"0","positionMil":"287.94290,696.04252","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"287.94290,596.04252","isAnchorPin":false,"label":"RX"},{"uniquePinIdString":"2","positionMil":"287.94290,496.04252","isAnchorPin":false,"label":"TX"},{"uniquePinIdString":"3","positionMil":"287.94290,396.04252","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"4","positionMil":"2537.94290,696.04252","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"5","positionMil":"2537.94290,496.04252","isAnchorPin":false,"label":"CT-"},{"uniquePinIdString":"6","positionMil":"2537.94290,846.04252","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"7","positionMil":"2537.94290,296.04252","isAnchorPin":false,"label":"CT+"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Breaker 20A","category":["User Defined"],"id":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1d90a712-93d7-4555-ae10-1782f839eba3.png","iconPic":"e5551f5a-2fb7-4493-9527-57db21faeaae.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.69291","numDisplayRows":"28.74016","pins":[{"uniquePinIdString":"0","positionMil":"192.35433,2457.96024","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"438.06850,2463.67441","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"446.63976,289.38858","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"206.63976,303.67441","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Breaker 20A","category":["User Defined"],"id":"a64016c8-4d9c-491e-ba46-f626b2aeb38c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"1d90a712-93d7-4555-ae10-1782f839eba3.png","iconPic":"e5551f5a-2fb7-4493-9527-57db21faeaae.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.69291","numDisplayRows":"28.74016","pins":[{"uniquePinIdString":"0","positionMil":"192.35433,2457.96024","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"438.06850,2463.67441","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"446.63976,289.38858","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"3","positionMil":"206.63976,303.67441","isAnchorPin":false,"label":"N"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Robodyn 16/24A","category":["User Defined"],"id":"21a0a3b7-bfd8-4958-92f9-fb21adb71ce0","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ae036c7f-e258-4627-a75d-99715ec815e7.png","iconPic":"69c28b0d-a0ad-46f0-a190-03e6ecfe42fd.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.62205","numDisplayRows":"16.53543","pins":[{"uniquePinIdString":"0","positionMil":"136.34803,1024.26654","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"133.35945,895.74409","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"133.35945,758.25472","isAnchorPin":false,"label":"ZC"},{"uniquePinIdString":"3","positionMil":"127.38150,623.75433","isAnchorPin":false,"label":"PSM"},{"uniquePinIdString":"4","positionMil":"1974.52087,1326.14528","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"5","positionMil":"1965.55394,818.03268","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"6","positionMil":"1956.58740,315.89764","isAnchorPin":false,"label":"LOAD"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Robodyn 16/24A","category":["User Defined"],"id":"21a0a3b7-bfd8-4958-92f9-fb21adb71ce0","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"ae036c7f-e258-4627-a75d-99715ec815e7.png","iconPic":"69c28b0d-a0ad-46f0-a190-03e6ecfe42fd.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.62205","numDisplayRows":"16.53543","pins":[{"uniquePinIdString":"0","positionMil":"136.34803,1024.26654","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"133.35945,895.74409","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"2","positionMil":"133.35945,758.25472","isAnchorPin":false,"label":"ZC"},{"uniquePinIdString":"3","positionMil":"127.38150,623.75433","isAnchorPin":false,"label":"PSM"},{"uniquePinIdString":"4","positionMil":"1974.52087,1326.14528","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"5","positionMil":"1965.55394,818.03268","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"6","positionMil":"1956.58740,315.89764","isAnchorPin":false,"label":"LOAD"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Current Tranformer","category":["User Defined"],"id":"2ce95dbd-bb8b-430f-8511-f580783f914c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e975526f-cfd2-4a7e-88b6-747cffbdf2da.png","iconPic":"2fc28fee-789f-4880-bf44-0d05ccb6f4b5.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"20.31772","numDisplayRows":"20.31772","pins":[{"uniquePinIdString":"0","positionMil":"1662.52302,948.25432","isAnchorPin":true,"label":"Negative"},{"uniquePinIdString":"1","positionMil":"1712.52302,848.25432","isAnchorPin":false,"label":"Positive"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Current Tranformer","category":["User Defined"],"id":"2ce95dbd-bb8b-430f-8511-f580783f914c","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"e975526f-cfd2-4a7e-88b6-747cffbdf2da.png","iconPic":"2fc28fee-789f-4880-bf44-0d05ccb6f4b5.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"20.31772","numDisplayRows":"20.31772","pins":[{"uniquePinIdString":"0","positionMil":"1662.52302,948.25432","isAnchorPin":true,"label":"Negative"},{"uniquePinIdString":"1","positionMil":"1712.52302,848.25432","isAnchorPin":false,"label":"Positive"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Comment","category":["Basic"],"userDefined":false,"id":"458264b2-a399-d1b4-4e83-61faa437620f","subtypeDescription":"","subtypePic":"8c2f1315-cf23-4ba8-a920-becb97f13280.png","pinInfo":{"numPins":"0","polarity":[],"pinType":"movable"},"properties":[{"type":"string","name":"Comment","value":"text box (double-click to edit)","unit":"","required":true},{"type":"polarity","name":"polarity","value":[],"unit":"","showOnComp":false,"required":true,"flipComponentPicWithPolarity":false},{"type":"","name":"backgroundColor","value":"#FFFFFF","unit":"","required":true},{"type":"","name":"backgroundOpacity","value":1,"unit":"","required":true},{"type":"","name":"textColor","value":"#000000","unit":"","required":true},{"type":"","name":"fontSize","value":10,"unit":"","required":true},{"type":"","name":"font","value":"Courier New","unit":"","required":true}],"iconPic":"6fc4b800-efc3-4a5d-827d-9566cfd108b3.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Breaker 2A","category":["User Defined"],"id":"5ce5e9a0-0484-4e7a-b171-46d0c4edfd48","componentVersion":2,"userDefined":true,"subtypeDescription":"","subtypePic":"a038ca8d-f9eb-4e93-ad0b-b831193aa106.png","iconPic":"3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.66667","numDisplayRows":"28.33333","pins":[{"uniquePinIdString":"0","positionMil":"205.23810,2513.33333","isAnchorPin":true,"label":"N"},{"uniquePinIdString":"1","positionMil":"485.23798,2507.61910","isAnchorPin":false,"label":"L"},{"uniquePinIdString":"2","positionMil":"199.52403,293.33344","isAnchorPin":false,"label":"N"},{"uniquePinIdString":"3","positionMil":"493.80975,287.61893","isAnchorPin":false,"label":"L"}],"pinType":"wired"},"properties":[]}]}PK
     mdZ               images/PK
     mdZ3��C� � /   images/cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.png�PNG

   IHDR  R  ~   �,  0�iCCPICC Profile  x��||eE���6�ѫt�q�"�����ٰD�ݐd�b	!��l#[`a�.  m�"M�(E�HS�. � MP����ܙ;�w�������w��L;s���;�%ɾc�,�3��$s�-�<��Ǟ{UWz%���K6Jt���-]]	~���{,i��G�i����g����a~���a����_:`���'�}�s��Dc���!z��G��xrzS����
:�jKf����d�:�Ë&ɪ]�i�=<�2���м����3�Θ�$�A"ɬ9���>�Ɯ;����I2��E�ó�dm����}F�5k���6)�L\R��~��.Ӻ���nU�2֜�ff����[��78<4�M�$%Ӵ)KӁsY���L�M�M=Mف����n�ٻG�e�'+�iIW��d��-��N�˒f�J���֎�5��׭�Y�`2���P2�l�4�]�3�M�^�����gI�Ԯ�� T'~{\ˁs1�Y�ѶE{oR,���g�����u����C�f/��@����jM$=	�Bos��;}l���-!����b�$I�`�!������d��c��$k��$��@�y�S��������������)�9�%ɵ�m�ɓɫ��6l� vmاaY���6<��ڨ5Fe���:d�e��]����G_<��1��sژ'�n6v��+��s�wĸV�x�y+�v�MV^��C�LX�;�<Va�+�:c�?�ֹ�]���~�z����rͳ�Zk��������:����i�m����w����~a�/\�aۆ�耍����M��ț�n6c�7p�c��_L�x[�_j����O8cˁ���국��f�/o�����iv��k�}�/��u�|~�8X�Q{���Nݮ�ӷ��C;���_;�岉��>:�;�<y�]���~���t����ԍ�Zw[�}i����O���5{��k�7���ߞ�w��o���)3���f>��}���y��_����^�xs�p���]v�w�:����>��#78���s���vܣ'�w⸓.8����O;��	g����g�t�%�u���Oν���]���W^~�{������|r�S�����r�W�ܺ�����o��󮻮����N|��<<���?^���lz��g|n�秼8��^���]_�ፉo���x�����^�тO��_�?����ڕ\�|���pݨG6��3p�{�ye�A��w�J3W����*7W�^���[��5�Ys�Z�}�:����z^��>�p��&l��&{l�x�S7���W_nL���MZ���լ��ns���������=���7�x�XY���כ�-l�v[5�~�vޱ{����������^8麶;w~l�K������n�!;w�2w�q]��vo�+�+O�j�.����=��/���7_�֊���޺�}��͘3�p���3����{�~WϹ}�C���O�W]�ɢ���/����Z���c>c�%߹��������#�Q����ѳ�Y|�����q?<��.��U'^{�/N����N�|�����?9��3�8�Գ~�c�>�C�=��_��?�`���h�O�^<��/�x�֗�}E�\��U�|�Օkֽv������冎w����C7/�ղ[�����κ��;����~s�o���߽|�w�{���������~�؃?t��w���G��g���������'>�������̎��n������^���F�<�o+�����������vx}�o.}��^����<��'�����>��Ã����n���c��_���a��Fm:�Q���Yc�{����ݱ҂��]����U�d��V;~���8u��ֺb�׹g���{q���0z��7�z�6�}��7;a�K�������Ҹ�Mh�r���n��6�|�'7����[�ro�x�{��-���JfU��v|u���A�زӔ�}�e��C[O���kv���Gwy���]+_���ީ�N���{^�6f���'�����W~����ӷ��{l�&�dm3�����x��C��{�~�Ϲ{�S�^_����٢�Ż/�}�A�����:��e���{�*�m~8;���ݏ����>�S�=���w��p�9�铞;��S^:��察���>��3�;���>�чgp��~x�G���@�%}���.��%���ν��+��򰫎��q??��3����+���w\�����M�����o�ආ�+w����~��o�;w�]�]�w��Y�ιo���>0�����!��c9�ѓ�x�c�?������'yj��s����������em|~�ƾ����x�ٗ��ݯ������?.{���/~�7�x�ތ��ݿ��ƿV|�����m>��x�'�$:�%�5Lj8���Q{��{�}��1?��7��m��+����U6Z����V�r��V?s���<�K׾v��ֽ�����+�_�x�&6]��M�?S�ŭw����O8g��zh뗷�x����m�X��+��˲�ٙ�"q��Uݣ5�ؿm���cvXw�	;�u�̘����I���z�?M~�}��7��t�޹tʏ����\��	���L?b���͞��⛛|K~{J߬��?}�+n����3�����7�>�o�9��m��������?|���.^��%���_?(9x�e㿣���C�]r�I�_r��G>~�kG7�ޱ�/�k9��=~0p�ܓ�|�)�N���CO;�G�~�ǜy�Y��踳O<�sO?����~r��_x�E����G.��e?���+����ّ??���9�ڳ���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\���<���O�磟9�/�?{�s�����x�{/��i/���K_���;���?����o���Vo���޷�}��w��w�n|������~壷>��'� rX8��< �8!I&�+�jŊ��N��]e��X��I�J�s�I�����I2�KI"�a��g�ly0�j9.͹�g�G��1����Ã���צ�L?h�C'�Y<���Z�ޕv�8IF`��'�utT=`M�?���iI2p�{�14��V��@���u�5x� ��������������v`�dc����ߍW��U!pS�0�0{��_�+p|zT/^'����gԅx����xm��7z{�~o�~��ܿ�~��W�zF?�W�3&w�ok��9�v2�@���z�3��i/VJ������hq�>�[�P�Bp�OH%8�����/���� \�������p�e
Ҝ.p�j���|��n]	��Š�o��?If�����W[2%iǘ���|�|�En����&��[S�p,D�2�:�L8�=Ȁ�Au��z�c8���!O��e���7�} �s�;�5-�:��g��?�?�2�\�M#V���+i��A��"N��tm�Aw���$%30����@f$#:W������S�7i�D�� ����?�!� s?�4�@;��J�8�-��SX����e��|�I|�?o:��1� $�)sd���2���K���gA�qs������l��g��A�s�"��m��j�R��������;����2<k�9���9C��/�?���?<kpQu`v���м����������ۧ���:ch�������޶I�ƞ�E����Uf���N��$sՁFL=�����������8�����e��JO���m}��;�zzۺ�'��vv�M�n۳h� ��:z��;�v�u�uU�'O�n���tOn��k����=��mJo�q���E�ա�:	K�ӿ�kx~S�u���Ý���7���|]}�{v�aܝ��zv�6N����Ll�i�k�~��J�(�[OW[kowKGޭcZ'�6;���Z'u�j�5�eƤUkk�k��j��Z��e��2ejwgKG�^m��z���ٗ�i�q϶�����ImS�:�����abwKo��)}]S{z�'v�y���6�TİgGGD��=ugz�Si^Rm�v�����܊ί��D�ڊ�\48�z�Т�A"���k�fk��?oF5?��Ξ*�e5�Xm��a�����)�J�L����=���Y���H�A�;ZZw��!?:��)=nW~3��sw7d�������.�8�����3��z �jc3���s���]F0u������Ӷ۴6K�qjWo{'���	c���S�4�T�2eZ�Ķ�>ld����I=U�E<����og:��JOKgW�S
��n��d���I������������#��i��fZ����A?�c��V�2���'[�F�
+a�ҽ�U�jt�W���^U�ƅIU�����~�������8���R-2�YiҊ�����~�f��k�q����O�����2��~�	f��ʚf�[�O0�
Q1Qz��8(���8:���'%�JM��=����&2�9�Ei)h�V)�T���c�e�k<�R��<2Z�Hוl�����AGͳ*�]��(4�M%�2����*�)�s]iMs�Y4�q����u�r+5�`�Iiy5n�E�م�Y-�)�@g�٪�%�#�%�_������Ό��Ԡ<F�J�J��X�05e��T�B�)����U%�%�1rנ�*Nf$3T/�i%C8ľS�v�Y��̬#�J�F�-6bY�܎>K�MX�6�1�HJ�H�U��&�2l�p�4[��M-5�$*���NA�� �Ժ#��e�F���ƪ�fRn����I�2G.�R�H��
<P�C�G%�Lf��5!�$��j�x�י��5��56��@���0�)l�8�z�k��~��R�Sk+p
��Q�:��Ƥ�ր�{� ��)�T�[��^G0��$��e�TY�#f��p0ZV��dXOp�T�9��@H7�R)�F+s�u���I)@�����r�
$�tMH:�z��mKx��ž�K@�p�D�G�%���ʩ�%]C��T�
ǲ�Gs�Q6+SN�����~*���L���p�8w�9iwRA#�5f��	%�AX���K�uRKK�uk3if=�Fa���K��*\U��y��#2���"�'����&�q4�xMl�i���'~D�T���@+G�$ͬ'������ ���B�%�ZU8|,ܣ%ͬ'�/����;�m��>�"���N���a�dA�t����,U�YUX�ι�:�^��#��0�	`��FA�֕�0�j�:~(+L	��CU�q	Q��u�Dq,����p���?CGQ�h������?�>�����=PH�?C�_�?�*L���ʩE��;�:��*J���+58��Iޖ��	�LC�d/n6�FC��� \��_1�?�$U��N)"�(�4����@���#&��I]�)U�6�2�)p
P{سդ�������z��� ��
�C����{*qR�JM1�T�� �42�U�hB�TJ*t��b5,���h;0�\��Z�F���*p�Z�!�:�t�jx		,��a�`�FT`)��| �#$9bFhf���Q�ë�R��%ͬ'$ia9Eq˒$�TFp\W��a�_G�,Q��$�#�Ru怈�HS5�@)���76�R�Zҹ 2�,�R:J����4��pE���$"��(���p�_G���r��>��P����j�PX��zB�n�w��0#�8y���(�؎$�'�0��C
cB�"�R�iA3R�z�0	�o� $CZ�f̠�p�v�u�!p}�5�#݃[� �Z(|���	x�a�����G��j ,*J�d1����%!�B,a9�8�]E钬!Be��'&���2� h�LI�gD`E��Q����.8 9�([����
�Ԡ�O"e*O%� ��d:EG��e:PFX�i�s�a
���X!�F$�.}0�P�9e,��c}G�U!(kd�FƁ�C&������ܭ�#�i��)�%�j���QĎ��8 ��A�=9X�/ WS���wD<Eg9X�?	��=�ȭ�;

� ,���{���P �K��x�@*�@� Dq��<+֋l�>Y�R�g�C���	r�W �b���A`��SN���D૘+��()���@�vd)*�������� ��)���BN<YuT�Рd�Ry��Dq�jd8��)2��(J9��*3*�0#I�p�BW�,�(���)�T�j2�3G�tQ ��W��(�G,U��bV!����?C �A"�/�-wE�k�b��d�qF p�d�>0� 5����%�*V(��F�RR�wK�;�O��g� "wnX4�T��R��1+���[0��+#sQ��+p���W�@(�"ׁsd��Y�G&+��x�(@ #C^N³!X��
�W��3"��yXE�3tP��U��)����������TE���U%�R)�g�	�����
�е��=�T ,�ܣL��(��q��5 aԹGC�F���pl�{,:
�r�F�s:P�I�-�J������Pmi8a8��Sa���f%=�bIU��gR���TH�>����mZ�6��"���'��DO^�[���"�g�[����� ��(q�Q�3
v�%��(��:��eU�b`���� 	E>��C��YVG.z"�d 䒪3���u�3����w�(���Ѯ~(]-����YVK.zr��T�#+�����jmy�񫥴�CH)ὔs͚`z%+-'�@��`(�%���%�	;��e��ؓ���M�@�=m��=Y�(4�� �1�p�䝡�����KL$J�����մ(u^2@��)�T���2r`K���fN�3.d;��\�I:~$=��@�{�~��*�5z��t�S�V��9�jڧ.q�q���s��"�	U6��eSY���}�eS��)�f�)0�iKzFϔR�I �`��J�+S���@ rZ6�D�ŠU~8��L#��� -���/!o�ی��-[Pi�ϴq��2�Ig��D\���j�yY��y ���%=#A���i��Ǩ"CePڧ,�q�������T3��%
�SOU�5�& ����kAu*�Жt���U���dÆd��	dwH�H��Z=�Z�QIy*�Q0�&+���%^3���q�yBR��w*qpNz�KӘ��`S���K2��Pt��A�����OQ�_S�q�z�(iNV�M�$&H	��1
WlDO	� ��L�Qqr�Ty
��H���cJ��D�7��(�J�¸K�0�0�
=Ed�?'���4��\������`t�L%(9�qZ˭��P�3���� �!����U�'�g��g��=�}�f�P���L�H�EO[�f�����J�r���0�(sy�@���Y�t<�aj�9EV�

M��)���r=YfiNF�G�A�c��KI���I����U�HV��q�Tw�u�J'WyOn4��(K�cOzPĀ%H��H�)a��\�,���B֨W��j��J
o���Y���+�g�łzl��i�S�`���p�����e��}Ҝ��g�'��	�h
���.
�V�;r�p�6��fȊ���,3��	�
���~��C����2+�QT��/zR%�S>'Ҹ~H�����V ��* ����J	�J^�o�O���(��;�×t�R��ۢ'E�T@[2*S�(�I�"�0���#f�̸���P>MZ=DOU�3n�����:=Z�甔��2?�Isfy��V���<�8z�{R�R����K�?�ׄ��ZP}Or 1:F��q�TR��cq����A*0��W�e`��SGeR5��%�z䚹�^=�.iĞP�Y�F��SN�9�O�}~ڛ }̃7K]D�H}��J���(!��P�	 ń�"]D"l�dIt��Đg�(Rq�Q\d�V�ʒ�BfX[
���1����)\�t�����vȅQ.H�o�,�Ӕ��� ���'J�����)[�
MȨX.�#(�ڼgF�L�9�x��=�|�t=��BBz�������&�bR���a��F��q��PyM
�i��!�	I��F����pʤ���<O=	�iQr�q�����N(���)�)���Y&�
27�dqѮB7?���%C���
۳����ڭ�O�[��Mb�rÕMVm�n�y��Ӽ��c�y�u�yfF�~�mD�Ȫ��]:���EP� ���!������&z�Dw�4E�j�������.�=�o���Cs��1���s�.l�6��3�r�VYrIR�\�����$��uH����!��-�G:^�g\DR���ݓWJ:^M7��+i�Ƚ礥��@�x���8�Z�*����ע��b6�K��缔���$2c�tňx��G{�UѩOZ�	��2�-����Ll�HCT�=�����jEh1:��N�|T��2�EhE`t��������9�@��9^ZB��rFO�s[�/�uG��J@�@��Μ��;��?1��N=���%u��RbǫSzt�Zm�]x+��At����n��A� �����,�W�7;���D�I��'qX��E��}+��n
�:W#�V�zU~��x��|H�HԎ�~rAѵM/�@��٬���Đo�n�1�I�9?��x^�$�Z�6�df�r��B�疛�k�I�
z��0������9�L�d<�D��Gb�\�	"o58='��|7�e���,#_$] �����ߦ�3"�d�9��7$��V�$�~�5Г%��*52�Y�u�6�p����,_B� ���U�nЄn��x�Q䭈�~��":Jߍ*z9�SIתa�<�$��|~!��f�i�Pf<)����s��]�kuY�$N%t�����Bb�0y�I-�9�)�r^�?^�V���Ҧ*��X.3�^��`��ZA�����r�_�s��z�Z��yu~������a�s]�ru��_A�xA7a�v�㕩7H�D~�#'�)4]��ym�g��iH�Ck��Y�n2o��o��S(RɜW��H|84�TOB�r��(Z�V#�
$g~�ty]z^�_�r��MV� 	�)��&�F�DM�9'�nN�y�5�\!�N�<
��<	��K* 3HV&��|Λ�f�ji	��6���r�Z%z�@ʠ%�J���7����I
���`o�\+�_�� �K����V1(�w��/�$�c��"ZAx�J2+F��+ϋ�٠.ጵ��S9�k=/9k�j�)�u� (�t�d^��N&2?B�+���
}��a��;F:Mu���v�c�tN�:��PQ&���E� �˱��@������q/�\x���>P+saϓ�z�D��܏�è�U3��PH��IN�]�[\�g��=L��K�)q��0�g�,�"��|	�X�j��_I����\�X�\+�i�z�5{O 2�^�"��­	�2V��~��� �e�_:�˯��7�y�,d�ݵ��D��e�C���r�*@�6tC����C9�*0DAfE�������'����ޠ�{2]|��I�HH��
�L���{��/�� p Y�ܤ�j�N!�d�y��t��n2��0L���u [ɘ�![|΂yO����������0Z"���D��x��0�W��đ����0p�և[�ڛ4'o�<bfl���OhE��yC�@��Z�'��1�GC�8
��{.FW��-0�7�HN�7��Uy_�#��Ⱦ�C:������EuӬ yȬ8��a8D�'��&�V�}��d�0}7�9��1�#	���p~ǰ�=o�a�՟0���1CF��/���{�2{�~܈ahZ�Ρ�2�Z��1��7&�T|���6�WO��er�Y<���_ʲ0��>BrJB��"��xx���ӄ���[`(��a
S!i���+)��H�׳�a���%G���$6ă�D�)Y�D��8A�q#��p�ޭ�L�ԑ���[`��F�{؁��WD�i$�QyI�g�y��g>nR&�]7�����Na96+��n=o�0X:��v�]<� 恷�0Xm�r��y3�yC��T�%|�IY�1t�� �t�6�,b��=�a��>��F�\[�#$��I��ﱧ�BR�UP���h���-0��2��T��c1��[r�S�1kU1�i��R��I���1}އ$��U�5���ɽS �¹�"�z#����,���eIoC"b����Z:pR���E#$���J��] x�*"��y=�T������[`,'�E�	gA7e3�[`,�ER#汧�F�'D �O�;�֟E�0��4��U����ED�� w�n\i)�-0]m�NL�B��)��F��X��_*��AF#�_xCY�&z��-0�>�f�e����GɈa����̼��TH��AF��2���T�j_ޗȈa$2'�}���|��g2b$����&�t����0HWT*�$���1��a\��x�g�"#������0U���x��H�UэPYNbX��2b�n�R�Rg���0�"������K
�y�)�O�%9J����YDC�\�NC7�9D#	q�@j���F��
�xT��XЇ�a��yX$\E8!����1"w�- m�:�ce1��Oɛ@Zx�9��FRu1LL���I�fàՆq�����~܈a�¸D���G����d�0hաbZ�:ݤ�k��R�nP�2�𵷋�a0��A Ï(�㐊FR���`��i�3�[`��S���5ؼJ�x����JB��`��U�0��/sOʀ�1�J��-0ZC�H���С�i=o�a��m`���%�>��������-�'��W�u(�[`�����w�i�k
*bŘ�ABk��MK_�P�(�Wo�
*�}*=��511}ZW�����*b�L�+�����n��T�0���+}���	0��uZ1�E�U�;���>`�y�(�{�!z݁��>�Q�(�[�ިXx����1���?�ʐK��k�y�`AA� |�Qt���Y�0��3�a�*t=bEwȳ� |ȧ:��Q�F�9}(�=F�1�k}~���xo�ȭx�F�3�!X��Ǫ�a�e!��A�@�P�V� �����҆ڕ��ޗ�A�p��V|mEG�+}D媠}p+��a���ح�礦˙��FY�@א��R��ۦ���D�=�?71��k�{���)�C�atV$m��R+��:b
�,�&�&���ǩ:bڭwx��T���WG�黩�s�9i����a�d�^B^�C�<>��h�SAPT��"���k�x���`��l��?�À�{��X�Ky݉F#��O�#���5D�"|2K�T 9=�p��`
�Y<��O�Hn�`
��%@g��@執�a0��nE+���Iz^��FCS���B�J��a�
5��M~M��sވa0E𓚤Zu�Y:bLa}�Hw��,��5DC_�ࡄ�¹�}~�#�q�گ�(N����y7T3<���lz�c"���)'?�:���8d"�A�

Co�2C�R¸�Ak�{����5�bW�G��5T$	�E]��-�뺉�Z�Ã��89o�a���!�׀��͛�a�5���-OZ���Z=ޡ'����%��1�� a�n����/��a{5�C��X@Z_G4��W���W0o"���~oàU�:�!�/H�k�&bËg�=4T������pև(�:i"�!��^ʇ�� �L�0`Pa�z� ^7à5�>�X�¸:�L�0��Z�;��ri��Ɛ����4�<7À�P�pB*?,�[`����-��GHz��kL&b��3���6X<��g&b�{Á��C��x�D�PP!'�q5�k�&b0dv�CӰc��#�1�e� ��]<\��+11��Z!���b#o�a� ���z�J2��[`C�)�Y��z��o�0�M�c f�&�k��+ۈa,}Q^�fC}�����1P�!��.Z��f=o�a�V�<�����]�����{Ɲ3�!7����E1��a�p��`0�c�����Bɹ��l�0"!B
̛��/����0����o����(��2�����xa	��q��_o�0��*�W�����<o�a,U�Āj^�ع�b#���)��R�y%���җn�7@��Oڈa0��
2@*��5R1��uK��wA��<o�a�G%����K�d��-b�3��ᰃ�4�x�-0����n:⃔<&���%�;pt�͇qrPao�XCߐ�I�t֕�r��Xz�x���[��Iϲ��w�Z,]��֥��Rw�$�_�Q���d   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    R  �    ~  ��    x       ASCII   Screenshot�lK  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1662</exif:PixelYDimension>
         <exif:PixelXDimension>338</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
���%  ��IDATx����b+Kn$����r���f�����f�i�m��,�(���@ �)��3�ͦ�D��2#�@ h�駹,�y���Ҷ��N�T��/�0���Q^���g]���yL�O���g��>�~��?_z����~��{�z�=�vl���/����>&��]����c�g��K��>��)8�+��ֵ���?ȱ8�y�����t]��+o^녟����k@�;=�<�{UV���Q~�Uf�)�;���������b��8w1浭��k�\������1��F�n��ֳ�ɦI�D/��+��4�a��M����M�,��g꺱��up|�5~�{�9��ƞ������>.k�k�;/�x�n�-ϝ�<��a�	��z./�I���k������^>�/�k'��/��<!.0��%`�.8��|�ȟ]�g)/���V }�m\�W^����<���B�nB�
���(�~˵�X�\�i�r��m�g{�׮�*�n��"Hl�s�z���-� Pci�3�$���P��j�Y������`��Y�� �uRl��
��s^���k[}����4�5��s^���|H�����Y��=��'?7{���WS���1��%��ǩ��nD�{��n�=ޫ�x��!��s�����L{yPy����ܗ�lUf��q@[v�i�޴*��S�vv8�oi��_�j��K ß����(����d�~˹��(�z��1�d˖�k��h�5?����//h�����! �8����R�;���ႁR�K� ?������G
58m��B�Z��n�<�	���j��MWe�8�U)�R��4,L��?��)��)����T��� N�$��(���ܸ��
���p����}�����s�+����m#���i�Z8[���D�lw������{ �ֲ����"'@^[d�,�#���^;޷��k�{���k�/���6�y�<.�ւ�З�g{��w�{C|&���u��o��ۿ���?������o|ӞgS3H����c�'��� �`F���Y7&|��X��
H7�NVo�q~��<[ V�Tޜ,��z�d85_߹�r�s/�c��1	��^u�Y��έ�iD5~|������aT+y��O�ʺ���f�ǹh��GL�Ȧ�2�j��\^ݨ�����|۵���i���T��=�k�齯��kǺd�_�K���l7��wm-�kV������6�|���]������w�����8��rk�-0�vn�sE[S�ப�V�b\-��z��߬�K�Z��>�=j=�����_�O�Q�����p��{yi#�s�����5��%���r�Sv�l��i�s���n���X�u����j�v�a���	Hi�ft��K q�Z�7%>�X��ސ��e��}\������?_z���fs�����=�@4.s�y�f�����js�ڶ�o������Эq�;�kc~�ҹ��o���S��֓p{+�.[�d[�������,�:,Q���9ߗ �K`�?%9=��6m�eե���[���2��XK�{N�w	L�g�ݗ�+(��qG�� �k�*�V�z}�k_�Z��Ā����D�@ʓ"�:�����۽�1�����*͏k`�?�__{ϥ_��㵽�;��ݯ=�Yp2��+V������U��k鋅��V������g��va_s���[���}�r���}S �_Ӽ�0s�>����`�ãi�E[5@ҕU��LJ�!��9^WWB,؊!�J��$�t\��	�?��.�g�_j�����Vhy����w�z�cE�����ϥ�9N5�.���Zq\~�	ەh�r<�N���<??�?������j�� ��Y�����_]x�I�M���Z�[�Nke9]�ޮ����]�?�o�&9�,�8�8��{/}�{�_�}�Vvv��h��r׬.\>�}k!^;��{��9,@*`*^SD�4P��"Ȗ���z��=��ɭ��&��ʏY� j`����Z�[�����P���p��5���⸎��7�n����Rz]�ȑ()9T}q�/?�ŵM�T��۵�aU�Vr�ĭ���o�z�~H�<�	,�e��+@���ɟ��ׯ�Ŀ�z#z7��U�eS>,sp�[��53>_߻5���o�����߽���O����um���)7�-E���^s��0�f�^�k\[>��Z�Ǿt< �C����kns�3S���]�K_h�o�Q� bx`�������
8���K�~e����k���������3�%���#t�M��ſ����Ks0oa�V0��B3
 ������?|/���hQ|�߾�ͫ�h\�5���M��M�$-O�(�_�|)����<��wy��ϟ?�u����o�1�y�d�f{[ �fM��[^7/���������-��g����}�s�&l������|	���T����9]Q��D%]�����߷�l�� U�iT��`�}�/��z�ƾ�t���J~��wN���[��Lpk�*p���פOЅR� o��c�y.�7�YH��+�R�V��D�=��:���� 8��������[����������bm�������f�P�������{&����i��N���@1���|������O�������/����xL���% �����e����v�̟�<�/��[�,�j}~�g.�|�k���5k��ud�k�.�5������\�k�5�c���cѵ��5�f���Tt�/9�)}��
��k}������I���3(��j<m#H(r�Z��h�E:��� +�\W�A28��]���փ�Au����9�6����[�
��������A@���S9,�#����l�jL߻��6�µ�7�W��'L�.;\wX��<� 
`�k����(�v�ǀ�[`�.���|�^r3.Y�|�%���?�|�f�~˱��sڂҵ�o��K����K����t�����k�@�;[K��wl5�[�즶l"��,hM�8�9Rr��A�O��r���c�f�͓Y]�����9 �C���[. �KPŵ�v��7��V� �H�8��0���1���XO���vӸ���Y���Ҹĸ`�������lN?~��\��sMA}����X?,�mr�����=$x��Iw��' V(�F %��g^(/&�y������3@�w��@���U��G����k��%0�f�^����~.�k����/�_�^�����2���ZxϷA�Ks�7�ɬ�������۱��K�!;���1�L�4�8�2�b]?�%0EVT���V�1S�U�i,���(�L5G^%jIgQ�֖}���΁����<W��(O� S���\�E���>N���_�"�����W-�YzNr}�l�%uu�E�oR� r�t��{��xps�h��.X�E]r��m���3~�[�@���\��luw�k����ϳ�a[+����e����.Y��6�Kחݳ��l��K�|�\��˟����f�G�:�Ų-�Cω��I���E��<�܀^�����q�	Ƹw�.��s�k JnځT�$���V�<�H3-�� ;��W�w�1QtH��Z�d����F@
�	��p���*��_�B����Q�����v��`��	���^�e{�(,�X�kq�\Z#�<��i��Vf��&���Z0�I. ���������w�iN�j!x1h��H�AVYH�5�E�W!ݴ1�y4�^}�U��)"����rIULT'�� �9i+�]-�q���Ť��}��|��)i��-������@�q��Q�"���@I���>��ܶ��������ww�]�A^"c6�[�q�����"���:��"o܌�F�ە5��3����'rs�3�<��%���(�n�%�F]�xv]XB�-���� �tVeV+�9��t�_ɽ.UTh��'���yۦ�u1����Q��K��R4��߻�b>v��J�s��R9`QzTl#�Q�}�s�d>��+׬Z�h�~�]O���HYxD�⨹���0�vlU)�q}W�[�ꅠj�s��r.S���㳸��>�ݻ����$� V���-��$�;�QO'n{6ĵOT�]3D�,����iA�_����?���_��%2R)��^�L�����տsʕ�P��/^�t��I���r�粓ส8�g͚��D��A`o	>Zk���B%�3G�H�����xE$.�m\,����q2�.���;�Z|X�zUD6�:�:�����\^�@��S�}/;/������tNހ.�t�G\�|�`��r���r�q����=Z�L���x��2,ݻUw6�1�]��l�J�4q&�%DW��@�/7鵋��%F���B�a�X4���{Q�h�6_p�8�����=�\����3q�x�"=с��5�+xb�XH�gb��J4������&��f@������9�x-�_ �����'z�Ј��p�;1d��s���/<q휏s�N<��l��x��������������OY�쨁Ù�����7�r4
�՟̒�*�֪]�cȾd@�	�믿���������?�ub�,`a04��ˢu�{^�"��dd�_&[?�F��P��@�������V|=,��U���t�67��|��y�Eۗ�2��ʀsX�mc;�����gV��1&&wV��cnn���]������J�����p����\�h�X�&��.����bjOgD&o����r^8���Q@��'ۜ��agr��r\��g�P�ƣ���SY�B��p+����mX5��,��QT����y(��Ţ˙sZ�M%,��\�ae��Ƚ:��D�X�@��u�ߍW������
u�U����\��w�H�7-&��������Եt�k�b#S���5��#�)�4ʆEQ���(*B�����ƌ�ȓW���o<�5�������h��6q�
�
��F�2.�����'�F9����
N���{��y�0?���8��~o��A�Ԯ�V3�k�|���N��_�o�k8 �+����H��E:{=l(��)�� �H.�T�Z��A ��ڐ\ x��鯿�Z�d���.�!7S&=n�IM��tu>����d֠�v�q�`��ЬĐ��ݻ������?���u�1i�]'v��w��n�I ����K@�/׵���r�K>'�N8̱=���q}�D����r��)�NE&%\��[ )&�k-�EKւPm�ܲ��j=ʎ�'��\����T�`�y�����ή|��w�qM��NT���R�\�2隶�c�~<?�eAcǵ �︻�),��;��[���C�V�.tq\Xj1	O��H��Z��4 j.�i��ԂýQ<x9f�,�Zh��$D*��`��[�7�Oq�Zʹэ�	�?,dl0��5}�t�X3�6{ә�8�}�^��A
�XE��s�}�W��a�Yօ�����4W2Ns��}�!�A �[�Ê"8�U��w;y���{\�����9�fe Tc9)k<�6�c���e�vK4h����*�B��������������1�$�f�	zN���`��/�8�1��fhM�em�:==�el';�nj�<k�-6�v��*7\���' ���x����_@�m�5 ��?/�ݾ�	�Xz���2�9����Ų�vbk)�_IA�	����c�����0 ���Í�V&�y���E�3�(x*���\�-�p7����,��I.���ݸ�������r	d�zvz�.x�w��	��q�������]�ܟ�T�!u�.��t��sc̰h�Uf�HĶRwJt�8�Y>����y�Bw�y9�mo��.s���nnj����:X%s�0�]���F�C/��kx�t�ټ�'��~T��*�� �eRY�zϭ�W�{��4��{d_��{j
�1&������\��,�N��Y��܃e�/ks$s���z��4���� ���NU��G�	�t����|1�a����ʼ��}	>3|+��5fh���)�0�u��ū p�:��y\�r1ޚ/��*��Dj󎻾[6�[�4�����˸��&���.[�!�9i�+���7ޡ��>Λ@z&�~�,�������ٹ;l�.�|���I
Z��n7L..���ﰨ0��� �#��d|)^��;n ]*LG¹i��,�O �e2"�@�V3���l�o�-_�.���pN�Tª�
�T�����Od.��Y�j�+ ~]6'<�g�Q���_��X�ߗ�~E�د��u!������2x>�_����<?;�M�O-�
��/^ �Y�j��g��C8_|?����tX��YqP3J��8W���M�Z<�i0~\i	 ����<qH	���])�+[�'x6���GKQ��,�έ�v�W��R��)f=�}��bƼ�XBM}�J�:��;c�bQ�{���㒫��������X���|��B������&�� oB��s�w����ߋ���7�W7u���Ÿ�g ��`G�VL�e�T����ͪ��w�2H�vIj�����h-͋�1���.@{g�����)f���'�y�c�(Ć�sU֤]O��\�Jw������c�� �".�^n��;e�H�h�%u��0H�X���.��eq���-���?L<�@�w7�X�}�w�Ggّ73K؂(�5a�
w�E�+��d����.��k�b 7��������f�Ҭ�����(���f�H!4l_4ݪ0���p��Z��w���������o2qZ��1I�;��^8��U)��1�O�X��S�@1�!�%J��ˤÄS>\-/	&}��8��i��y���� VX܍�	�; އs�Jٰ����+?����+X���0/H�)�����W����{�y� �r�O��86��x����������<����\	�3fH�h�������|^Y� ܤ�(��ȇ��#��ViL`0O <}���픑m�/=@ ��oI��u�t���4������p�ܴ��R i�<�	�"�~XE�{:٘H[�"��tTSb��>W���Ov}��'Z��8u�Z�輺�?���J��-C��zh4a͐�ˢ�l�2'�f���D?�{���_S���$��w���VwQ��W%E �j�H�뱝ޅ�EwSXn��oL(��N&���4��l���jQ����yH
�� �ާJvsq�d�܈E2��]�'��؝l�0�p��ss?��t*!�k 5��1+B΄��8l��y��˧f� ƞ�w������P �Nґ��t�צ�h���PЍ�@똠{��7��M:��P�샎�͝���"R�ND$Q[s[=�t�Kc�, �QW?b#� �	��̡��ks��J���������X r�đD������V�S�餯M�@��2�m�K��z�R�Dc�6�D������D�ʊs �5��\<��븩wb�1��ʔ86O��-��w�۝ݍ��k�!��[!�y�@�Ojk5q��x ���U���Y�,\@����NoQ�������Q��Z�x�4w
��rW|�"�������"U�Ckx]�E� ����_�R>�~��@���(�0wZ��p~P�B�9�p�����?�M�HA-r�EQYvS���%��K�r^X�p�>��I�ߋ���I:$8&��fh�������&��^�9��WKe9�r�ɸ��� ��N�Q�*��5�a���ir��%�`L9Nuc���z��|j�=sqޝV�0�Mp���H�1��-�b7kʠϢ���Y�lŮ��&�N�,!\�Ԙ0kJ^��n�s���s��@�p}#z7*�!��W@j�'�Ż��&bR:��+7V���`� �2�b ��� p� ��R����\e��J�R�pKq�l¤�X� p�V�%�v��~ۤ����u�z>0T��`o<�h u���4���H�����eó]����A��ė�n�77E�[��l�٢�����q�w:���%.?aA�E�I�T4�J4�	|�#��6+��j�u� 1��]'\�G\�&�� ���Y8IR	ʙ��2 ��7}X\W�Q�����~L�]�a��G$�Tk`����hgsC�I����*�����{��r���e!VP-�Mڗ�Ȣ��y�I��E�� �y><(?��a��4�9�ɤ����M<4Тꁮ]��l�,� ��W����Veeҥɬ�N�Wr����e]��ﵕ2@G9���c�,�we����ǯ��È�9<9�A�-�&)׃~�<W"|��8x	�ڂ$ͨ���N`�;?('~R����o��:��jZ����ѧi�8P�#��g�;}	��Nܵ�C�_%�P����7i���k��=��\�5���Oi�5)H��g�����5jr���Xy��,�l�V>�z�:�2�h��B���f�7����Z�;���v�ɢ���EJ^�r�;#�%�4���g&��]�8X�@�4�K��3J��߼VZ���4I�~c�s���� ��]����ν�t�8(�bz6�J�gJ���ANº�>BS�6��dt�ܢ�~����g���4��$�d4��>�7��Xu%����<M��u�����vu�޲X�%o��ZW$a��X�hx���m�7>C�oZi�l(8�<�Ώ��,�#�nl8bɎ�G�u�v6����GS���r�B�D���+Ξ����u�(t�A��g�<����m����p�SA�Q�LK:W��%)1�j�{Hml��:�je�ǖY1�"}����ϕ��=�W���u�q�5"w@Ć'�lq�������r�Gq�(�厫)��v8h:'O�|�=̚�����ãg#�f��%&�,��)R�XuG���s�ӈI��8Bja=�ƀ����>�DA�G�9�S!]bn~%�3�טe;�({�E{6KB9���D��e��� � �����Ь"U��U�����&���h�Hnj�,��63+؛��(]�n��F����>XY��,��`)ugy��V�����5�4��yn�腄��C�D��4�Y1��3N.��$P��k�ܯ�=X�'w���u��믿-��,���1"��U�a<�s6�X��{��� #�2 m�����Y����p^�� 7
�s���x|f�0S�*�nE�)��poSp��*7{��y���{�(9�9��֍S���h�u�p=�-2,�T3�|��W�)Ċ�f�Lĺ?{���ʴ����;�M����&y*���#���EJ0}#j�rP��/��E&ԕ���s��Ee)��f=..�ނK��� S�KD�6�1uy��}��ew]���&@�I�dL�[\��;�t%��I,5F�w��gia!Φ�"�"Év/��4��d��2^s��E �IWn�gW�ke�G�7)6�tA���Z������}����(�=��g#��L�o�{#V=lt�I@|�0�W>:8�
?�����bs.80Xb�E�u,)���ҹ��A��{s
�5^w����g�\��o|>0�R�����-WK�����RF�����{Cr��7t��.o�s핣5�^@ײ���������s�^��H��1D T�#2����i���G�}]�s��B8l��v���=׬�,*5��JhQ+A�Z���v>���j��4%��ܑ�c^��5 \��i,BO��+źtci��w��Bg�5�@�A��n��ViH��{�ʟ5�?V���X@��ʭ�j���b}q0}�"U�xp��w�Y,mT���(���WΛc�&��E:��"w��Y@ԄԚF��p*���T��2A�1 �U<,�2ɊEtլHD�L�T�s��'+%*X`��������H�ĸ�HI	��]F��F��V�2���`I����Y�Q-��@01q�,RKR1qݪ�8�4\B���3��RY�p����D��o(����΂߳-������΢���n2g�:)ťX�)�<؂�v8�BaU t��7�)�j�ߙT�\�2�R����?��P�v�@?K"�U0�ň��i���;���H{I�T�F�饸vl����;d<�77cX�C�s颟����W�d�$b����hWXM�����P�:���)�F�>�j���N�A������3��h������z[ߐB�kB�3�S9�弻z5��G��'�c
dAUּ��0֞:��d&�nm��`2�u�tm��M�����7���|C&^gS�N����.�*������_?���V3o��o��T �D��CuTy���J�;���$�fՈKb�[�ƩК��s!�[dTS���x4�B'����h!��u!����K��+~G� d�$t����W+iΓ�	,sG�=E��T��VC�����g�	PGը�V�	�6��F���k�T����,,)�;�Ɠ�.Fd}��-F��XdC�J���R�=6�\�LK���Xq\�I�;C���E��z�M���g��v�`�Y2�&qh����j�����`��s@j��N��R*�u�NI��#��0J��V��7n�3Uz�l ��,�-ad������Vb�^e�W��mSWHH�A'�@�.0=�X$F���%QX�7��,.?Y��˭���4EJ��uT2�[\�r��7<2G���Ez	L]G���)\=�|	�t��b�Q�"KK�E��Rɓ�Q�!���E�o�trkV��a�ź,�nq���pm$U�`�MѸU�b ��Ȃ���H[*���!�q���"G�v��q/V�B ԕ�|'�,�K8����T�F�����������82����(�H��:0p��9�F�;<�1a��/��Z�`�z$9D^�2y���?	� ��F�Ct��]s9\�\���Wǆ��@��WV��v�B���Ϝ\�	��@$g�c��3��͛��T�v�sg�cP�E�=��<{K/1XUZ"n�+W�o;�!Q#g���*/��w���w,�䆍{�h�ws��\�D�l |�9X����1���XO�҈�M��97�т�b�@\�����h�'\dۄqg +X�4�ߎ�Ȣb��H��t���*�p���{4��V���ݔ�u��ؕ��e^!�l��KV��1�?��o(�,n��0�+�!��	�­�<��5�0x�L�^ ���}��u�7�������s�ZN�P��W�|�Ny
�a)��u҉X�@A�IGwe3Hc���\���,�M��f�9\�b��@�,���ieV��&f��r�9F7[P�rB-������W��|�ʻ�;�wf�<���r����.���ad>"���2�(��)M�8�Jk�剎�^N�iLo|��]�|�jY������\�4�0��4�Ҽ�^u�X49�7��������)�����fM��ߤ�TH7���h��Tk�=6�O=��Ѭؓ���=�N2�\��9���~���d�q0MY ����2y��B��lƣy6)�P����Ò$�B+��Xs��qTl��\��-GJ�"k��k��A(肷d�#{%t����{�#N����D
��kuR�à!��Q��Ē^�Js@���I������Ѓ��o+p�Bxp	U2�9I�*��e}`�a���R
xYt�TaM�X,�&?�v��12L	P�2��-]�:�QW�N=X�yN��WR�B�Yt����3�i�3�Xr���O9'�v�)G�׋d��Z��ӓ
/Ƣ����̽�H}�ua%�S��[���M eAV�R7y(ůW�?�hI��qZQ:��Y��`Jc%�%��@��݈��q�S-QKv��&����F��/�-�_[�杏/�W�~ P�����\��3�r���%;�[
�,���K l�C�u�i�b1gw�=[�>�{I�U\ŢT阧�I`ρg���Uҧ�P-6"���[]#Q�F���h`��1�RH�[��i���p��m�&� �3��<��{���:�u���<�+#<=�d���~ٵ_�O6Xu����lN�7լ����Eц�%C�v+�>8]�� $f�<�kf`��뗯�9F�]�ٶ �)%�
��U֊�u�n^G��J�U>�&�t$����N�>���8cӤ�!� c�͗A��GP�)[1�l1M�ù`q�w>)2���/,D�d>�$��jVR*L#��U$֤D��Ľ�h����^����wi�p�yNV�lE/z�=,>�G�Y	���|@c���be=y��3��{\/�@j�&��l��>R�Qi�t`����l!�)rO�{�fM��3�MJ	"�Q��m�iu�3����5hG�ȍj��J��w���-竅N膻++�r�EPh��C�`̯�A�Μ�`R6S�U,A�Ӻ��������
ߘR��u���)m�e��K�u��Tk��������v��^��d�Egu���r��g�1Z|��-l�W��Mמ(Xj��쓆@jBw�529NP��5���u(��M�b'ǂg��87t�1PR@bpb��+���=V��o�0�Vid��pcΟ�,@�,��dգ�:D��\�]�.Ό��k�{g��8v���1��d�E�e!-�딲U�2�H����'Y��~PW�$ORXD���� �[Oo�9��]��6�k��q�|�&�ʹ�4Zh��0o�	u���(0��)o���u��;6Nl�qM���� @o�l�p�nM�U.�@��1Ƈa�Q����Qa}��[��e�H���y#c�>xU�W8wՌ>ʆF��vjQa��z=�\�['d���jU����$t˜[*үM��)�ԅf>����cLG-�"��Nl�7M�T��s��^z��I�N����aD�u�InJ�d�<.+{�n����ϊI���d��ΛrW��e%�z����8��A�z�ld�H��N�:�6"��8[a�~�1K�k��h����U~��]W=
��!���]��wM�S'Wg�`�9u���z�(�h��^um��8gr~¶ksT,�k.�˷�h��;���i��*7��c�B]�H�+V������do�z)`k�uUu�1� �� �ǣ�8�Jj���"
��x�.�)�A�J��<�Kmջ��?�Y�CZy�< �?� �B����	�zGL�z��廏ߋ����</�S1`�nS�o&Q�1_;M�|R��5fa!Dq�,JN��<y��}�(�w�ڒ�� C����|�.k���cI@z0Z��Q^k�3�$�ۃ��a6y7u�%��4�FU��,�X�A���"�4C*��+W�T�v%�,RD�ihy�H~�z��Z������r�L�	
��U�ȸι_�`�Hg�71��zQG��~5�ֻ����8^D]7.�e��јt�[�.� �'.�I�-���{���:����6.Ց� bGС6m��b-g��)���ּl��PLN����b�ձ�����=���E�^FUE'��l-Oȥ��dO�擻kl`G+OK�=�UK��2zͥnl���4�����h��ڂۉM��A�� 0)����`���Ǧ[E���q%n�zL 6h�s��G�\:��;1���3���𜬯 T�<[:S �|Z+l�!�c7�S��hp�qa�EZ�
ƵG�w{&�d��C�ylNz'V5+E�j��pݣQM�)�qI`��1��#jo\*-��5� Qjk���i%#X�ˁQlL�9-��Ѳ���jG5ـ�h��$F��^��3�7*R��jgJ�� m���޺|̰`�8��dԉNv�0�v�e�?��� �,��}+#�+`����+�|��3���[�GѺ��/J@�&-L~K�QHY@E�"�D�.����e)3N��TR��,:���oZ�q8x�s�����I-��zq���4��uU����$y�*��-C�u+%�nk��d p��<�� 0k��cD?������H=X݁[[�fF~�Q ��9ϱhzM& hb`y�K�Y���+/Ӧr���Q�jj5.'����b�aQLN���,���lW�|:z�F"݁{�1
%���$�ι\ݤ"[k��&�Qm��hiC�0���$dHu�G��3M)+ҷ~�O�*�L�A+6�76�T�rȰ48vS�[�bxo���

��k���4%K�ܻ��͔�A�{��=^ǵ�������WY9H|v��=ߝک�"�~)֗5mU���oi�j����d|z� �ƃI�Kو���3zpNL�Y��q��Z��˒%�h���!\��5UO��]H5�;}��En̓e�0XE7��(����q����P)q:8��ߛ[�L����Y>9w(E������ߍ��)�	���P���dV-?�yb_l	�,�,vw�DkYw��R�2���Q�1'O2z��}��t�GK	�Vt6���F&�&V�;4�Y
N/@�q�~�J���-uQH���;<@�Q�x�����W�`���]������������1S��mL��HaT�ܺy�g�$��8F��AwS���0�J=�1��2uS������,X�n��V��ƀ����
��b�bĸ��ܨlɖ�[�9�Eԟ-0f����-/����<aHV�g����q�(��Z�Z����r��
L�.�*ӱ/aP/��Y|G�H��=�B*ы�B�D(58�=*�$y�0$�<��W݄w����G�E le�f�h��9vF���:5�%yb���&I��f�>�&�����R��n>�%��S7��AK�ꝵ+p�xN�o��c�N���k��XA8w����P[-yGk˅ģ�:�Jkͭ���Vm�B���g��7�l1�YE?y!�;N�$������cX\���ꏻeUp���k��A��� ��nR�{�4γ��6� �s��xc�U���y�X�s��j]�ʶ�u��A�k�4�9s�+Yފ�� |�q)M�ͪ�ַ��Df��Z����A}�b����c�ƆŢ+���f]��RF�J�,2��f�'��FY������l���Y�ō1$j��0Ƣb�����^RF:f�S���U�Z�h$1+�����̳d�5��8��Tۚ���VH��Q��-0 N��d�W�@qk+�/���0t6���� �\{J8L#�.��Z9$�彰T�O�r7�VM?��a������2kA��/J��J�Kv�s	��{KM��� �1�Ѣ���/���՝a�5ъ���X����;=�E�e����X�|�.��qZ��� i�d�3H�*g&n�l�뽽���Ƥ�5	��I�{��0
�Un��L(�? ���8GX����w�z� ԭ14�U��c��/���&<(j�Gԛ�F��ei����2�E�95�7�T]h�)=˜N�(�\��������:
��y\vև*m���}�0�D��2>��Z�{���v(�(�B��EjD�`4���~�����[��� i�31ù�q�B����N��7� �;K)�x�q]U���p�YmI�NZ0�����z� �~jBWT�˼lB� �����`��:����gԞ�Y=�3�|.${t�W<���+ �&��nQ��ݬ�6n�r��ɕ;�B�q ��	����C&Z��n7{��%Z���,��[6��ƪ��zDo�H<>}Vyʤ��rJ����}^����k~�O�/3�0W�y�k��	ԭ@��Z O�#o-$����1�;�;kJDV��X�+�DZl�C�Zڤ�e�"+��à�.�g԰
>+Qy�q#�����h����x<�z�t����T�T�� �D�����_ʓ��x?�4{1,���RWUH�,��VJ�'%>�7��;knҥW~�%�� �ȝ5sd���<mEì.���f�^dk�{a��{���;��"	cd�	��A6.�@��U�vο�c L��e� ]��b;��,�<���Q��NXJc��n�	�Z��d�vֱ�Fj�A�0K��:����jӞ[л*N����M��r]�K �� �y���f=5���װ�eY/�c�����k�6|�\�U9)�l)tQU&�)�KV�v
e��f���Y�r�K0�)�����Z�z�H����D�/�������4S�m I�x ا�Hy��
g��eAU�]Ŋ�R��@��w���K��VO�����9�k� )�SJ��Z�J"��Y�T�7&����Bp��E�gY3��tk�QX��ts%G�ւ-�ъ~,��_�_��/�?��?�/?�R���ߗ�֪���{F[��sDe'�����|�/_�3�j�Q̀S�i��G�g̀(5no�zƀ��)�Am�`J��`��q/03Mn�)�]���{&�Yu�Sa�I�j�"�lC�tV�[�]��9l�W��3i֝|'�+t,@��֊_���l�2ԊSy��McL^��S��<��Ϫ��(L��ܛ[O����h.aOT�m��"JRL����lY�B�9;�2}��D3��Y��g�B���'��XmaT�!K:�.�f�f�.��
�L.L��z�|��^���~K�K7� ���
?X�6�#��h�.�H�l�f��P#(n�Is�5	 �`��T�B�;˂'���'�,�n��̈;��i�I�`N�W���fϓV��� .�7(wi���Vζ�J7��.��9��N�L�G@��v��㣧�>=j�nB �,�R��tc�10:�{s�q2le#R!���TV:��π�dӉ̩�6��-Zn�H�Rq��*=��
��|��]�kp}����Ze�U���q�+�Y܋�0��b)Rg`yb�b3Op!�נj�ɏL���%��0���8{��������%n=�nz����N1����֨�+"�>ͣ{�DşE�f�2�ڸ��.��ծ�����}^�D3ff����E�֤�������4�5c�.�Z��Kr�I^�<W����D�����Lg
�/n�8?���0xAj����U0z�Q�Hd�<.�xy�^*g#-���NNO�J=�Fϥ8����T�j���P��Z2��1d�
���/,N�F!�3�&n���#a!ª}�,.�`Z.�Si�ڒ[d��62��STC/v^��d֎���h����|�H٤���A����6�q��ĵ|����ճ���H91��j����¢��]V=װ&=e7)�;][G8��Ӑ:������ާ���1�T�l�,�ϙ�a��$6�\�����ؐ����C���*u�,n��_�^cl���`�֑Qd8.��֩��G�Q��9:3�^�he@:,ލ��d��9f��-�
d��r��O�0��&�4�7)�����t��ǟk�M�2��^c���Qi�:�*J�i���L�7��AUf��	=s���6.�4D3}`�ǀ˚X%0�W�_|��R��~�W�b�u�'w���]Z���lwf?��}�:��Mz���.P+óT�r����Uf�7-��ohU���цc��5Y�Lc�U�m��&�`���O�N�f������?�`����i
���M�q�B.���m,m��(�L�nj �a��:��Lw�^���dAS廿���g��o�����U�f y��/�$���%�j�U�u2|P��epP����#�f̖
L��,8�w��+ 5����J�����\48�O?�, 
.����HE��s��A"2*I�T״L}��!o�ns�@R�Dv�H��to���d-3��ʸ��M�.#�b��rՠ�@!t�I�Z��C��y]�y��B��x^�esր��M���~��8�Y�P�����`�E(O+���z�s��u4s�X��Y��	�x4�k����,�UZm��E8�h�ؔ�TК�u��Q$(@�4�nj�8��-���"�G�������0L�

���g���嶀�cN�7�~[�ԮZWB�P�)��t�q���lLr����Z��fK����8M�*��1�i��za�������W�v��u1z��N���0V�ųq����hG�c-Ց�~&�#um�:���S�@-�.�bF��8k����[?��借O��#���X�X�5��k�E�g���53�q,�=��,�Lk}+�ք��DjsX���d�)�!�{t�p�4d4�^X����Y�.ߩ5���>�N���T�a�W=�I����5�9��U���,KĜ��#�ߞ���.-�� ܨL?mr������Q���m+kI�k3S]
l���
��XV�{/	���ݟ�(wH��9콤|���xD�Z��\b��Qj��s�7@*��z0I�M_�~r)B�j�[U1h�iDfu=�v��Uu���b͕/~�e+����񇳻h�s���qe��(��A�c��t�f���'�8x�(�@F�%ɓF��J���8���I�����˄�F�(Y��e����X?���D���&s1���A�@�g��_j�f���Q2�f��ꃖ��&R��� �Cr�U�f]��z,`A�m��u��бӂ�8W\�ϰ���u�m�*^Z���tŕ�iV���D�ժ$q|��И��#�ުE�Z���'jJb��o`Ѿ{��GX�����
��8&b�Z���D~o[*�;كbO��O�R8&�[��ip��*�SA�\X%l�é�N�`CňeԅEF���I��#�yK�,�"�>A�@��>s�Z*����'(#�ͽO�i���։w!����pe�&�0ŕ`�>o+�8���<��aH�@V�d5�q/��-���+������9'�YM��k�(2�Ze+�$k�nb��53n�B��
Ms���`Br��1�T�}ZU�Е���6-�'E�z���R�(e�D�jn.�w���0儤���,׶5*}����h,�§VU���^R��`I���n���,X�kSb�B��,��RU��#��/�
�Q(���7�����\�����//� �K��%*4$��,����2�S+X��7����/���T"����I9�k?�6���!���߂��
LG��3K����H߿��)8�ުJ1���\*�X�u���A���-��l�Z�ٽ�\������%$��9W&sW���Qfy�d��*�j;/�Wl��g��/�57\׺ �I[����g�4Cm2�����I Q��䛼t���0̩ R�Z�&�?������+�UvΝG�c-g�U3�M��Ґu8q)L?��{����
A]U��$��ie�
��.|��2��V�@���w��5�
P���^p��1��߇�#�D1�s�QvlX2�|��m��!��i���FN�_�-���y#��Ux�Uޙ��\o�]����V��BP�����+����Q�:�dp-bLD'�闉���S�^h��*�ٜ��ֽjmյU��9�?J�S�pm:���dp��f�7wB�@�`�+
*cӑ�I� �	lN�e�V�ѽU[r��	���~,�BE -R���"�5�DG�������/�������
C�?G
l��Ŏ���,�y.�<v �M���V��'��E��J~s�}�r��vQ}�Zе�k���v{��3P�uD�i�jO'si�
_ZY�i�	�XU&�RU�V��k] ij�X�ww�N���;Z@�-�iE+ú�9�L�TË]�e�R����I:,`^WQx}^=W>�d}Lۙ�|e����W�?���s]�d���Y�\����u���j�P �Q�����o@h�������Ug<����m5�V���p��%4�&��}�}�r��Ҵ�OG+�i�����e�P	� 8,�&����&CK���y3��;y�ܓK_�-�f<r�V�{���#_��a�nY�8��"���I�b�,��%��~!�Xu�s� �ј�[S"!�8Ǖ:�Z�ɴd�R�O���=+Uͅ��p��R#ʂ.����F2\o�eWҞ�Q����nnҷ�f֒���M�"�Qu�D��*U���J$�?Y�G7����:q��E������1�w���&OLtP��F~�*�?�e��{�˵b!j��N���+����i����{�R��d�B=��U���7�H��ju���E�G�r�Խ2���6~�|�\�Y�U�aډ��e��#��<�)d<7Ԉ�:�kZ�zs��y.U��Tw�դ"�(��+��cʂ�1�� �E
�ZJ,ڊe��9,����l˛V3R"�7��t6e�hJ�`�Yp�E�,<�
"��A�O�H���݈�"�-Tmf��a�����0����ɭE���wnA=��m�j�@6��	���X�6y+
���!V���/�>tڳ�ru���l�ɩLv3��n][T�A ��L�0�j�)�V�g�!�ՙ%��<'����o�2H� ׫�'�5�1��k���5�=�ԥ��Vyp��b�����:��B5b]&0�*6�۹wŤ�,�W�cq0�x���*<5�)�k���i�JMѲ.������1�;u�m�t�X�khr��:Vk�*�5�G�@W��� �a����P��8�����!����Xz�ss/���H�z/k�q��œ�h"� ���*��8	�h��¶�2(Js�P~�XQ���:�t��}��xx� �H+dI��Q[���h@cwc���<�U�#��MC Ъ	=������R*Q�~'(��p��hP[�"�VZ�V������h�7{�v%7?	��[�Q^�lhў�>(�:R!�),��:^j}�Vst�<�$��`%{o)A����¥+���wI���ɳa����[����M^�])�x��K���C�N@�q>?�����/�N��S�D���P,h�nB6�D��nH�`��2*>n٪ԅ��bv��w�;��r�W�0~c`�9��e��HCɒ,R�Y��ŭ�u��2GƜr᦯�<kk�k]x��p��|p�y||��8����K��h4�E�[x)~c��=�ִ��Yf<�n!�n7&���q�W/SD�9��c�W��7Q�y�>��9/`����]��-�t�e��9u-���)���rvCȩ���;V���xHa�be,�5�CZ[��d1���t�[D�p1WMx+����1�p�N��)��&�6A<e�p㓔9�9�O?W|��u{����cU�(����"i+�4G���Y��(-�!����I܊&��[�J�{h��@�̡�f��of�ϗ$6��Ra��֥��X�a`cD��}�PG�,�GNX,Q�s�G]ʺ9��Y���8H���+ei�P�E�Iq�t^���'��h[u[���ͳ���Γk��	{���d�םɆl�s�P �l���x�)�.�͓�#��A��Q���0m�˿G"�jSXA�zJ��*��eN~��.�_��]y $�&��5�U˲[+֧"�:U
:ywO��a��xqE�^E]j�Uhdp��&a�7I����,u����>��C�����>�A�Fˠi%��|�XI�C�3XXҟJgsۦqW`��{=���;�֢�t�d\�A�B܋؛Y;�7N�2���Xe��2x�.��C��:2��Ff��l���/GQF�Xx|��`��xr�*�֦~Zh瀯 �9��i�.�cb��, ��3�hyԤ�,��"ܨfQ$hKj�Ӻ�={F�Fn�(�.����A
�U-`�|�Ȳp�;��Z�&D�FD�@	dIё;�nխN�9�l]�Ǩ���U:�
�p�.
���l@�<��	��FtZǲ��&C����E�b3��э)Zѻ9�$���ԅ�Gv�ޖ�xOS t�:��z=�T��鰪E���`�����o��&���տ��^�~���@4���{��k�o͉�C껜�]��e�,�\��#�h~T������*� L�>�m���kL`	�����2������,���:Og<.�ֈ�<@p�
>�z25:^�|����-�qL����+�|�؎*���g�Ï?x��Y�^37��vnN^�gK1 P��^���Or�pY?�?H�i�����I-Z&04�-m\�]�G��h�Q��U0p��7��/��p?@�:�i��*1��|8�WQ�-'T�p�9�3
��3s?��IY[\��NsE�|��(w��\ub?-M�@p�Χ��`���2��ë\��9u����Bk�>\Z�4�bU��"%�H��(�{˺�;18�ef6Z9#F�uהh	��qY���R��b�vsW�E��b���jD����qF�KK>�g�0��誅��F��&TJ�H�d˗���4�Qǆ>����os�ݵ�aZ�9pts�ɓINzue���'������0A�h���4�� ����Qg\ ���8�k�v�Ĺ�@P��2�plT����O�����@@�2�p�C/�N ��h�tb����H!�X 	�/�H?K3�L��u'��6�L��Z��QM&����O� [QG������*T�,���� ���yC��O?IU!���ڪM� ��i�2g2iͽ�U:�I��ڑ�XTV3v״��N�-�쓼J�Ś^[���,�.�, `�J:g1���o���^�H#�z F~77jϖ���"�lI2T���"&"����u�E{lԭ�A�"���5��ɁV��}2#+�!��h"��p�(��Z�3���wF=�FE���I6�\E�Y�q�Zc���	��Y�N�̖��[��]�7�w�PR���	�4��3c�T�y��ֻD�/hY�7@�iXU?�@�}NM+M?;��)�x�&��c���亀�
x�Ѓ�ʀـ�.��j�v��tV+�5N"�/�BB$-[	g��,"'�����U�����w��l�ȑ�~Sۻ	���v���zʧTR����G�q	�h>m�h�O�� �r|��7�+
u` D(@��`a"��h&7�%�����L�/�`�Q��{#U��PK�l��Z��.u���%��\����	]	��G�Dp�qM���n	�x���ԉYp�G���8y����K���{� ��
,�_�Ż��|�l���]�Af���=H�����廏��&=I����vvoXUɯ�v���{:�$%�x�������9���w�Ǔu������n��&\�X1���>O�\�CJ����
�J��3�xn(��Y-�z[n��ճ��x�nmv�?C��6ɓp��;�B$��N,�y����}�ׅ�I0�C��H=-R;�4��a�:�:zH���C��]a�M-���ֳ��bra�m��0��r!��:�NL�¢��άOrx����O̪b�G)��xS-�܈��_~v] �Ѓ�R{�Rp�DD_�<U���Dtwv;�k�����E�y�h ��"����? � <�djd��k���,����e}-�ը]ʀ
?�RX�O�ZP+~�\`�bsf`u����~\�U�� Rђ��t��#P�}���} %,;p�8g�����4 �n�%	)c!��j��Υ��[kwV���L��������}c�b$����g�M��F����-v���Ng?�d��a����<�@�|�;��Ki����Z���:�K�֚�5�|Rg 5�TE��b�.e��	q�j/���h���3Zؠԃ�V)ӴRAhp��rE5XrU�M7�y$A�4@�,�c����4�,q��=�A���*�M>���b�±��V�<PX�8�u�9���b��Q���$j}�N�7�5�&�D�uJ�%�F�t?���$� �O
-7}��������̇@�ߩ�UkV08,Bd���X��&�~^@;�I������Q�K�פbύ
�"�-F�B���_��W��뽀($6�{��g�FD���6L��i�5�b�<�4�)��+� �p��#�c�i��P3�f����R�p�)��D��֪w�����Y�&b�~V�h�[�2!����.:��C�R�t�b4��0��|�˿�M�������3�7@�·y�l]�.&顡��:�X�ݘ'�{�g����ʻ5�R��R���� �w�w���0���ØP~��:���`��>��*���	^���Q��T�Q���Z�оBiG��b�.���ޔ�	!<�j5_���F�d>���Tp��"��͍j��kVE���'+����]*iI,���OKR�pcЍ|o���Ւqm���"�>q�K�2!���E���R�쮑q��v�K�o2IKi-W!�X�Y�NԬ/<��S��V�9��S����ϣrdg r�]~��JME�t+�p�Ά�Aq�p30�qs1�-��5�8���̗;�]$�mǯL� `�+v[�*���]>�9����6Њ���R�8����UF��m�`�sZ�f�N(�޳W>�2��ƅaQcB�c���
��N6B[�@�rp���kĽ!7.2m���-h�M���`	|�Jy����$pz�1w�i��<+E�2/�9�s��h�wP��.���\�K,D�����A�,���B�Y,�Ӳ�� ���&�4�:�^���}�ڼc�ޞ���ƚm��oG�K��׺1�f�)����}�'� i��=�������#b����m����Y]m���쾦f�5����Rd<���>&�R|٨m�U�b/aqk��8Rw�$i�d��*au�q���DW/������!�b���U0N��,���E\�w�����E����]��������wޤ_ˑdM;�Kuc釻X@��<���֞�Y�e�b��(nם��p�*�6�*D?X�#�,�O��cY����Z�$��ϼ�7�XȍU��\��NN��!@f�\&V�^'8\0<<3�h��Η)�6���dd�*���e�A�܂YD��>���-�L�k�p~b/s�C�1�E�=ͳ�Qg��&n�a3#���Ζ�v�x�=H����4-M�7�?$j�xG���:d���2W1��yRۤw�I�`�\e@���+bqE����xܰp�q� RC75���ܔ4��h�Ԝoy�ng���^�y�Tk��Gs>��ɼ�aEG��IAɛ��'�Z���p�Ck��dј�9*��,��V��}2��&~t���xl�6��`*��k�T�A
W#i\.�A�dň[_Q�;Z:��<Օ��9���4 ��
]�;͘�ϝX�YXJ�^Ӕ����+˽���+[��.������2]��n=��w�� �<��"���#Hoﴄ��.^k>4��B�+]ױXI�y��~�Nݿ�=(~+�o����y/�}�n,Isi�bU��j�=�d%YQ�hc���p�q�n�����L6ĠF�gPy��$3�"]��	 �a���\)��՟�j�����?��F�s�XUQNN�\u��ffɄw�^����%|}�"Jd;�>���޺�j�r�bsu�{K�"�f���h��g,����mndS��wV��J��Kֱ��σU���Gi�RŃ�h�GZ�5�C�+`���zb\���X���a��˘8��R@�ڼG���jy	>V������(�X��:�ǳ�rKxs���,)�Xa�*iE�0Y���}�s��װ��½̀j��k��6�B��L���0Lf�Х"��Z��}�!y_�동%z�ψ�/`ڞ}biq����j'�(6��6��o=�Y�*�W e�r)���[��Av{���}��|�o��&`��o��`!ii=8m���]_��	�������ಖ�5D�Lj���I����௿�*���_�&էif;d)@�|��I9�`�3�3�PUt�U�A���d���c��Xf	Dq����"���E�,<�VЧ�^7!��o�MAՊA���叿k�ҏˆ���X��ِ�xa�q��R�z��r���x»�}�=e��?
��f�4��Sa�d�R[����R��^Ưb�QՀy%r$X���z ?e�lo9��K)���1k�>X'�I� ��Nb9�
`��,��~\/��ϋ��{��M��f���:�2��FO��F���"`�7��3ZS��e^Z��{��8����5�,K�2��Ԥ��Ȧ�F�d`�cd��`��F��c�R�B��ˀZ����3�E�5Ϻ�Ӧ�v#�,T���"^��Nƅ��0�JY������`�>���j�<��j�P7��b��%j��b�e�NV���p�]vL , �g�|zN�8�d¡{�˿2G6j����Vy]��C77���H���]g�w\��;vo�M��߫��N���0b���+��������ɤ<X�\�HɒZB�<�mϋ)~�i��\��|���d��BP�a#��Y��)YM+�ͪ�l�u�S-У[��4�E�����St1�/�KeQ�ײ�2�Gk�J"���_�1�qy:>zYA�)%N,��H+>k˛��(M�R�;t�˾ؘ�(~P���e���.HHY�y6�F��`�eЊ%����&�R�\�U�V1�wL�%���,O�=�����}�_o���|c��Y�6@�_��6�ɩZ�x�Jg]^?�{���*��lj��N�#j:^X��ǫ����֟�h��6S:�s1�Y@�:k�#��E��U&�7��b������gӊ�f�D����ȿ��7
�:�%��k��gI�V�������U }2@,e��"�`j�V84�+�O�ĞGI �=�Ϊ��Z&�^�N��ں`z�@�Pf� 0y�3\,�����z� RXKHՄ�@J
����m����ZvR��U�?��k�r�6�b��H<!۱��b�9�h6���'��v�¼q.*����������}R�b6����o�L<zDNI:rh+��E��<��rlyz<�<���3���/�)	ܠ�
6�O�d�$��9���l����7@�g+�[��$)�''I�/Q�v&?],ӰV�K�=�(�Ǔ<�nn���M!#��<�1V@�j���oZ(5m�\�<�:�H����v�k��t�9���5��Å�J�x�/p׬Y��v�e�	�L�/����m�	GUe�oP�l���v0���}X����N�*�{=�Ț}W6�*�òz3=4�FMND�z5�a!�ߛ%y��m׺����#�
7�V�]�E��Ӣ�l�w/���oJk�����8i��p�O�Hv�|���5���� �k0K¬u���d����y���C�����?>.���$\�dUŊ5�=i@%jQ(�=\���h�YEs�(&�4x;��;õ�l�,��~0O �:��L/�C��Uӱ)hK�*����9x-h|t�+αiZ�i�z��ì�:"�nX/ԁ��ZV��&N��!u½��a3�c]ב�&�"Sy�O�\���C q㥼 <&u���sN�yQL7���w.F�X�E
P����kCN"P}��@kؤ����m-���^ܤ5xne���Fp�`�*E��}Cb/�!u��U��I����Tq���(;�h XU��o����K������U�U���:G��s�ǹ���e�K�<�i�h-2A+�)�mJ]��5��Y�q�S4�u��yʩsy����D���u��w<��Z�uU�8.?�"�9�%7[2V4��3�sD憖J��BO��N�@F�6�f���Ho'�*[ �s�e��%�j�S�I*��|��GѼ�vek����՘;L13����6`c!o�5NwBH*a���d�Y:�j*+�[����N� hXĄ�@�8��nj,2ȸL"�@	��*(wC[�*J u�y���WB����Cΐ�J9����x������1Z��Xm�6�&��rR%v�^[4�G��eN͖�X���V=i ��/d�-o�T|���y���ۘMO��u"LΧLF��ٌ�h���?����U����ִ������T�iT7�--�Y��Ά�d��ڤ�jY���"����9 ����zi�굽�F�|@������RU������,��i���n��BR����q����(��`�0�sC�L��2LO�W���11!~����n�j@�+f�s�z�t�XF��I���Vf��je,������h�p,&��1��,����"��."��&!�o�>������'�}Y,&X��rJ��Bd�I1�$[�,|�MuSrէɀn(6��>�jB*O�g<�/��r]�H���ʳr��u@�Qg��C���b�}q�eO�i����V������SaOx��YyU5�g���d
P:Ʒ��Ⱦ�cm!1�#�����Srg�w��F���<+R+R��D����1ڜ��c�>�1�4��6�3���uf-u��o
�֨2Qp�n6�:��fEYy{�����u����щϾQ�Pa��xhj:5����+��mj�*;G"&��2���!�Ɯƕ��Ճ���ӷ>Z�(�i�o�A�������U_��k�z�]H^�����u(�8���=Z;�:�<�L�B���&^h���!X���q!e�U������'�rÒ�SS�m��X b��|��&]��!;�<{ƌ�ܢ���Q^���r˃EZ$z,"��w� `�A2C.�AlO���I��\Q,row�i���y:*��,-��
Pj��E��d!���#����xJd���eH�r��)�-��d:'>���;����`��̠ U�V���mE�04k� �uT��4M�� w �f<��F�������d�9m�l�GkU��0���	d�z�5ǌ:��V�l�g"�C�(>�&Dm$7ٝ���?l?2;�a�b>���~�f�V�������%S�v,�@X�k7�D�b�cށsv�L��Hq������}0ts#��0��e��ӆ,��S�;G��֛K��y��ۻ�=�Ju(�V��2}��� �ǣ�(c~P���ޢR����@���ft���Y�F�Z}
R�$cP�|}�\]e���y��|'�����Q��JA���R,%����OU-��źā��*5�E���ɲ7����{ʁX�]A���\�l�C �e�He0��k�w�b� ��,-���,O$��i��V�¹���1���,<�i�o�-�����I�Fǡ'��Ⴠ�6���2��n�,&��kC3��B�0���6M�e7$ = Ǯ*�<�$ޫ�`S��J��IrD��ZXf�{ �ů��" 
ks��\xxH].U4h�^X��>�����r.¿[�����g�,��8���l�|�N6�/�ƚ��gSOX.���⫝̸�`R�J$�̡��A��Yͫ�*���k~Dm�㳼�VlG:+i��A��4est
�F都5���59���,E��]��Ȅ����r����H�E:9mPI�6�v4��cQK����%ܜ���+��Q{|�{�Uq��E�� p� �{��Q��i�Ө�R�SI�Ԗ��G�Z���w�mč�N �#u�]ds�h�"�W����,4惣en��9jiD0�`-݉&�����|���2v����Q���\��`�x��
m�z;�Iw_;�N�#�[��%����{'�9珬�c��l:r�Lb�¼2���5N�2��EB�����>Z�� ��w�x(=�\?���Jz\[�Vlg�b�TJ��E�4d��b�!��wH#�J�[׈&�f��p`�fFf�6��ڍ@�����w�{X;����XT���(�x��N~+:T���:��	�
Ny�^�%Vn>����1�$,N	,8�"�N��| �|�:Kj`2Yj%���t��F�"3z�U���ͱ��&",���8c�%M��{36�;�h�j�UW�#�s*Ni-& �0O6��-{��nQ�F[�w�P���e3��b� �R��-s}*��0��B
*�2�ޫq�&w�ש�`�;yW����jR)UPx�!8�AL��v0p�E�j.ގa6�z�G9�F�A����Ң��b�ܝ$R+u?M�'���x�"����I��e9�U����ֱ�O���_K���kv�M`z�����?-��r���í�uF�t�����wk�Ɣ�dY�J�c�1�yp�TZ�ًwP�P�fB+��U���H�{.葽W!b{���ƂMʱ�w*#��HA�,�ld�@*������ʤ���UIU��1.y�=�F(��Q>p�NX�8�gQ�ה��1�ai��A��0,�\xy�l�l�<�2��/U;P��S�}�R������<{�U>����C�@�պH�QG���K�o\�(�H�\�&�#�\��	X��V�V�͘E~kYO��>]�s��_7Y_����t,]s��z}	��kJ�5X�M-lm������]�\Ǒ�-3�zC@�C�/:z�����:3g$��譖\byann�7��M�R�U�D�ů�����#� ��rրٔ&!����X��hbrڕ�x���]I��+׽0������d|	�4��Wm�<!�S�?\������{�^RB_�t������;o�a�=� �葪Ur&��	,�x^Ҡ�]�!5j��9N ��=0;��X�l&&�Euj+��l��بxl�zVj&���U�~e� m$>������U�nt�mLz�RRY)�_<��i�<R�'�ў�M$6xRi1#j�}'v��ÿ��^��-\��������x�0�',�-�������xSN�Jm�Q�p.�#��������=�0��`-��xN%��L�4���)3��41`�#��&<��^1:�BoA��2����DI@$���\��o�-ś+�*F�`fm�x��r�"!$�,ym�z Ytb��y��y*�c���;��wh�����b�(z�{�Q�[�����D!:!`ͅ��^lY���bc=���M����9�'�R�\t��y�j�Õ�HfMb�x��m��b��u'p�KHoBi�~w��,�}$T�8������exXą[aO�L~R��ٿfy��w���O��#U�T-r�9
�ڨ�uR>��T���>�����W���Aԩ��?%�7J��YL,$x]�a���y�87�iEuR_"b\J���V6T$h��ԟb2��SP}��:�Z�Á�'��f_ �\�3$���d'��6X�O ����a�'��.~�s�C�.� �<I�e���(�['8'�='o��G�vq]$Z�q��X��K���s�)�a�x��&m��=�j�:��5��7"&��!k��{B��t��{�
&�ޫ��ދ�jb��{���tC����BnҮd��rΚzP�h!�J�\ͼ��.�"�T��cN�^�n�Y�v!�/�\)m�܀IV��]��WF�ɓ0��t&����z��א��K̸�H���*����6���/��͊9��yW-��eF��QB	��h@�$�WKD�u@���]j��������d���Ζ4��,AO~'#1K�t1\b�D��@윺���r]L�јY��ML��=k���v��m|�:��Q=?)#�����&iR��c����Z�۪�7�6!�F�$�'�q��(]'p�¤~�.J�D����hS��~»C���_����~?:u��*��2��COvDh5�3��Kv�6Yx�+ �g;Ο%C,��$��~j��.�qŠG{��J��>�����y��Cv�8�t�d��~�I�,
����&��^r��ѕ@CӜcm/ա��0LQG��W�ܸag�L�%U���*C�h��;��=Dm��؏�e��cV����3 �%	���G������G[O;{l�;��m�EO��}��?������0~V+�#�dE�ɾ�t�S�o[B��0�U�V�Q��Ѽγ�Q���/Rü&���%�����^[�#��8�B�J��:1�D�7�ʆ���A8��c�,�`@���_�YV����C��Nk�;��1&���8Ąѐ�V'�'Z��Ε!|��!�ѽ��j�:�9V6Z�ic<�lf��g��G��9B��k�q!����<�U��2�I�E�AY�,�GVڙcd���Y=2�ΠP��tj�QY����ƻL:O�I]H�:d��E>�:Db��)6�H�*��nL���������:���,Fe{�ƵQ(q_��Rm'���U���H���*����zD}����������E����YQ�'�"��jG����x�Ӕ8��m�c�7ŝ�KQ���&������~�-Ϻ��*'�18�$��H��LS�S�;3��\���ȳ�,����x}w׽���x���b:/�/>n}l"�F���'R��5�E.Ae��Q���H��֠ׄohE��u�i�$I���Ʊ��
�5/������v	�ur�L��9xE�A�F"-����Dw��z��V+ؾ:�e�,|
C���E�Z4�����{�F����P����P���!����N����1`tL0�Sy���0��|���o�GPӨ"��e���"x���h\���Ԑ\'�#øj1[�F�u�uV�t�Р��mdb{T�g��H|�����!u1��Zw��8�����9�oܠ��O���|y.��0�qD[~�.�(A�k�f�h1b�,'���1��Tm�/�,�G�j"5�SK�ļ�U�d LSUW�ռmw��H!K����pA���o�!ݹ\bx��W�P䗨�XU�e��,7a���&���vvj�'�bm4f�����V�����2��v�urm�GSvTм��6G�N�q��n.�n�֐>��
�R�v�4��Y'���������^8[x�E^!6�S��Ͱ0���駟�+�LY���8c1�qN hN-y�4�r.C�2�@6�B�y�&xE��q���E��e�^��7/�h�V��5hZ�;T�((�(��ׄj�ucb�T��^�{� ��w�f�U��86�Ň�p;4�r\zx�a�[}ڨ꫅�%�4����.�b	�՘���3o�Īʺe��?�C;zh\�9|������0O�!�&�^�:�K\�H�E�:�;*�g��ĴP�a���Yޭ���zx� R���k���g���&�-(A��=����p}4�3�{V#]\�� �?e�w;�#Rf0+�XյdR���klb<t���}`�	+�Z�jiyT�-��<�'�b�\I'�e�"�����q�[;�ｙ�8��6�/b��"�KB[ު����|~�������ܣ6��8�������5U�]�g�g�^ӧ�	j�L[�|�9E��"�؏A���*�!�a�H��h2H�0�lPw��&F���Bc4� �j����y�ڜ�l�u�
�'V�D6����5S,�̹��9���0B��%<��3���3C+lr�a�x�<y�F��Q^_�M���f���Ä�_��1c6���~Rub[ԙ��L�a����B8��4��Xlx�y�&���VB�c��/�BcX�z�Þ�[N��p�b�{�����5ʒ���O�����f�L��CHu������Kld}����`Ʌ	?7��S�a@���!&sp��Dխ~���eyȉk)~�y�N�7�������*�a�OJLL�ǆ�}vu�l>�Et~-H��X��&�CLQ�M��Vp�����t�f�?��T�O�s
��*���NC*�#�P�h�H�s��S����������Z������ap���>b�M�\!�ӷ�H��u��joTɚyJC��y�m�Y?9	b�^��3j�S�a�>XK\��� 
s1����y�p?ۂ2�$�F�ܱ��C��V9�p2�h�f�I�o�:��J�q�ZiL{`fɤ�ׅ'��C��'ǌN���X�0Qᢼ'z��H_X�Q,���v=�΃������!�8�%_��ҙ��^z)�Ѽ֫H�J)Q�(CȪ�=&�ư՚��Y��;5�"E1u!�&�
Go�l^&��Ki�F��%�/k(�d�#]X���)x���5T��Gj�ӔUnHƿ��ѣ�ѓ0�.�O�9�v!��e����l�؇Hs��a��?/CO��� ��v^=�q.�T�F��[�e�?�qM���z��7Zĺs'�q#n���k����3xR����kO��7�g70Z�鮒�sC��$/Űϕ�O��F{���SײTc�z2����=o;��\�p�)��[��o4,絥l6����8�ʂ-����}��8�pih��գ�ˌ�RJ$X G�j���s�%�w,-�q�C$ar�HE�=���|a"�O������YX넻�O�9������~�(�I/��bJ�����Mx�
���'mS_��̜�d-Q^�ۈ_���Nx�mRA�Fs�4Q�x�5��;O����q4�=ʚ+,�����G~8�87����$^�d��[�ko:^(i9�gQ��lrgU,��Pˁ���8JE���ǽ�R^�Fx[���%�Ue�Iq�j?@="̣��1���=ǌzu%�m>��>5������q��:��ļ̾�V�&\mQV��'S���e`cF/:����Դ9��.�zݠ�}
Q�������^�+cT�
�J|���M��еp���۳�N*eyh���9�4ȕ��o`���{��Pڈ���]��Dn�˵�!���y�۵�*���|�X��`"�������6�c�K�%z�%������J/�T�e��jG�T�fo�oebf����Xě�}r�S.��4Ҡ�i�{��`���jD�(;#Լ�0�x�]Jrp����� K甴m9o?��Y�"��/r��� �}9��'�"ђ1�Xm�˘�tƟ[�0��prN�ic�'����B{f�S��,ܹ*hpQ��0�����x�m�Y�	�0Y���[&k�x���81>Q�X��:�z)�s�)Ts�a3٩"�V���$�����;+�H>G�l^�������]�޽�L�P������LF��6"��C����sw�v��Z��9����>D|����Գ2d�bS�_TU�E���k�HPS���}j�*�ѕ�k��ũ@%
��FK��_{�_�R��}ꛊ�y��N�X?n�u�p�W���[c��%�WSM��j�	�+��{*�8f������������M�l�)	i4L:0V��l"�}���;��%W�n�k��G*�K�2(R����[΅-&v��b�]#��ő�u�Nh���g��_أ�K��1�s2��if=510��7�7���0/�Bc&X�k��܌~?GV~v�p
�Y�*O�)��
�8yr�lvC���������pb�y��z�B&��1�?��d��+V�*�F=���aT/��d{���+�4��F�޻��$=��% ;�D�i�O���0���]�=E[�@r>������bc-�d!D�W�K�|����PL�0���³��2��Gt��,�e�f~���A9.A�R��T��Y��־����Bw�����d[t�%�|�S����'F]F��/�׀��<��_��_~�8�|Mh_��ֿ���pÖ�8gG�}��6H<���bۺQڅ�&d�t�/!h��z&�zE��y�\�0d�0�kV#���Z�UY��q
�<2���pu�]��� ~�(Y�)NpyP���1/Z=��7|1�d�`���AӠ�Ӳ�&h�����.\��X������%怂�Ml��/��=R�9��L���ǸisTa���<�#-1���L,�`St�s�:l7�fP�hs5q������ߚdX�g�&)�M�����YZe����9[�DG�06<R$�f:;�Ƴ_�{aD��ߕ��T����z���}�v'~� ��1]���.l�r8̞@e���˙sH�U�p^�����T�'�Z<I�CX��mo˾c4���I=�[�杩J�uh�$��r���e�>�����������:��(�^J��x����M��.x�ʵ0B��1����:y`c��C�Y,�<c`-[X��d�)WCeH����:����6��������;''���%���I[��j�[W�Q��H��pJ*��=�ND��#eѦ�f49/�5�N�W( �?+k��P���P\����a��kum�PD|O�[{
�_��k��6:=�ţ��Z�p?b JH�dp~�j��hԉS��W�ę*G���q�T�S~)k��*���:��Z7A�(��
�6��e5��<+�x,?���Ex?�
�CC�F���Z{
�b��9`,��e�rث�	��D��v��6�$11�W/<6�5��4m�[�;e�hC�kQ	�A��XlC���.�Ö�L@����[�Q�SJƉ#Ne�^�Y�M�<BnV0����84:7ICD��r�K���Q�w"�O�}gc��������kXM%�`�,J�]e�u�@u�S���:e%˟	�Q��*,�1}��!����+����/�#*l��]�a$n�/T���M��Kq��:I;ym��
g��~��*R�������R�nW�\I<T����KPEwo��j�l���8�*4@>�T�W�YaPA�j|Iaq=V�k��mʀ^���`[�����-��K⻗�14bVTU?*]f)�,E���6T��;I�0Z��t�2,��^ᘕOa-�gpu�u�!J=���Q�n-���$zA���M�88������a�⌆���+z�4�T����}0J�"q)5v{=�*��UҒf�<��j�tt�V�����`.����ګ5��A]�00��k<rB%�@5G�9Z�!;��0N�)[�d+�*��]� �<�M1���~���%��v٦?-�;-�r��.7�j-R9�%��*��-O�j��{��S�U0�L�u>�>.��(#'{v8�wz�e�
�����Z"��7����?-Uh�lߢW]�ʰ��d�l��ڽ�`Cr��g��c�A�Q�3�rq�_x��U�[c1Z��Y��#0"$cA`�C���33YmjiR
������j4�]�Fx��%�1��*oSkc�5��A�Fqlhp�T��*T}Q#<�����D]�r@��/����gB���96��%�C�ɴ)��>UX4�x?�i�i�
������>60<旸D;J�(6����֒{�М}��r�4(��}Q���Xm+�E�+ͽs��v���#}��Ƙ �?pAq������=�����	ii����9ۄp��ke��������eV�^�%�.��M��U���H2�{O�8�{��y{3�{W�W�fZ=��&	a�X7�Y�7�P�n����>��bÇ����QӁ���y�8F�d]�e�����̚��&��B7�5�HQ��1"`�V.c�D�̐���j���7:�u_yֈ~֨^�Hݻ�|�j�3�����RtJ)#:5�{p��y��zK�d�4��I�ZxOYD�J�����㧨�)nr
r��z��Q�1�)��B;�ir��l1� OmH8���:K�H������/u͉<����ph��X�ա��&�ar~.7:\��p�?������Q�X9D��ũVY�<>� b�Ȉ*�=�w�!S�wG/FJU� �k�D��>�
WG������6��Cn�ݱ�27�˲���W��D�V��VO��]�
�����_\���»#EG-�����߱���U`���a=�橞� /��C��������f��x�/�cOZ2��E-�Y !j��^J����)BK��@���q��^�!3�P��0��#ᲄ�t���b�R֤����,�ōxmrF����6��/<�3���S�{�~��6�[��Ux�8�
Ee�m0��3�>x�ų��B&��8��3����ԃ�%Ԝ��I�,�d>�O�t�F�:,F�:a������6��C5R�i����^V�Vɬ#~iz��þ$���-���` ���w����m�|M[8.��{��"|w�D��gñ����sh%�V���x�B���$�y�Z�����vUE�,��0H�����B,�ˬ:�O�����7ՠp�(��^��ƌF(�Yv�;�w}x���g�6'����Z�ŷy����y�z�р<d��5�Nj'��ҳ7�c��e�C��iC�Ϥ��ͫ�:��J��r�V:�Jzw��<*/����n��c��x���H����1�J�l����tfƙ��1hs��	,(�jE4��hE����`�h0��<U�9C�֡�5����t�w<�Ns���G+���y�N��}�2稒S��%#��=��ĺ&�ٔ'���J%_�^�!;'6J^(��";C}�|q*��{��$[+3�S��V��ճlLXM}�֥:��{�Y�^>�p���S�� �]'�?Pڷ߻G�ifu�ɐNSbZ0�M)a|EybR��>T���:q�֬/(%��3�3`�O��K��R�p��c� �E9-�=(W�Q5�_<�H.�O�1�>gӄ�؄��җ��E	���,�x,j��ɵc����xn�_���X��U�$EBT��A��ۅ3��Fc�n�%�|9����#'z��z��r�Y�E�(*H9$r�j��=E|��zP5^P`&7�y��1���|IE`*�g�p�Q����.���q�m�#��;.�lXJ����S8?������'��`�L`�+�v������k��,��z�P�������y�L0�p�0{���]�qza������Տ��s�#AW��ɓ�r��;�/�oSk��j�57�H����u���[{�/���*��S}��(oD�H�p�L�.�)�2R�U]�^)OzQ�`\���1�}X����0Jd�atL�h�3l���8��:a��AM�v�O�-!�o[�M,�z>G�[�]YS1x��G��,�EC&O����՚��yj���Q��������}�]p���?y������e�F�޺��Φ߸G
�"y1T������C������&f5:\��ۇol|��po�V=t��g]�e�;X�Zb�� %BzU�-�mR#ֻ��c��a����s�,{����E|�x�Gw�l��
/�/���;CW�؄=q����"��q&��H�5;�dG����#�I���j�8�G\�WD'�u���?�P���d�0�'���oT3;3Q����א�X��OB���X���N]\ Ƌ"��L��P!�cL���	j� �A�Ę;#������6�B�sX��P���S��3<��jc��&���g��T���V� �7�1�1��H�H�`�Obn?:q�?�.�H�2��i8�%2��9y^�gF���~c��/��4��u3��׿n09e��]Q�(����L��E�ߌ����1�R�Z�٩��Y�K�y󚟻,��d��{S)}̼��;�� ��
)�E���0��66.�;]���f�����I┲��n���N���&p��Ơ�K�����f��.�e��'_�A�!��5D;����D�a%'����om�gf������A�xyk��P46/��Ͽ�l��9P!ø�7j��3���b�/�P�3��2����Ӓ�[�����+���5K��mq�s`�[MV&�|ѐ���1N/�B��14Ou��D�Ԟ�~ �����e���i��{��A�R"eT*w��1����5�H���W�Q&�?�:	ѐ����=�X"�Q#��`��yd�b'n�T�5��}��U����iHk״�~.i@􅢌�d`y+FQYo�9֛���+����y�0�*0L�ѹ_'ǽ��)S�d��~g!��:��	�{\<��wʴ	��N�]x)�`���Y�ƅN/����Z=��!�r����|�M�!u� �|�#C��M�<8����^�mX�z������NbO�ؽ;^���D��0�6
�aE����7yph����L�5Ż'.��\S���Z�'�2[��uS��s�Mc~�1w�2.�yIKIm�Kx]0*=Og?���VS�������o����1[H�m3s���b�EG��Ѡ
�s^���~˒ԤNe����I:7q�>C�:)����m��TX֏�N�6��~�a�Qm���jG&*�J�����Oj2�K˽�0ܼ�6��*�&���aZ����E{g&��(;U�-jYmO����NU#̰�Ru�����dlaGa����>^{��aP?��r�6/zƘ�@�y��<������Q�Ð�y��<e�=��M��dOr7�Íp�^4�������-$�͒�m<�� =�ʾ�ln�ML�r���Dm,F����Y��DLa5:�g����d��8��_ܠ
8�D�zS�t��Qy���K��>�/����/-���A
u��x�*N'1�l!�0���˛�c��S	C*�S�k��r���G�F��{��&Bz���/lC��bob���`�7��W|���e-_<Ǎ��(B�D��=�9O��D��z����LTc�{�R�r����������P�b��8���+�g\ǎB-��z����d	A�S�����Y	��5�'�Kx�C��a\$Wi	��D��8l�	����ޫ���%�UF*lB���䀩v��w{�|�z�3��;�O�@���5��й�s1g�̉#t|�`�`���zmH�K,���Jks�o�?��\�>�����T�L��40���(1�4xt�w��7<Oa���PWHe��wVJ�״�f
5��ryW�V0��!	0I��8՛��a6#�J1�p��Yܣ�! �hL2!z�E-:�@/Nc-�,#
���/�����3��N��U�m.��i�J`��	�:8��)���r�6��2�T<,S��^6�'�p������Fx�֮'����[1,�tB����:sC��%�����O*X*wduZ�^��Eo,S�9[���j4�m��6_Cd�J$���dD��_b�K�F�7�zC��!f�I���Ŝ$���� :DjfHu����U)yA@��1��jh/���)T��Ս,�܀ޯy�M���/�ϥ(pɾ�:u� JoT"�5Kf��+Ѧ����dᎈ���ɚ��SZ����T��Q�f�?/Z��PJXy<�0�� kM)\\Q�X�}��//��7N"d�1p Q�alY�o�c���/y�O/�5���tTJ7��{��Q�(b��7o��]���׾�'�F)԰��[g���P��d0��E��ް�H�'o�P���=�.3�u8ӵ��K'�*8p�cп����\~����l[<���1�2�C��%�Wj[]bC	�z������.��F�jh9�%� jR��
Π����R���5�𭋵�܃qҚ��E�J ��ߥ80i:���ƒ��|��Y&z)j�Rx�f<'�2.F��F/�<[�Cu�(�`�G�!3�<fe�go)]T��3��D�����3�e:��5<P��@���ָ3)��̣��sd�	���	�'(���I�D�A�����6��)�f�XUvtƲ%3�W��%
�֖��̳�5�I����z�Z����*�+��C��Y�����fϦ�xj-2G�����S���B�O�f�0P���.�;$JI�a�ؕh-BvIؖ��VC>���ۄ!������ :���0�2HN,P�#�G�\��FDF<�h{3��������`��B@?��`���kEbc�l7�}l�;)��6�wVf�ɾ����Ӑ*a�'��Gw�*�@�^)y�X!�kA8uK�,s�~O���&)[�;\J�nӒWUAF _���xYhPsF��/7Zk4>��9����tP�RO�����l����p������$�C�J�l.�*�����hU��Kx�T@�v1CJ�sDe�"od�UAm|�_�ͣ�c���E�5˦�iɲl#�7,��A�[0`4_���^�5���Mi���%��1���&�7�zEk���65;�V�1<oi����u�7��o߆��9�&�O!,W	�����P�5&G7����J:��e�S�T��@�kr-G�5Q���/�G�Q`Ѐ���?�:�ym����
X�FG�E�8R���k�*6)�h�&I4�F�*>���]#�������ų�<�aP���%���9�_�Y���7�|c}h`�@���{����}�"l�A�+1��hkR�j�ӝe�]�Lџ��c`�)'���J��ᆆ前P���e�}����K)W�_��T�\KI�)d y�ڈRG#1}�e��ݣahmۅB��f��.>���#{s�����A�sw��8Gr���P @�#=�w�ޗ?���������?���s]߳-ek��&�]�+��1b7H�b��g��MGB^gaD`olŐ�n0\ޓ�>/kؕ����������?�S�{��ŗ/)b�8��Ƹ�B?c^�="�RL��YNV"�_�P�9��b��W<VL��J%�H@�~��N%��~vo���(cu	y�y�S۷]�M��(_a�� tʕ�D�V�N� Y��U�H�N�!�Iv���6��r["��.����9���M[lEb�xRJ�/߮���o����?������u���6�0E�-u��x�����iؗ��>��("�k�.(�J2�7�2y����� �p�6 :�F��߯�~5o�.²G� ���}K���(���7r.6�j6� �dR�~뉦R�� aК#���~�UUh?{��Z�섑;)��(��FΦСA��j��3%%�:�q��� �,����Be�;�ڎ��5�Ю�39�X������eRy&6�;+ay�����簔�G�i"�/<�r��[�FKf��e��^���Z^,�?3���Ǯj�����}�{z�g=gh�����Si��R�rb���ـ���j������S����H Ó'���8��kJ��b��Q�D�+�a�4��Y��2���7�����u2!<M�8y��2����n�y��N�!$����0xƭ�
"U+)���J�������H`�~��5����yx����0����iT�D��\��t���R��nz�j�a��Rj�dl��F%V[�%1J�1VݾȖ��K���V@Y l���ٌ ��yA��b�fl��������h�0
|]N�J��z��V�vC*o*�E����2ň��%�tx�T�O�{4�k���L�JZ�QZhT�C�LQi�eF���fE$V	�Ⴭ�c�h��!�AN���\3�A��;��&�����>���*�i��WUr����?k^�v:?�8?ɲY� �#�!�?�o,d[H-�,V�h���!
\$q�̮�0:���x����TگD�œ��H8H���L8�ơ�O��9Ws�ugbV���`��^n-DEp$�NbR���Ya��PQk��9)Ǟ��jD��s�4��Z�n4�ީ7f8���(eE�����T$)�ͦ�jUR�#E(���?��_=Q(-���������,�����}�wkx�/�`�#=>E6�d��s1zzФ���\���MV�'��Ï�P��P�0%���~�nQ)��5ԻI�ʊG
u���+�Wo	��ݻ��~���l�Ta�a=��E��>����%S���?�`�����qoOV���^�z��������qfV{x4B�4����59-�T���Qk��jۧ(��|燽�w^���Q�0�a���(���0LTfS��d�1�f�5�Jl6���GG������k���m)�Ah\���6��*� �e�&|�a��䆅	\�W�ְE /��[;` {<Z��2��#(&��p�����B�{O�R���j�R�V`SE��#��R]��s#��7J.q�g�-t���_Z_����\C1�ʔʉ$������դk���p�5
?B�Ԩ/~
�	Q+5e�M���d���G��'2=)�&�:Ϥ9Y�k2Au�S�#0RfY�8���EU*��N�_���=9��0ޓ���C��K��̋���k��~�K�ʹ^QHt�T���{��|�l�� �����_*{'���E�1�K���axjH��"�Uޕ7j�U<�\S^�M�<y���
�a���"��}�O;�f�>�F����&�g#1g�c��J6��V���s�����n=��.m��d����4O�����]P���\w���g���5��5�}��C�\��Uh�^_�0^m`�dWIM�	"��$g��8�P�.���j�*�?y�T��.U>z}P�E��C\Պ�*57�xԼ�j�?���=���ڗ�o���l����A2�B�D:�^�^��/��g�:#�Ā����xo'%]TՄ�`f�\�p�����������]+����/�j�'�P�����K;��;;�%�E)U��G-���<Qy���\���q��	���sZ���A��o�?&�両QoVO��z/��"�i��RR�,i��8cIƐr�=HW<��M����s��P��<|�ȲN[�^���Q��!%�4j��9�i8F�s���XY��T��yD*���Qk��.��6�p^8pj}��k�ki=����Wo�h��2g�����AE�d�F�����N�U��gS6�-��ڐ2A+1�M}l��}��x8O��ٵc���զ>C%��(�9��C9���w�/25_�����p]уڱ�\bǃ�������>���d��̀b.�$cy^f/�X,����H�6�X�j�[�(� HFi�E��$m�4��3� ��?�33�F!ZԿ�ۿ%Bэj��$u�1���CM�T�d�j���o��mA,F�Q�r��tل�x���=z�iЃpo��l�:f>�Gy�u��W������g�y�ӺDH�<�4�U�Q�~�`Y6��>�+m]�k�l�k����56�u�F�F5�l���/S��M[ym2��dK���-R�ғOYH��z,�%n<���f˵���t���t�.4���,{�Ui˒P� ,���lE���C*	J��{��9�S&3�����M�Ç(��UF
xH�{a��Qs�J�,����ֺ���b��!O��f�ȸ*/�WF�$�g�����J�~Y�W��N�Pxs�^Ix/�p�҈j��̬� X��ݦs�H���htSyGm\A䕔&d|���?��&����Y>��C�����aSm5�'���]P���8�<0��γ�N��VZ�X-
�A.�k'�D��EZ6����������~�۸x_��-�1%W������$�zԡ����*�qK��[��!e��5���}��os���x�����o?��%����ŀM���_E��8��#�����*R3g��:3�]x�˒xp۶��ԃ,�8�5���I���7r5[�V�Ϫ�g~~)��z.��,��b0j����1A�	b�0���Gz�p���̵���wV��"T�*Au\��1pYǉ9E��"�ݶE��������z�=W�@�W���,_�T��yђ�y:g�T_21YfT���>�u�\u��m�`�cc�<�&<�*6�����a��g�ЛT�q�FM.�D�6��jp��;MJ���,�|Ө�����Iy��CS�g
U{y���w�)�A���u��A&��[;`LL���,��t��d�Tߓ�|�����qRx�&E*�N�0�Vds��"[�TRx����ʛ��Sj�k��-*�u),y���CYV8��{��c�	L6���k|���$�4��ήC�9��9�/�Wɪ�4������o���{e�����@[uq�-�EU3o[B)����|�ј
�m=�a�)��m�EV�Qk�<�}��O� �"�X�%�_��ˎ��ͳn$���^g�/�<@Uuw�������[F���6�+%7ږ��(Ө���S�K���^v�5��.�w���H��b�mS���]��5���%�QTs3��m���R=uTR�i��~�'b�D�ׁe�Y����L��)ڡ�ЬJ��RR�Ι��	������>�^�ad��O��t����g�=�0}&�K����k��u����~��(�w,EU4Ž�4���W ��{;������8����ѡSP|�m<¦$�n�6�������<�K�\zf�Ϭ��޳�uN����w��Ѳ5O5���e��f܅���>������y~�uO��_�N������9X�񴰼0���>z���S�]�s!o�`�Bk���)Zc�'x�ƍ�:�')\ͳd	�ͻ,��(I<���H��d<�ǭ��Ә�f�I.Y��
�dD��J�Y���=f/g�KN�|�g! y��n쬍��Ƚ@���\�����w�?2\i[�|zAQ��9Y��}uF56Pf��l���2�c�q�QRK�{_��x�0� ݁/�0���]���S{�I z��f����.<��m��jj��։��k!Λo�N����1�gAx�΀㺻�ǣG�hj̵���C*��@;�ܠ�%{�,�i� �\g��?�5U/�,��#����:�������mq�/����G�),�ijH`)��[��g$� ����_��z��D����F0���H����a�f�=�a-A5Ed�	�����9��;Ab  ��m۠�,�N�`jT�D%���:���e���,ڲ3�`�/���<�hH3�F���:ǿ*!�(�to���GUx��n�`:�2���9�:��&h�����춢�z���X���� [タɾ��(5����zM/��g��
���}P�z�Kl�����T�I� �yb���l2�]��|���A�������3)��~�'r�՜��E��$z(�l
1���t0j�rS֛�ґ��/���:��Eh�R�G�Yz�2_�D&�\�;CƮP紤q�P���fk�6������^��ɇ߿d�4�ߗk���<��Ry>���"$�?��5�N|鿯�v�Yt���p�嫗���K+��]3U*O׏��bSֹ�&�!Q�GIFZ�d����^G��=f���������ޟ{�v��_P�߽��b��9]�`H7Ft{�ͧ0^��*L�s�����۶�I�>��$�������(�p�!��=�H����	�6�U�q!lD����F�Q���L�.?=�-7^rz�^T.e�I��=�.�B�]�=ʠ��5��C#v=��ڄ<��9�U]cnO�jK$~�����o�_����B��}�*�a�ݨ0#��J67�y�!�Ӌ6�|�e�.C�.<��������@�Y�˦�\T���)a)\�2����S�Mc]o��M=I�J�\��2����#D`|�47}����9w{MX�8Ȼ���}{����Du\[�y�y�m��*�2�����^)u)%�w�ړ�[Qa}��t����ڎ׼�� ¯2�q-	i9(PJe@����'�!~
o�E��Y���z �j9�f�S\�=��%&���K�Y]�/2�$a�	̒_�.�
�����x�'~��m*9��`#-�ё& ��������߿3E&^w�JTzbݰ�ML�w] �g
Pj��!=k����g��2�z�ԙ��)h��&4ɍ zN�Tj2܆�	%w�\�mUR�
��p۹h0�ὥ�w�+��Z�� �r!<2QrQ�jC��p���~& �q��Zy,v�F��:k��?�j�����=�K�qO��~�Y����_#=Ϭ�W?��1��-���`�>~�3#zO1���\�2�� �:
��Ȉ�5l���Si�d�+W��M�>S&:�����ob/TPP��_��'�imD�ƴn�7�����T��8��������s������Z��[aR���t�q�φ�zj�I��ٓ\M���N�n����D�n � #�k�ɸ۳-Bk��l��Ҥ� �#�Ab�a5}��m�+�	]��Cx���l;��7p�~�����ӵ0�ކuMɹ^�k�����t�`�4��L�Z?��1vk�:�~kH���L�xf?�N���\�7���6"��+�� N n������E��5v��f����x�:@I�����EFpI�6wy)|ގ��}�w��j��g~΋�����>�Mua�{�YdH�#�������nE����o�9�l�h9���>DThw�c[U׉J��Մ�EFC�)���,ah��{��e���)�k��\Gj[�?{�~��p���B\[,�ox���Ǉ1��u��K��6�_?�ݶ�Z�6{
�Xb�0���tlX��i�:/^�0$�@�Os�>"�C��%�-���j7�Z��T	��E�D*S���\@&2`���3��|P	��q��h1!�	�R�=I��8��߀�d���2�{�H��⎈�ެ��2C��� �º�
�\d^���Xn����|�Q���ŸBHd_I��k�k.�x�}ˌ��-�h���U��x���G����^*���;/N��2O�g�9+���𪖆j[c�Qᥳ����S�j�#61J�?4��9|�Cl�S���	��'��z5��k�������Qׁ�뷭����gHf�����rx~���xi3�$lR<�F�	>�yB�2�ʢ.�@l#"���ʺ遂��2�Q]Ԕ�<R��7����c��S҉����S�uR{�)x��QJ�I5_l�/A`�n�y��E�j��k#k�ƴUx�8(�~����N�L:y�3/�!��.=�E���}����32/�g�Hޝ�m�Z�2�rc\)���ы����~�'Զ�%�6�Ѯ���g7��;��( �0�x`C����5�ľw���b�Ra���4�d� #����YE2���i�s���6�k������ݳg���>�_�w^���C��u, &b]>n������hS�ή���h*e��	*���	��A�`[7*+���}�����zzn�9�'eT�u������Fg�C��K0$U��<N�����	֙r��k�^�r"� �����k"���;���~�zޗ�h$�����q�ޤ�6�x��iv��h�v�����~�}�5K�� ��7	��d�it�j�ثطx�u�=��U�e����i/��B��8k5���G�7�F��6�^����$�\#Ֆ�fX���6ɤU𛡽Nؔ|�z�����#@@��:���i��n#Y�~��O�`�Ïߗ��?��cB h|>�?=�0�0�777�q�GIVGI��B	
��x�*6��z}=d�.���!<ٛ�ߕ��D�}����DS|aY���;���w��tvR�1c8�3�q׽�F�r�EN����g'{/�+�wN�i�r#5˲��Ն^}U��BC�WLM��+�~�N5�P��E���f���v�ۭ��t@����h��H�n��F!���Cքc�]F���)ڜ%0��~Jc�ؽ�6S&�����WC��+�����rv�����6�밐�)3�M��w�N�X2
�yh�E��Ӿ�0\ڲw�'(��8����E��0��=`�T꬧<�ө����7߼1�{�N����l��,�����!�B��MW����RaǙ�O�[g��,��6�+O���3K��L2��P�o�H�V��F�q/�*>�>�¥/"쒘N�Ŋk�*W��	���I!6����%���)<4�C������k$�,���w�J<����ь�鴷�%������wc�����	���-���,� _6��ڍ��ڪq���R8�a�=-�z0İ1����G���D�B�V^��p���]���g[ǯ�R[�p�u�|����ՑD��a��x���i�kFG���B���WzU��[ٸ��D��]�n\V<��{	��Rm���lLl�)�#2���Zu�K��������*: �Ǭ[pϋx�҇`��<x���Ѫ�umŪ1�X�GI���C[m�-F�Y����~����Z����UKl���`�K����_~|ޘn&��7��!u<G�I�|<F�H��j�n�%q��i�S��R������l�א�F������x:F�a.ZH)B{�,������o*+�0Xʶ��=I�<O��?V�&�������������?0��TyHV�HKF�s��?���~.�%��.��nO~˘
.�gD��.{�[c�}6��˦����w��:��Z?�-{��3���x_0��0��#x��޿3�K��`늻���e�N	<h
�
|w���q����Z�N��]NB�fztE����|��&��S�M�T3���'��CH*�#��&�0�L���S��ĺ�G�L+ `����0J�:H'�5��gc�Y������_�m��K"�l�s��5�z��%�V|��wM��+���襂5.O��ZR2���QkV����M?�?kH9���	�|p$��K�g�9Jʨ߄���'M�ݝ��AkI�!��в��JZ�!&��W<D�<����vv-0��;�J۾�a����j_\T�Uow<�$~�����(
����W�\4�OL@�z�"-Vi�I�eIuv���|ҧ�����i�~iq��m�s5�j�=VM4P�Ҿ�\��Q�YT��g:�yȃ!o�k���
�y��[�&���a��㽵��|i�#�v�@$��ʏ�+C��_�>M���?���[����D��S�Ph��q�}4��L��H�@������]�h��j��k�T��x�&��F��
��+���+�z[�D�ΨOԣ���{B,�E�S��B�m)5�=�{�/>����C���({&<���
z �%�ǣ֊s���|���_V6[h/l�	��8+��W2@ p�(iX�q�e�I��{�+7�G"<g|���ntU�{�����+xv��xdHS�x��Ű�X�a��P`�]E�z��N%�b��ՅNA������WqA�'�p-<Ykr���^m�8��]�x{2�2���x~��8���<�*i�;@�K���,%��k��¹Y��ģ$��;�T!��W��dּ�bg���v�l?��'"���}��	����%�ty���9F���.�5%� �O��&	VOz�F�J���N}mbB��r���*�n��F�i>5���)���&�(3*m�'Ƒ��K�\�S���QF~ㄵ}�����]�ѽ<Gӈ-�l�v>^����{{/��T�@�G��F��!I�hB�a�N-u�4�M~������m��<cH=y�y��� �	�,�a�I	'�H)�
��Y����8����;��kh�ɺi�$߄A���\8$q0��}��ou��?�P��O��X�� ���io*�mk�,��{[/��\�>�ԑ)0���:a���`-�����j+l!���1����}W�X���&��Z�z�2<�R-C%k�R�o9�©r��$�ԙ�O�1r!�uk:�/�c����j��Q9����?~��ĸ���>��C'1h���F7�C�eI|L��T���G�?��PQ�a���2p#ƥu�c�E;��jc��gi�+FI����u��$��1 �|�ڛ]�6/Fܻ�2ECΗ10~�(
�`��T�}�(��ꥺ��TSI�q?b-�ɅF\
��~q�e$��E�^K�	B�q�U�ᯚwQ0q!]���1�k����J��`z�7m�F�f��a�˕u���My!ie���n�H�m��.:�H$h����X \��.G���;V������)������B�}q@wMلL��5ǯ>酵 ��$�����'�FM����B��<�9}a	2�ܻr�2����@�� .��
W1�tro]���[���G�~פ��&y���!�q �]^q����b�}dI�6�,/`pzp�* B���|c����r:3��}�m��~}o�u7}4^�%��6��L#&���u����:ϴ�fJl���z�,��&�h�\�o2ۙ�e��6<�h��Oc�H�!a���!���ܰE��U�u��a�1��3�����@d5�d�ԇ��j�N���s���!��Q��	`�F?K)�{�&�_ّxY��@���Z�3�g��9��M�}��k���'��5���-�4��R�B�q��'��B����]}3�v����������=/^�*/_�`�����1�>��74hP�G��1Kltz�7~Z�{�!ԅ���t{�4��u���<'�5AL�K}�C�����fg���:{��PxX�'�pqC�!�H��Ґ>�w@9�o��,סni3X����.T�|�,(�IpN�0����c��zT�xU��m.H��~[4�CT��e��}���2K��a5պ�,!��,Y-���2ySA+�`��r9/�SX�y�U'�,O��?�����W�S�8&8[Sf�ü,�T��vC�gC�I���������z�1up��%>\���͕�vN�e��$�ޯI�y�돲���6�����|��Fa��7��L%�]�Ԙ�oݙ���ƞ	�&�W�.	�W���M�t&J}���7����po���2ʵQc�_��~�j�ƴ�W�2zҜl�Z��`c!Iȷ����s�kC<1�h��vOH�y���0t�G�νRS�V޽s`�@�Tk���<;�35����Ƶ�c�7��)\H�^�8��"�q��Ę��{��.��Zg[8U����Y]��U��_�����5[�:�b�V���A����ǹX�e9;�6�W^D��6�H8�-.��FK{x��0��a$^y��Ǹ��ޕ�>ءz�y\P����#��u�{e�^ǈ�θa�,�Y6�	��>j���a���l�jm��so
f482���:�I���$y�6V�'�sa ���]���y�FW�?[��S=���\�����������~oUf�G6[�Z.ꟄϬ�~���!�����Yu*�h��r�oy�dc��0�{�tB��+ê��-Z�p�+���4�_멖���:=RW㩫D��M���X��`����#4���)$W��fg���^E��
�6��=����ً7Jv8=+r�D�T�,��K*�*Aөj����~��u���wi��B�~ 	��z�[�[`���^�@��t O����e3�u��TF/cMf��:����V�$=�9�>S�A��i�ݷ���ܳjj���I�ѓ���6�I�hK���Ƅ!
4^�^�[&Z0v0� m�����u^'㪹����Q�`�p@�L %������nn�M��:U #�C�,���]Q��Mv��23�J��[#����Z��ֿw����K���*�bQ����2�|��}�*��}�=C�y}ݯ�k���,듪f��}/�={2���@�������o�i�uE��� @�r1|;�߬wG�g���qaT��V���N��+�q�S=�9�s��[ҵ׏�6�%�|储�+�N�m����8�V�<K�uR�)�l��m�8_�3#ƞL�s��wx[^�zm'�4e���Ι�e=��Lw�]��`Sb1՜��0ػ04š_�"�b9��2�SQ����ߛ�ђ�xK����g��K�W�(�Kũ&CW��6k�b��mxV�ѸAgJ��O�ir�����_�x� �S�|�� }��˅�	�`'��N�^)�C�t�L�������׿��OѺT
�Z�#��SF�nm�1�%յhL�͉`�zt�|	�-i�E5��s2"���}���~�N$���cv�JcOyE�ED���?���$�l���8�^�p��d��`�`�T��'���?��V�v��d<�������h�[Mp�I[�}펵!����*#;,���D�"�T����'M����u!2�6���4��E��{�Gy�����I�))P�;���>�x�ڄ�)}�))aצ*/sw�0�y�3d���m��3�h��@9�t*�|�@�/k���@,(7�~_a��H�:ƺ��B��'6��ݧ�l��dz+�"��gI[��ڂ^����7N��y��c��4������B6����M]����ˁUsF���v��Ѥ�=C�ٰ0�
W����8 ��9����Eb�a54�}����s�XcqN�:�,����a�	��:�2�0����Z;77�9[�+��?E�z�P�\�
�K�5h��OV?Ǧ�]z�W!}R�+���8
1�l�������6����_�Ay1���(���+
��I9M�Q���A ���������oj<��{��lq�H)[�}�x��{ͥ���Mh߇��p��@��ZKM�Ab��a[��(�"��$F�p��nq�Z{1)�������h-��!�㞛�~v-�_�ק%W�J�C����;p#����#�(k�;�7�yYͱ�ǀPw�BU��L?Oo�m��,|}�<9Ί �"2�g_\�#P#��'�t�dEދ��p�R��0�d�����V����3���Ɍ��j���:T:vˤ�h$N�hۨ+��C�g�s�0�ҧd��Us�s����i��c�j�W��T �zx�{�j��:��0/J]xh�V���`7X��v5��*r�=���=l��bks�.�������A�c�غ�P+�1����4���C'�O<���=���1�Z�'7WS%�,ٺ�"V+lD��&�l|o���b����ԅ�I��*cx5��fj9Ep]��;:�eb�S}yK���V��۷���z�1AH-��~^���z�l߮��#Z#?�x�0H���ץH�s99�S�v�(>^�mj�<�q9��Me)_�EI��?%
��	)z��;�'��Vwb��	���t&֔�S_ͯU��k����C�iT��{����)����򾖪�o`��bX�E�zz뺤;ǌ�8T����S�0�%��B��4~){�6��H�Ń�?%�|�1JO��(�［��fkƗ^�����=��~����N!I&H ��x�U���f������O�Y�tJӃ��_*�<����� m4�D�ǟ�:5��/)K�z��n�o��'�� 6Bx�Lj�������2���6�r|�<�u������U^"���Bo����'�莆��*�0�5�Æ|L�bd	e&mz����y*iHc��4��sat�s�3���E�-;�*��k��5���,8�h��;����d�_�_�P��~���{��|�͛��Ո~�z�߽�f5�k�#���%/W���yU���1���桰c��p�d�^S,�X�i�*�{�ƣ/^
WjM
;��KTN��qq'�Y((>����g;���*�{XXC[�u���J-���%^�CB���*n`c�-�L%�����
����z�P�!�<R�-�sÈ���z��S����#H=��V����灯�m�|;�V�h��M}S<�&Xݙ��nnrI���.**��~�:C}�ϫ���?����𾝱h���?���'I��t�pn���Z�5V%�;�R�a9��l�c2���?�d	e~��/�xv��0/�~4�=P����9ߠ�$	_�
YB�<q;L��U��7��}[~��7�>-a����00'�7)�ū7���+3��6�/����7���
�M��[5�"g슀�*(ı�%<@?(п�]�m��F����Ê�W	�[�4[�`�Gn��#�󪽊M�TpM��<������O׻XvQ�𙱽m�@��Y�h��s���0�	��)�-��3��u��}�!�HN������fh��#��l��(~�rs����Eg�KTm��@��cS�7�}0��50o�#��x!eP	a�5Zb!~\k{�A�܉���3���gN��ԸmdG7Q_�
#o�ﯢ?����X� (|�#9qϬ2a����k�F���+�)(B7�����Ƀ�I>M�eS�l5�2C5$�(U��g��0�%�)x?BU,�l��/A	qҌ/
|o5�	���dg;��{�<���pn��@��9DeW�eo��ɓg�xhL�B�j&�R������4U�F��һ�߫��ՈvٗI"��>�@���b�v��u�+�<ކ-�1F�e0��}�6!�[��s�r�BfPD�Е�p������٫�nn_���!Ex�Ǳ�Ͱ,�}�ߌgeH7-�}-�&w�큃�do\<<���0��1�B�n�ub�/kh8S�z�0=�^�ڽe���n�a?Z�`<�Z�4o'&
�Sk��!����؂�lk��:�UvzNU��z`s�f�0����.��uYzz�翷�-*����!�m&�I��tj:�`�-�j
u7�g����U:�	iU��3��~E�]G��]=��־�
�TZQH_y�T�P,捌���U?�.��
��gi��t�T�MlmHEC"	�&&���N{���D�=Vs�C��Y_���v�ʫ����Pv�d���XI�z1���`q�z�g�Oمp�ทԨ>�~<�:l�:��'�F����ͬ�uM�ai\�d�S)�Dq�)8�x�`�z��<yޖ5���g���:f��	��K��V�|�{7��J�(���8���ɑ-�q�6&=���Oo?���J��I����<�j7߫x�γ�G$C���臜
(�z.}�m)��P������[� ����^ �'�(Z�P>�_���/�%zI��y����BScks��`��~۱5L�fr"��S�A�����p)���%v(hj�#��ΓWJΩ����5��h�Q%���^��B�j����W'����2zM���IUjj.d/-7�짱��i��r�(�����}�-K+!�#�z|��G��"Q����r����a���QO�L⚦�;<ѽg���-�G�N�V����S��5�+�=>ϸ��V�p܇a�R;�Lh�C�����n𺢍�] �����)_��\"�$�u��a�U�*�c�Њx�~/���W���p�Enc���{�)�0�]�]�*�������I����j	G��[�,{��K��D�����q؄��f�ø-����{�
���q�-9?�9�'�J�k�G����tj��"���ǣ;�h�~�$��a�8�?|�p7��=ڤù���|��5ح�^��ic �n�R&��P����>~�dk���g���h����(O^����4�KU��oڐ�Đ1�<?u�1h;\�O_����ԟ�GS�o"�%3�x�ˣ�I��i��~�¸��D6l��C�<�Y:)�6z-��R�v��WC�ܬ�~���Jg[�OOHS���H��5{]�x��-	���:mvUO#���u᠑!}��r�'�W��6�M��1G�7�_YH�k����M�Y+C����1�,	t�Н%ެL�6����d"o'��Xx����l�O�0ɑF_�����]�`˒����[�1��w^5t|���F�N%g7V�3n�]\����3������Õ� 
`�EC�:�BƧ<�An����EA��L�P���7�q�@k$)HKZl�&yX۽�=`����0	���XԹ��9��}�.d;�ѽV��m�2�UkZf���K=IO�����x|֐jQ��U�o�:]�Le��+��ԍ�"pe�8��:Fj�������$G?�I�8�n��V��V����[�X֛��Ӟ�"$+���%n��@�fPu[􏶈���������Gx��|s �SEH�?x	_c<�I#�P���2]�T�q~Fx<���T�øš3���{I��lً�)}��N������6��i�f��v;zU���m�,4���S_"�SF�a��ɉ�VZ�zZw�Uc��VY�aW�d�Mbn�k��F��g��Q�C�C�x�7xH��1����r*lS���e�H���w��Q�4>�2K$Xk�Ѣ��:�*����Ō���p7�����w��h�<Z��Ǭޓ'G�	-�Z�[����՘밆���Y�嘱���Ko�����v�.��=��ߧD�`,U1���X���kS����:z�7���]D�G�ߒ�R� *���;�u.�<M�S4��:.�&1�a�U�ʙ���S��I�\H�8:���U+��z�B�e,� 3�a�R�ur��1�W�1���x���O����@�J��+:tpm�3>��TWd����YA�Ax#@�1�����A���U�T�eF�ZN��|k�%Յ��YRĿ����{���F�FzL�ǥ��5�扸���W׀n�����DJ�̧��@���{+�w�r�n�%�ߥ��P!jI���U���K��6�v�{<�~ps���7���-]�`��˭�z*9��^����J1�M��õu�>OA_b{`��3YǇ�z���t�~��mU+ڡ����^�W�b��L�g��rн���b^7��w�Вp���6j��Im%��|t��IqҺ�k3B�"�
{��G����hb9K�7+}��<�GZ ���VGk����v%[���Ґ>�MS�c�[�M��bbY�Kc��E�-��h��I\U����p�N��F��BY*��;�(Hn^h�#���1�N�����3�xH����P��\�KQ3T%ImM�"
��?�!m���\փ���[dT׹}%�ߵ�!�R�Fo'q�h�#��n0�[3o��kO��c��o$�V��٣A,�t�ħ�,϶��#Bz7�%<����1�41�zZ�,��.��a��%����dK��١��I0���ς�/��&A�<^`���}]��ɬ��z��#;3�Q[g�%�B���rI�Q�?�&��H���(.>�w�5���ZAd�%K�gF���=�Ti�Y��.V���hI-�����B/w�=Rwȼ��?��E��Y7Xx��P�	PZe_Kt��D}�i����U�(D�gb�aR��A��3ި�Ɂ�&�o�������=;��v�<�L�R�%�#��mSxN��ncd�qS<q�y|!�r-�?|�
��R�BHxt�Ulʳe�3�ә��dۚ�):�ȓ�$M[��a|�ε�RL�C����˹�� �e�!�2��^�Ņͩe�]D۰0���M��?סE����W�5B!�/J�F��S[�+�-n_��x�H��Ŋ�J�^#�}�0l��Z�D�!���6�mb���#(�g��KR�z/>��G<ؖ����1 ���z�;�j|�a8s��g�m����KU�X�/Z�M�}Œ�h��P׬��Ɠ�S�A<,Ό�=	�(�&`��iCpO�@����â��<97�q���4O����CKDrqp�y��#aH�p��՞NxK�'O<�� �[x?;݈YA�p�ԇ!�\!��$8'VIN'i6(EX��&��5Ga�E��ﱘnt{k+94��#u[%�'���&X��<�a���mTZ�C� ��=����c=[o}Q�q`/I�^�#m������AE!��O^���}L��s�-2�&p�y-�q�guk�D,���qL�.�<Ѧ,�	��Y_�j��7��v̓�7T�<`Fu _�1�4֣i�5������L���+z2G$���M�9�D8ӷ%��R%:JR�k����Uy�vJ�~#�S�z����j>y5\�D]+\/��p�%��G��ݝ�	�-�v�EL��P:9˽��K

����M�`�=�FtF����AuC��vgǋa�ޗc�:l)�9�ʃ�rB5\+;~G���L��x�B�.W������k�0�?���о^<����K��5�&	���0�S�N�BY�pwwon=x���AR��Çμ�RDG΁%���]mW�*Rk�߽3�Gx1�>����w�h!T��xd�|�zM��^X)�+���w�ɯ�Ŏ1�h�p�_Q�)?;���#�K)YC��T'!70l��Sk F%Ų�Q9i��X�}�3"y�A)�8&�"q��Z�|��[X��JO҈ձ\���!��;���kg@�ˤ�l�f��¸��0�:�>���$<rZ�)	�f�Ή��W�zZ�u�\Q§���4�Ȉ�q(m9�5�����Xs�&~��U<#�Ak�� �7yѮ�e��f�VF��f�A���
�F0-:�a����@w�P5�Q_�e�O���h��9�=U�G7�5�b
g��L��,��z��c�Ԕ<yĥڷfG�ߗ�JnV����oF�ia�����_���K��*Eo�$�:T����M�ӳ_{�ɸ	������XH{�P�Q/�K��{��?:�������877�P0� ��F#��bg����Gv!�{��ޅD���AaD���k=����@�WtIˉv��X���i^8��g���l;*F�_�l�V3d��ʛ0v���.�k��P��M+�H*� ��w����TF���+`p//_������8 ѿ��_����:%<"X"�Fp�8�������3zrI�yY��<2�϶BCu�%�����!�|�%JK9�s�-&�������sd��{�0��C{$?aws@Q�1P��pD;���ߟ��<-����V7�Vy�l�wrQ�U����}�zDI�B������]E����{V���L.����G=1�AT?c�d��١�?��˥��"���c%�n����:�{d��Y)<�R��(�~�F�l�u�h�8��V���4�tl�=E,�gc���ΛgY��XX�I<�N��`�����7o߮^�k�p��G�c�#��1�AV�����G���7�"��Q��II�=x�Yc\?����<A���K�����c�i�nd�x�ך>�+Z��ٔ(����!��^eL��Z��4���1k����!����`j@�fLCX%����������~��{�P9��r�޹���߰Ė!����SON�W+�	��,9Zs3��*ˌ�^�y�ۦ���:�:PT696p�7m|.�O&�|��2W>>���v �M���D��R� [���d�� $u`a�\�Q�����3�����jp�����X����,����u6�?qo�`�q$	F�* E�%�L�η�����B���֪%$�:ޕ���f� ��mi�u�
�ޑ��nnfW�$D����>Ӵ�6�_���3ez�>H�8$c�)��qmV�Z��Su{B@4�6���RJ3��d��usV�5 X��z��R�[�!����G<~�G�/X��W��u�39�����dAU��s0Mio"�8����3/b�����t� ��3�0�ҧ���;rG�-N<�#n����\���7���~�C,�S"%ā���?���ca"�ÿ!x���1(��<壖yC*��C�M[��ΫZfk�����<�r4A3�������7��F% ����ِ��3�r� ��R�����;�Ϡی@��o�-�}��5#�_<���O�}����������Ⱥ��}A�(�vk�n����<�Iu��,j.�J����L��z� �~~ޘ2_�VXq�o+��\�MW9&,�Ƙ�ƿ}@[p@��mZ+�a��xL���ѡٶ>�]T/ʯ~�uz�Z�}�����g��!��I�
���B醜{v'�s'��A��q!�-f���X��&S>r�Ћ�X���j��2���PR�`�-�5�9�*�";���y�c�����<�Hۓ����D�j����&/�O��Hc�7i0'́vCߐ��B���4���v�.M�j��i/�-K�B�����
�<��Cn4"�s��m�~ ����\����?�Ok����+��S��T��� ��^3R@
������Vi�I���8T��_dg���x~>�hJ!�^�~]6�K�=���*��]L��F�}��5mO錴����h��=r�C��պp?��_���oH��2s����on�)�b=��S�|o޽��v��A=��a�3�`0�̋�_��h������Q�}Rz<G(�����16�h�aȒ�\e��p���>R<<w�k�]�8xD�s@B�G����V�mh^��{��6���#�Z����H����DSt�ƾ^����I�iӠ<Ƙ���GV�VFcr�l��qm��{���6=h�Ur:'�U���/�9����[4���LU&'�d��+˳Y#z6y��^�':����{dF�`�I,�~�?�$N}�04����?�H�J����1j>�?�;q�T�iF"*c<R�+Oާb����J�T;��(>�[�6�0`n�[eA(;��SՎ�X�U�ˎ)67���O��~Ɵ� �����9<n�4�&�A9(��E��Z9�x�������]ܧ��R{�,�&��z��q#�b���A�ԗ��h<̽x~�>]~����� @I��+lp�w��!����:�����c�]��l�����#�P)�x�N�$��J��4=ʹ��t�
?�U�z�d���L���2%���7�9�r��ߦ��kt��,�D	�]�H"G�P<J/df��(k�A�CA�W�|y���k��Dq\��Bk�Sd�A��8���!1/�=�1����6�]YVOd��I��"��r]2z���HXce��[�n-y���g����M�뻪�Bv��9�K6z��d��{	,��ڗ���3e�u6�E2W��NcTQ��&��'J��{^�����k�Ë����Vz�������=�#*bF�Z~�Ġ:�!�;����{�]�,����O�߿[3џ#���詍4_��H�#�m�R�T���n�OK3
°�Tg���b/��Mm�<ސnR�Qa�l"�XX��Mg5|z^s's�93?h�g�{�lIM	�rd��U�~��?ň��Ե�/�^�nDk�`���T;��∐/��������nt��Q
:���v�w\�3���)*Ԭ�}��{�W�$1�)$��b�Z�\���lc\�ZFnΛrA���Ȫ��[��2f��O�>����J>�m^�R������m]�E*�S6�kmȇ�2�Á���ټ���"�W@p�D�6ڤ�l �1���_|�5�X�{R,"�k;D����=��,�H<x���O����}v��THQ}7�i>tR��T��l�~(�j3�NzuqGM�Iy���l{
�N�ysǸ�J�>�x@�6/>���HւƆ��+}]d�o#�Ywy�ҲG�Bs��WkI����n�_���@�GRe6���9����"=s�v�i�r�5��A�h���k�S*>$�&LĔ�n�کn�P�\��Y�SZ�Ţ�����.�+)�23�t�����(7�8������O?�_?+��M���`f=!(�[��Ys_I��DY� fp�����4�"�9 ��L��pm�i��o6YJ7^2H�� �@���]�<E�34�2��:��$����q,�|� �Y��/����f�G���dS�IcX�7T�8�c�4	�-m/^��}���!+�h�3�q��p%B'�!�K��"�ĵ��7{����տH؁�"Kƃ�S�JY#�@�m^n@(;��e�<DH��Z�r���y�U��Ӈ3"�~�a��M5��kVJ��\�_�U�[���6�OR
�=;;�+�7�=���z#xj�Ԯ�R��!'�2΢̘����p-�����܇��>NN�]���De	-�Bi���6&�/__3ꩮ�j�M˥���-Wn/��^e�H}xG\��~���f���^�y�i���>�UDj���|d�#��uO���A��>�Qܟ�l%=��(����0ZFU����/�J!��g+���B����kX�p㹹��m��b��4��ī�p�����xnѷ��-�4��;����OB\nH�@�g[��d���~����:e��S�̹����!�A-ڷ��� �fveo�3ek��z's��3��)�JZ��ޖ��<�We�,�7ia����{Nՠ�7�/����'��M�i�4�U	v�!� �����x|H����8o7�k}�s�kԅ�'�v���� �C���\�gi���24�pq���7)Kکv�w����{B�����-��s�n�s�b1"�b�F*r�A���ިI��;6�M��@�Nϙ�:����ʘ�.2\�P�| 5�"�4j9�2�T�n
GY���mW�YAH)լ�n�	�I�,�}t�*�;��M�����{j������{�π&�N������q�O��12����=B�x�0�Tσ��^�0}�=jvl$�{=:>%��{]e��Sl�l0]S��k�����fecY�����61Q7i>�0H5�p���QRٱ��!���4���-�6����?�4�ޮk=L��sBi����.ޫ'��9�NM��c���{T�x�!�Y2֭�E��Ԟ����6�¥t2�>�}�{��r3��q����QS|(t]�R56b0��k�w���$����46��$x�"��0������@�ߜ�=��Y��"�DT�x�x���V�̦�S�9�
������z~�3�JPl���s�& #�N�(����;�N�h�Zr]�[M �ϻ>�(�;�}�V���w�:(�bL�ʙ��u"thăA�Yd����Ԕ�վ�'������4\�ƹ=_����n1Nd���6�&v��.x��&6�9�/փ�Z|���f����7kP���^���F#E8W��4��/C)����@�`&��������^�F$��L0��L����I�n��O�Z�T�]^�[n������7d��,�7���=�{	�&2�����ʩ�6x�P+ݤ;���8,4߼}0	g�sE����d|�v'M���m� �Pj�Y�Z�)������T�_�q�";��O8�"�����[[�����i��GA���*�g���n9�{�� �03 n��������c������{>���ށ4UH�(]�d�.� ���i�L�Q'���9ڃ�Mdf󼨣ΠlФdX� ���k�nx-}H�q� ��,�2�c��ڌ������.J���hl����7G3�xed�k��x�i������@�f���gE���1�GF*l��S��x힟��xT �Q�E�ꪂGTm�4aG
�ǟ�Ok�#�c��Ypx�k���W/��,ܦ&h��^7ҫ�)������/����Ӱ�&6��}Nv����f�Ζpwv�d ��Br����K~��G�Ƈ���W�E�����H<��e��f�i4>����);����c���Ư^
��E��E���i?������J�����	_��%f�[�_gg�tI	��#�;4�( �lo��25G��~������x-�.R2z��F� p�#��,��^�qP �?���7>{�|%jE+�L�"��F4�~�k��y�'#c�y����׏�bK����F9N2�9(	���)�j��p'�P��\z��J�\m�,<�CX�<�[>>�bz�C������v�W�� ~��.�lnY�x����_D����W�رP5��+l�H����M��q,f��,�ܑ[vV�WX��Q���  ��IDAT�j\A��4�އ���Ɋ�e��N*�^�:SL(���%�C�����놎 �n����Q���b�g����(-���Y�?c@۰!�S���������*�����t�qܬ��2ޛ�A�t��=�Y8��Iy�RX�2� ֖��G��#�����Z��<�>��sj�FB�Q�acX���5#��6L����Z:IUT(�x�Y;uW0q�l2�a�9�X��0ݒ�~�b������B�lKX۸gw��b�G��w���� ;�z!%�=28崊�[&2���H^��?��u��y�?�?��7�H�\��d�X@rd܉�*�q��2Iź&C��S�t5��s���ٵ�iP�'�n�M�A�9��dx���t&�]�`d��F�nr��Rg���� ��iP�"�̬йMdȝ��b�b1ὁC&(��S7�pQɢL,��nt-�hL1}�A����_)KJ8I�Y���yfv��o�	���@�>�6�cV�ҩL�'*��k��d��ë�laa�y�QC3Ts��p���娍'�	B�iʱ#��+@̀k�C�R��ɕ:�'���޺q�+���& J�	D�=�,{^+�=�����5�=��j2Ξ�R+~����-2���JG�F:<`�<��������{˹X��:���x�JSA�w�6�̾�h���ޮ���@�0�A���y� �HX���x��l���2[4�}��^�W�f#G�f"�L�ȶ0A"����IO�� Ð��!�H>&�S#<AK�.	��iq��=��zʳ{�Ѝ�\OW�)\��V�r�י�e�����]e�I%q>^�,����r���A$|wB�����h '�cR\�  {J�ܼ޺�<a���%���鋛|7�%>˕�Xt�Jd���үsP�:|5L���@�cd�S�)v�{�`H�Sj>�3}�Դ�_����}i�IT����	��@�>�lO|��͛7�0�� (�I\Vttt�)�u��pREBJU,#��9
:yQ�H��	i��yI�f�,��f\�\0�1���I���=��׍���w�Z2��������_��:�D9��%��c��0[��X,1�����x悢�����cU�^��2\�r���=O��Ll^�N"���fʦo�����̠�{�f�� |�7�s�P�IN�fu�E��̓<fUT�G;/�E�q-ll�����G��Á����o�M����ʾE��k�T���������3X�TwyEC黪p��V�)��1������N%;��B����	l�H�T=Mq����L��u!�y�:���<4��9Kݍ:��蒖EEE�~��E*���I���+PR`.t�q@0�d�J\ǀ:��̦���r��55�bZG�����ΨF��/���#< �����4�JƲ�.�-�Pd���Ȯ^3�wo)t�
 &� F�X*�Fd��׬�L.AZ/Q�u6P`��N)v����sZ-��c�m\����-���9�2L�qe�&�A#���ƳUH`�3�S���F�Ȓ�5<P�ny��L���n��_��:F����H�@6�7o�C�m@Ev���� �Uȧh<t���2j�s:��u�|МT&S�,g($*Ӄ#����.��p<���xh���<e���o�7VM���k5*�����!���5�����1���L�����Xz���61'O��_�;���S���̮&��N�^��@��$p�)�inZ����?//��9G6��	CZ9��������kje��0h�5f�Kn�]\������eE�4/^�����8U�4��ct��5�i���|����=��̑m>�'��=Ć��).R� C��Uû����pi����-ltE�Ҹ�!;�|P^�麉�E��8<��� �v��y?@� �TI�˒S�*5�Tv�+�M�
�q���^Җ:e��v�ll�f9��8�{�#�s�y�6]t��i���9�wg1�j���e�of6V��b�����!�1y��������D�C�v~����;���ohrML�L�%��G�<������/)?���z���l��'vr����sv�c̎��`=�u��0����qD�;Fs*+���ދ�CW�I������{ �Un1^�Y4Ҟ%4����vIw�s�q�l߃$i��TT��1�����%��U0mzBei�W���]���Y �򣒃�Y�t��TA���e�Y�,�m��9ƣ���v����9�#Q�pOO��>�^�R*O���i <7��.�Z�#���u���?�����G�Z��y��D���n�AN\��B�_<Oo��u��������)3u��~<t����pٜU�^B����[�.#�B�v���-7@:}^�����ݞ��δ�|&tXq���g]����5�.��΢��}���C܊�n�܈T�B��y*�����8��2=iNW����=x�?���v���R�|�EzM@ ����N������t#͎ME{LZZ׊�n�!@�ݰ��n�W/"���a���^��'��=�=9-G��$��)��,��|i����(�p��_��)l��Ie�N׌G��1="����dS\Ĩ@�H��o����߱�T�Wѐ+�C'?��0�������῀Q �J,]�"Z�/Q1`�R�!� ~H�gڮ�磃�/S�������{���δ����n6iO�QX��>'z�u��@270�} �C�$����(U&�Aa�G���$�c��͌4��m=OD��*���S� d" ���¥���w�}�"n"�Nx�?���j�[6�v�������ᵂ�h -(P2ƍ������1�mf�Sz[�.3�As�4�2��ͨ t�XB�0]� �d�;�ht�� W�?с��N�J���K�A�seQ,��k}��!��\x�UX/�ی@��mN�%�[q�Dr�{�(��D�?����T��D��ξK��<�!���ᷱ>�p��e]�U���ݻx��9���md�w�M$:^\_�}�bx6��ț������F���Z�>��;q��q>�]_3�ب�z)2�g��l�7�B�'M�6zf�gcȄ����DD�14W�BS���1M	FҴ���e8���
� ׆����g-Ł���5��H|��E��gbq�O�Y��/g��J�ַ�`
�����ũ@��j�E��:����j��l�4��倬I���g�	�IX��'66&2�m������{A�;,�v��
�������'M3�i��ٙ��(�PN�T�	�l�4��͛M,�ql�M�>pj�̃����5�.9�&p���΋� n�QV.�m��O�w�]R��{bgL9���[�ݖh�LC��������Le��0]_�aNp��
/����i�f�e�g,��4޻�nyz�z	�*��%�2siJzu�u��^S�ȸ�G���IB�$U�%�3.x����=�)Ԡ{�aX���0\�j�{�iQ	�w٬��w��~���Zd����oޕ�ݻ8���Տ�K?�����0�ǚ$��u���U��.eV��^=�3��5����<���:�������t%��J�ٛ$�8��,����s���Q��YKa����H����VR���5�<}�0�$�yw��7>�����O�0Dn��X��,nT(k<����rgӘƬ�4�_��MsS�,����ѿp����o�$bI��4#��.�PV�>�CZD�h����t��l�޽{_ǎt���6[�"�_��3�!�'F\��<FF�&��.���Pe����`m<�O�M(��g}V�dWz�ᘐ��\�l��t!C+X��/}�˹�"�w֜�P��4����Am��f�v�G���57���5��x�,�3=f�Z����+ �\7��þ>�g�lL�`l��P4����?����6�LLn�9�N�1"�$�� ��K0;�-F���x �	���0�9��M�C��a�A@CdȌAg������r�vڧ��d�K�䢝1��"�dr��؇�ˬ��Ԇ�BR�W�0���^l�����x�
ѕ��v�	�,�#\��q�A����4�)s�w�}�����F�q��"��v�������^������*��Β� �B8����E�e8�q@ ~��u����ct:�'~� �����s��N���!�Í��{k Mw ͕�@��cd�n�-�r������u�
���8;�8cB&�{z%2��I���Gn�x�:^�מ�ާ���E��Ѹ����3�������x�$V'���y��c-�Z�.����Q��6+����7�>$���웛8�Lg�'-�;}�%��K�S}ςr�"���J���Sx��]|�]��P����)�KxP�`�����p�1u��l���O�
��1��%G�<�5мz�����&^� ;;{��=�"ϟ��fS1�9o���Y@���˸��a7��rl�4U��O��ʊ@��e��C4./�Ĩ�y� �iۦZ��w<S�٧2�Hz6��Jj�:#�z:���{����G<~1����gU�J��y����
�>3T�j�,��z؛�Ƚ�=.ǘ�0�cVOu���Cuֱ��ٜy�5#�Uٔ�8�)Y��9]R�L����|�4�UB\t���)q�C�a�QUʧ���S�¨�}r�X�ȷ�>�@�j���P�H�T�4vh�PH5�Qj�1)>��JF���r�,Kds��4����bZ�N��(�;,M��< 7�m�I%d~��_�o��Ɯ��<�\��Z�����l��Ag3�)�h}����aVs
;��Q�T�C��Qg?���^r�
�P�B@o�9�Pv�!%~��C����I�C�ּg��z�hT^Z��$����&���@w��8(X(�;���7$v�*�%�sY�eLU�M�n/�_�u��E�k��pS*�(����~N���(���^��H����繦=y�l;�5t�ٜ˘�n7J�S�i�ɥB��|>�<��Ct�7����C��4[J�y¿��㫤� (��a[l64�Ѩs��9dN7���?r��ɖ�"[ec�PKב�K_��(bQ�ݦ\0�J)�I�L�����NA�pCe��y�'����%;5J&�8��ѭ0K=�Z�ob[E��P��(�����)�C�7|(٫�dj�t�.v�5�j=�c�_�j|~���ˀ{yO��30�[�ۮU�^>�PKD�/����eo���/��O6� � �x-�����B�_\c)m�4�Nj�D��իxo_}�yK���Z��rj-�/m\�B���F��1/u�iW����l��2xnwヰ���ݨu���FP)K3]�(�euQ�b��"�ʱԁ��,��8�zS�W��(�>��oo�z:��0yϢ��=d��L�ޏJ��0��[��F���DU�����������<[��&�%X&��s�Hm�՛�R� ����f-����#��w�%�mf����`p����F��w��3�m��/6b>��_�Fq����i�,\�r�
m����9�{c#+]εy�����K�P������s�A).�exaFCO��9;�x0�1�8�F7���szeE�#�l�q��Z�J�1wn�����M`�+\�S.i��k�G���������#���U�ڂ.�GIl׎a̦��+t�] �0�I0 ���d��	RB/Ѵ�B-�!��Ϯ�gt�c=?�:�������X�Vv�o�^{!�8Yf�H�'L൙�r�`Ȯ\���L�}�w�s�Ჾ&��zB�0�e��ե6�t�XQ��H�N�aB��%�Y���s�{�`�T܋���1�\��>J?o��g��_��j��ZB�\�i��{U����Ѽa��>�{�1�'4�g���|N;$�2>gdU�s.Ve`#��2c%�Z��a�%��\S�����7��ￏ1�(�r�[3�_46y
��4}]0B���>=A���ӳ�s-�Z���3�N�����aހπ{��@6�+��/�uV��R6p(��]������|?��2�*��ޠ�,���3�G��of��~U��IHA7��}���bd�'�X��(��p�;+�>iu5(��fD�7]����m��Qy3����=�������c/K
VU'x~�x�'f����嬩�;5˶�����G�:{�9���O�t0+����l��Q)��1
���t�q��G��s�N�S�A��B��%2f^@c[�3jk������F�P��e���{��{��QSh�X�����{������2�~e UF�~�ϊF���SV��HB�a��H|B��ף���a��R��1��w��t��m�T��S�ĝK��(�������RBͱ_B�B:5A���Ҙ�&7!o0��}N����Q�\��#����GuB�Pلr�E�g��%�C��8�B�s9�ij%�&~?��͔�c����z�b�Pe�<�<��TY�L������3&8��H4G�Sږ��Ĭmּ"��S_����1�|^|E��cx�yFv�q�w�cq�[R|��,� ��A�eZ�3*��hpr� X����c��=�mTmc%�p�5���������x�8\��#��# ߼�5qWvp�:��`�%#�J:��#.H� _(��a�e�{䁊;5��_v0D�nB�}��(w�=fۣ�ݔ�{r~����8\pPڐ�b��<i���X>N�\e9cpUCx+����9�me(�Q�p�;��t��:�u�r�ZV����c]&-��ԾϿ�1~.��#���l����A8-Ё�ۘ'�7SNs!?��%g:��s}J0���tȠ��6[�����R�TJ�����1/(�VU��S6d�
쫗H�-��d�I�8M(Qʳj����1nX-h,��1,�y�*0·�徳����o�#��]�FaZqO�H�����W)�c�������r�#tE���MP�ύ;�y�ҁJ��Ԕ�݆��5`v��4������T�и���$4�n�v��/Bݑ�q��UUZ���b�ڼ�ݜ\J��&��=�x�<:����x�~�ז�����LX�g�ꐥT�7�԰.�׽gO4�&Py��Ô��N=���}b��	�����nH�C&VE���z�׳��OB?�G:@� ?iƔa�pӇ���ZL��� ��*@e_A��TL�F)7e�T�'�NQ}!	��W�������8��"�MiL-��1�tQ������˥�UFZ��O�!��kd����b����垀�nwN�;�]��_���]d����*>
�r�\5���V��� ?H�N\�F�z;6�塵�(�l(�σ#�Hi�6E���-��-�#>o�q� �	v�E(G@�w��&�,j�=i�Tjꮃ3wf��m�%�NM0�����|%�p/��qp��%�������e�Ǎf����
)c�P 9P��js�Q�)j��%�S4q�ި��8���j��8d<6`眗��
�>�A�n�ڇ`Vȋ���L�m����&��7(OXs���(#?�����\p6M�A2�J������r�=wG��!�]�b2�� ޳M?��>W�XBi���Y�L� ��x09�0C�DNgһ�����!�7~�Y|с�=�=�,y9�2
*$9�!]�S����:�szC@bK��W�qV�H��
-��B���pdF��w�	�����k�ee�/��RO�y��V�:����x���M�bFK.�%7N8���� �XZ��0TR5���{m�Pf��?u�!p��"@�{�K�P�����h]q�,a#����3Iܱˎ:��o�(v��ZP6��j�b�4���0>�B���Xz�(n(�3#�n�����@66)l�'�����rB/jf�MCI���0\�Ѻ��t|I,�jQx�5�L��Z�u{I��t9�D~����t�4]�q����[v;�!e�Y׉6�8o���3)a&�#��_J�����=6����q���i"�i;^���]�3�����Urͮ�����CE$u
Kxm!j���BH�א���$�e{��i���ʄ���
a��;V7���J|�~��E}�/S�ZN$���E�Z�h�^s���>隆��8��o_
���h�$>ϗL���	5�X��p�J���Ѡ��-e1d �D��|�2�0���!�	�Y*ۘ��r4��BX�G��?_�_����E��!�3�<S��?�zU��(?��Ͻ	��P�!L�"�gGXM,���u���Ը����� r��������(s��zf�t&h_#8t=e��m�OFz_��D����W�	��F�Pcj�G~1���7�ƃ֤*#���r\��?��)1�]u��1ѝ�N\>��|ݲ�ܘrhc�b�Y��S��@��iN�I��	q�"31�]`uU)V��#������c�}�˄Y3�N�΂�#v��B�?����Db� (:Ճ�E�\L.�&0$�w�%-'6��jz�]�%e���+ߚ�C±�6��-�um�罕)�������<WM��x���3A
��eɑ!�B:O՗8̱gK�y��)�%���%wG�������|bZr�3м����%ٔ�Bt+E���qX��F��Ŝ۴��B
�c(��7"c;�?��z���Q�韙�t���mb�������������O���Wm[�j%��0�gR�m�M�X]��42«��
��>�9~�r��N�:�����������x8�Āc���Tp!�g+�rB�%�w�l��R��R:�BL��a��U�O���Lل�Bi�Lk/���O�!Fq	tIg�����MY"5Jc�����]��a��廏�1���ȶ1Y�-HP>�j�I
ZM���4�5t%�w}O�AI��ˠ��4�1��i��ω�{<�
�,)�<��b���+]�$Ss��l�Z��^�� �i�a���a���.q�U�8	 �x����Շ�,����ZJ�7q`��J���(�փ��o�%���{�@N�T$7�������|^�y!;�6&/9a��p������ns��BQVGu����g��Z�/П���S�|��l�'��Ǽ�Y́o��[�9$CdFzmc��,�MdtpQ���sm /������s*��De��!�x2?[��Q����_԰����됐��]W�J9���Va�s����g��8Qj\�
M��W?����bX�ǂ���#�ۧC��uh$�/�{h���]��54�Y����9!�g��.0�^N��
��E&wr��%���l<���ku�=�)�;��.Sy�J�<CC4�,�9����ơZ����C�ČRC�vG3����c�[�şqoBEt���A�b����p
Afe!Ǣk�(7,��تa�3��Rg�[���Dȧw(��w�N��͕�^k]!�ڿ�� ��!(����:�`#f��}�ǚ�ʏ�gE�J��,�7�����m�݄�������y�0|�V|`������)ب\���x}��K���Z�c�Q��"�#�;񍱗<`��{�HkR�_yt��/�t�G��5�Yا�x���췴8I_,]���r��$U��L3Z���F�;NSv�q!�Q�l�����Y͟j����E�,E���D������˿�K���')*J�6�lO������&X�y� �GC	c��o��>�(`��؜1�qsT�rLuFˋĩl����)�܃�sQ��}����bea։�첝��v�� 6�~a�8r����r��F��������-�{����x�F$�`{��{|�>4��&O�"{��)ǛZ�.�{ġ ؘ4{�!lp��gNk���oU�k��I�KWK���tY�� `�����n�"�k��Q�{ś����x
fs�oD�ǃ㖗�4¸�g��P�օ��C�	�����z#�\մ��g:��{�]^��#���a���5Fx�i�Q�u��z���ě#�jz�{8<� �դTX���cr�}@_�3@
��Р�ܢ�J/��2qH縠b����}p����}5_����	��<�Z����MYr�D�/��Gi���EnB��3V�b??>xdk/�'��\���V~�8�D�Y�����p4���������% k�S7y��d9.�6@j �F�T5�O�� e����Mt���Q�Ar\l4�ؔ�pѱ�
���AM��0 �ѭ��(���mw[���V�O��	|Q�f�tq8�\zPM�\�WHk��i����N�6��ME6�k�.?6�[�s`����׈�͑�!��B����.�~�B�4��R���D-�J17�"�N�܉[������q�w��ۻ��N8H���=�|j m�|���:�_��9������ب�7F*,��ڢ ��{$
8t.�SAv�A��m��� �ݚ���eɃ߭��{v�L�0a�X����N6á�i9���1���"��Qm��^r���������k�~%�T,��7`��#�l������������s.i�]R$fO`�~���8xZ�:��U Ŭs�z���K�!���6��ޏ����o�G���F�/Α��+�ÿ�¤��m�t�V��}ē�r��`t��,�3;�$���D��ɕ��(SW� ��]WUD�J�E�O��|j���I�<��Cᢌ��Ǹ�^	Q<z�عJS��D��7�؂���wmv��.�ki���8ib%�<n�W��p���3i�i��j��s2cVaw|���|�����ׯ����C��;"-�u�k�Om�$�c*P����&����	�x�`��P𡑶�MvU	5^�W|�m)�����Q�L�g��G��*����y�؊�X!���4�{漮��!��/�7:\Nɚ���.tB)�<��멼}����w�����a��c���Dbw����\G�8��#(i�d��s�R6n�U�M���ʳd���s��Z�S�EG�~����H/��-{��koL����#7��}c����7j�I_M��f͝���p'i���#��K���E~�ˋ70o�N��3����� �}�@�m��S|w �"ri?�ޱ��4̼��:qxi*ۺ�Fe��x+z�e�u��R�}��yMR�8Иa��M}iT,6�%�sNvE�2�3��XI�JM��q�kz�~r��9,���I�:��33}ln4�����T����TM�cvq�5�	O��bTg?~N�Lx^d�}牭�ܤx1>�����p[L�Z���$�s��e6�U��7f9��q��Q7DL`ϟ���[� ��g���5��E#�Xg����r�Gq������2{<��h(��7�_�M֢�g��rZh<���Z��٘��5�zU�3�N#��X��Y�ƕn�JKW���BW��o��/�F���v�L�Z��_f���k����=8[1�[$�V�ܦ�	$KI�l�#4��P�ؽ(;�]ՉO1˽\�z�N)M,���C$��')���0�қ�t���4�c�C��M�F��1ƣ����AP��*Ӈ���T���ث�H����ϟT��i��[>٘}��y��,�/�G�	����w��֔G�g��P�������4[��AAC�a#f3!Lg
�R����do�]��Q�G_�&�d$�q+��Xw'݃�$�08�s5Pњ���D�E�7 �M}x�>>�|t�#K���DI�uWk��H��`7��S/Ϛ,̹�b�&���k�T���P���)���ߧ�?��Pi��W�ք)
gOzX����k_�KӨ=-$�ϵ82e���n	pM8��`A7�iߌ4��:�=��C6{��)�L ��߻�@�C"t��!�.�PCo������!ƢT6� �_6-�L���4;�CU�d ŉ��<�v;�9{ub��)O�HIk���"�C�,ߦʁc���y������e�N	)D��4<�@J��8�Q�z�����r�V?o���n��?�ø����(h�`,	>K��2(2P��� F~�N�i����+LR�B_��L�75ɳ��6�L=�����C���O)����N���U)���C����$�^�xx �4d���(G�pFGF�@
���f�C�Ӝ�p���u�R���eP��yJ�y�do�)�ǰ�[����^�Q.A��n�`�R��X�R�B���F�z�gk7��������E�Ǫ�������f@�����s�׿�i��瑀��ϣ`:r�H�&�A���.�=t�'1�ݡ�N�T	���i���jrժ\j�4���Q��Ժ��!����U�:�*�0��G�Z���9$v�2�)�5��u~�)�G����G��b0��iɧ�0'�R�ύd���F��9{"[��%3�&ѢM������ba��&�13dΌYRX�%�����2�X4C���8��1���:�����^~��+�Q��.�bq^�H��"1�����Y�Y��_~�K����ğA	�m��e��D�F�&3��b��K���pֺ����ׁ��L�`<ݥ�;�Q���LK!OtLΤ����)),-���3L�w"-�n�5�����f�SP���gKS�ݞ��+��9y��bc���=�/iE��Lb�jB�0<I�c��)5�x�����C�͖ţL�E��w�ςA�Q8��
��_eé Cu�L���f�v���A�l��;�4����0�9J��ի7���]��v��Y\9�Fօ�&B��#;�χB�ar��`�$hʎOnz�y6����)�yl��oX�WVF�͹�20	"ͅb�ɩ�.���^�����id�S&���5��At��������С)u]�58�<���i�����������ߟ�)�쥧tiB8V�h)KC	*�d�E�Zӣ�[�պ�*쀅��>6�Q��(7���L(}4���#�z����nD���	�}�"�T xo�X<�`/�%��*��({�u�(�9K����!Eg;LN6I���=��'e�������f����qU�%��@K��UD=[���w�&~��jr(�F�$B��(3r[ٍy=��j�209�6��t���nw�TI�,oa��`G?P������3�M0����=F����Q��̨ܔu6ۇ��p`�2iO{�%#`T�Q0$� �eA�+h�Bh��e�}��jK8(�,�<M	�:����F�HpY�1Cޕo��:G��w�:2	[��.�4���}��hw7U���,��'2�o
Z�R���=�t��Ǣ|����o �g0�M⢥\�@6�`�W�:e�i` \�"-��H�V���u#����Pv�K�T�Ð�Sz��E�C&�Ax��A�1(Rab�����Z�bEc���6�u�;̞�]ދy�O�(�H�q!Q��.�ٻ��#(>�{�.)��N�-���m�I�jfaC���cf�n�~fj��cc­�.�q����3�7}���Ӡ��H�91Zl<6�ٓ��o������2�,G�ɩ��a�X3��6��z���	�ݚ8���M�떪�G?K�1�q� �ߨ)�,��}`�E��r��Ma�?GJ�T�M,g�{$*c�w%I�����HI��1u\�#G3���ڬsG��>�~�f:��2O9t�Q�,T����˹�#Q�E��[�\ީ�|*��KdȋꦮƠE���o��{笌�J��L�B|i���xz%��_+9�7��N3v�6�°d$��W��ZA���6Ҕ��3h�@jl՚�O�@y4�%3RP�`�L5ԟ�ׂ��SZ��ցy�]P�"���e<�}�����8x�_�|Y^~�R�Y}�YF*h�����S�zr�J�����^H�5��\P��{Һƫƚ��:�F��6j��s��{;�.�x��:"x)�O��tH;1��aq����k&���&��{i��4¸-�)��R���������೸��LG+��(U�8Q!��I��ԽF`�D�&�B`��,hj�q<hz�e����{��̢�s�3�Ѹ�T����*��$n��YM>�Uͺ}�0k'�*]qM�M�����9f�Ul�6-8��%OA[�^��e$>�yrQҲ����6�9�i3z��$~S���?���ˀ�{}�T�F4}��:�r~�E���/��긶/C5%��>�)��4��a�;~n�"���Q���gb���X���dUyp���M�yH[��a@��`�pD0M��ha��~�L�$���\�7oh�w9�=`��nG�~�\<72��*��d�4��t�s���l��xz�vI�����S;ez�k�ZZՅ���U����&` Wu�4 ��d��^�L��;�GSi8#Y�OY��qh� �
&�w�ְ���Q���@���'�V�P��"e���ɝ���.S�}��S$�i_���ma���<��e���I�gM5�����q�OfdC��ݣ@�<
���8��+��6��PP@�M�����J&��(�Ϝ����A;~Gzx㎜gE��E-��;7�5��s��9X!���`���Њ���P���Xe��	t^�~��`\�(?`ܣHf�J��������@M�&���(��%f��c�T�\�_���i��$��|J��b+2eO�R׼tT�	�1&x����t�� ���E�.�Y0���X����1�;.~�O�I��1�tC&�����3@*?<�����a�N����E�n#J��6!��jp��5a�!e��еi���:����2mU�����X����в�E�_��h��uF���_}c��f��ݻ�A��{��dp���Wk�r4$�~n�z	���.4�E���L,0K2�pVc�u�~�������}#����z�02&�߽KF �iQ+A���.���y��9���� i�}���O�l��oބj�Y���e�/�����|�T�cT3��ٷ���'�9��:u��\oBz-^~3����ԭ��V��k�I"�^��HT=9C��$��jBWnA[��y��:��nX���]����Q����/=W�>8�h��yW�y>/<F�����������)�Kk�r2jb�������*6_y�5x�M� ��e�jM{5��䘾�-߮����F͎��4N����zc׭��.��{�9G0%�T���/�L4��	����N9.�A4n�h/Tނ Η%J��Z]�8��C$���T.;ϙ��O�cf�X�W�eq�s�l���I�;�	�M��:[����{�����~-0�x��AP�j]�_��}͊������s��gr
��RC�1�(�ޒ�d������k�]sR�T-�u*���!�C���zf��ob���Q����&v�����Y��~�J���V��ր�xV��l�O�p��l���`
��hT��I�!p�B�|=����ൢ�h�?��<`'8��/�������
=��<�-x �O,�dӗ�ɣG�)�W�P2]R�Ŧy��yHG��O����!9D���"��T��ap����t�_�P���´q)�,���,U" ��^���S5F�dH��{��b��^W�ѶYlĢyN�)������b	5>���cӓ�ڟ	�G�6�\�	���b���<,�ƴ��]J�d�E�>2?�/&�#��	���e⡎-n ������D�v�n��X�c�N|?�8�����Nޘ>z	�v\�
��;�krΠ��vѥFP��B�rXb���C6"*��K�6O�5��*��ꌶ&"K��gͤ!.��F�-���8U^>{I�����0y/�w`����3���my*��k��yX�.��U]$L����hY�y�$��1��4���b������ߝi�����%�Fa��o����B۟42��9��>�kd�5�	��2�sJ�Sp	튏����VyE��(cܰ�M��(�Ү��(�������KR�ĩšV���N�l��9�����kD��ֿ��`̭�4d1����#��\f��M�8��Q陮
��93�(�������lr�%H������<�.��?tE�8�}��i���icȦeD���̹�~��ۯ�����^d���u�tW����5�h[��U���`� ����St�O������oٵ7vbɰ(���$ۄ`�Y� �eh^�'�޳��;n>6~N5��l`a�ൠ�ƅ����p���8ت_0��y+��bd��u�F��Nh�(Wy�E�-nt��iקf�x��6T:Dm��Fd�oww!��q�q-��Π��}A����OGL/�YDq2�<l��޼~CK@2��~�Ҙ�Q��W?{٤@ ��N���SX5��"34_e7P)�}��Uu��M�z�Aݰ$�n��ǎt��anbm�����gF���;���{�+d�����ee�9	�1� N�6ȅ��&��	�����#�:���`��N�L��X�//Od�p���3�C�0�:<�<h3��$=�7��x�K�q�{=���u��D�	�~H7�οW(%a�c/�ى�D4��-c=��N����0����cݜ/WI����e����9.��\��`��|g� �1�X��Q���}5^����k�\�'�Q: z�4�!ι �ǽ�y�ۃ83w�RG��P���^<_nt`}݇Q���$�j���'(�1+H��1:zs��G�5�y.[�M����T��� ںe�@q����c@��M�8k��J��l�3��D�i�i4���%���[xM=������\Ap�a|��2��=�lU��?G{�z ��7�Kғplnh}������%�B�l��ETdڵ�3'����q -���^oQ��t ������S�/�X+Qr2���`}Y]��bH�х��D�sC�9��Cڽ.��O�������7�+�â��/hj��b׷��NՃ��.J��m�"�/�||�]D1�ؘ}$a�,S�lOlP�̃�`���;b��m%4(j�у�%�v�	�x�{k�q�1Lu3�&x��m:�?�~8����_�"���OJ�{O�I�,�A��뱔a�k��|J2N�	L`l���sK��,��"�h��?���6�q�I)=n�w��@��2�#f1�s��4����*�?�O����\���m�gԔ�^��|�ds��U~J>���]�6��zrm��}(��Y�s[�-�4��U�^6�4;8lhA8�\޼}�Q{��7�|�	�'���L���GtP�M��/��|�k5}#������HsJ�а#l�o2R�Z�!������t���
��dD�M��N��2#��%O�c���ۓ �1�ۻ;f��#I�XS(ɷ��H�`�lKgc�c�nY��
(�?��� ��`���t?���#E������w�>�Y[��$Ɩ���S����*N�}.j��T��}�q���e�g��pRj =�S�@쒝�eI�'�e�s��2�T<��$v�]= �������z8��[v�C�+�DP��DgTƋ{eU�M����	�Nn���|t���PZcg=m�I8f�Ј$6obn8��}^[[b�o�8#0e��+
�Pg�R'���;(w�)�<^�;4��0��2&��ÔX�	f+���N4�1^�?�&Cʦl#OluLS�=Ԇ��Y$xR����q�)@�_�I|ɒ9���;�� �mܛ s8��/1/(:�}j�M��J%v������]HRw� ��l�����4�!S�hP,C�6鐟�Ri#����C����>ǛT�Q�p����-r��)�l�1�,���Sc���x^J/��yxZ4�JQ�d���d�}=���	���5�NE��~?�3�ɦ�u�99���̢��8V�2���2�1�q�^7m�`19]A�����
G�u���z�~��8/M�#$�rU)6�!M�s��fa��/�6h�$�9أ�h_~q����V���2��۵����Q2�}Z�7�gw�?�<�����MK����V���������hAW��p����X�7��8VsYq'1�`Q*}��12g�V!xpvc��774�؈l�j���R�q����Ŭ��'捌}�an�n�^a�M-�Ge�|]��j�3�M����O8��=yp�����x��������m�d')�Ț/�9u��Y��נ�t�}17�gR�Iɬ�$ek|�~��\�����������cuB�ы�`W|�%�4�b�kGl�jՃ3�����RG��s�Kof��۪M�8�y��.KTA!;@|Ƌ��p_�t�F6in�y��9�Q���!�	4�R�R�,k�#�Q9�ψ�4��f�DU�K�V�}�!�G#�t��D���e�r/���W[!-��}@Y���:�
D����U�a-���|��$����J6ע��xq�!p`�v#�NS_��zK)y`�튰C�Uȭ��B��ӱ�4�PyR&��d\5Y�i��_�O����c�ϙa�ţ�h��|����Ң�)��Y�|�ߔq7f�՚�0nw�fUW(���P$N̹���9�@�AP��as��_�%�hO�!�Z�,@��WLU�D�pn
�v�� �_����(�F�d�L�U��Qw�T�ǧ�[��^��hnXmЫ�Y����H�!@�M���1>�t�~�+�	����a�~����JdcX�Muc/n��������wa���ȝ� z^S��is�d�>��4:�ض��颬p��eI�/d���)��Lǥ�T�Ȧ4a����4�=�χ��V�2�Nc��gK��h�xl�骢sw�ِ3N�{�I��@�D2�V�H�H�@�n7���@������a�̾U�Ͳ����4�[ȋ~�4�麇 h�ܺb�����,�&-��@z�h�^6���=�g�,�ڇ*T�����8���:J.I%uR�Im��Sgm�ߤD��D����ʐ�T�Q\��N���%�k�}e����+�Ď��K�����)���;fn�k=�9&0=��?��(��m;g��� ����q������Ғ��P�A��]�;�=�a >��C0f���e={)~n�j&o_�=ຄaI�����G���O<����i�1�Z��*礃�R2�������Ç.��	�w�]���C�~���6����m�'�ɬF֌ps'��ĉﳩcX�%�+"��!b�l�*��G@_�v&��ϩ�$�o�=�T��3�-��NC��G
3"�Dŵ����#��(6J���9��4���*����
h-[��݁�Ҕ��	?���B���o'KwC2m�pC_�ޚ������Iσb
H��Ǔ����y��ɢ����
����b��������IQ���C���������w�Y�'ŽW� �_�4�'P�م%"��a襠	��.3���D\�;�� [QHJf�� �Lj�s�S����f�Әת&��������b�j=�5D�nޞ������r����}�i9�L��3d)vxږS�F�7�cf�!67����g����d�cOK? !����z���Q�^΀mI�S���n�l4�v)v��{Z�	�	�׼䢏Fƍ<�\~#�bT�o8����Ⱦ��2��x�~0	*�PʯJȀ�����od���f���zS�����ڷ�
��f��L]SH��?��$��'����2b>~�D�ᡏ�������f��p�~���Ͳ>9�X7�6	�o�S�̰fei6)NC�`]W�5PG��/�*�_5��'��w�<�&S��5e��$֎=v���L��Lj���:�����?������A'3�N����@֎��L�S�A�qe��c5ʐ�Z��i|�B|l�jWq�&]�^u�L[�cvGy�*ބE��Ԏ>tr�k�5A�2�cf[�n�"��$lȣ�'u�oB�w�qg"6����äFK�!�GYtW'^`'2/�6fj�A҆����q-��]D� f4}�q"��ָ�g�S�C���� կ�A���p�.�iL|N�L�����u��~I+,H�I�������5�cf\+eb�q�Ry�i��)z�mU�~��������P��ry:I-�Ϻ=n��F�M+w�o2��x��5��]t���]�n�@�?��{���͊���"�c��Ʀ�����^m��^��x�?���;�r�ɖ^�#���e��0~�����4��i�x�R�E���'�_�	�i�y߫��2Cl!���+m�u*�<�N�0���U-�+���9qddHo����`�򺝓A�r�M`5����7��:�}�{b�hMJ��+8���N�k�c�_H'CB��C��u�ĭ��߫�j�T�2jlk���6|���_yt������ĉ�<M����"U�xn惹����[κ��d�k�Ig�y{F�@NoP`�x]K
���et�=��y��ެ����Bd�,WM�	+D\4K�H� y��c�{�M�Ft,|8���y��7��1d|�l:��}ǟ9�cs����	����%�:�����~Ō���~p=0Q�w��}Ѕ�;���s��0����b��xu�F9��DS�04������1W���XL����`�,
��pAd��5�j��>�<�q��h��I8�!D	KP�L��<�]I'��n)v����>֐q^�>��r̪� ����v]O�@I�˗����-��yT������c*����)����Z���zƛ$�c}�A�&����6����Kݍ�$E�"ke���k�'ܻ�ς�A�1���%|�{\�����d5�aW�Ql�L���ȁ{[N��q�0��T /{�؄ډJ��{I�Ac��x߸Hc-�>d�S�b�:t�X���Q�R�h�`Z��+�xZ��;�w� ��s�K|���٩_7���M�K��fbG���$��%Zכ�WH���y�yC?Jb]>��ǩ|fp�N�0��g�N��{И6�J�EΙ0������6��
f�����3�#U4���Ej��%I5�I��I�zC�g����b<͆ґ����i5�����
no�'4nt�I�#��c��n���q���΋��~xJ1���Fc^.�>�@Ut����-�K�n��Ls��?��u�Yl8-KfBf�C���	��)�:���F:0�jCK��/8�[n��*��5�b�Jm��߻�9q�+��d�d�4'
�d�s_�i���?��жu�}�P{�̫������:�R�9�$gu������|�T�u�7��"��)����ڵ����]�8���p]9u�:��x��)�[�Mb����j�9>z}�?���3ړc��Ì��#m�<;���A?�]�5��Q?1nJ7E�L�֬!Y3�;������p��}�TcfC�q�M�k>у��\<l�-�p�b6��S�pn��I	rI��C6~lm�p3��w����۵|{el�w���y�	Z�������&����z� 
b�hA��Zv%��x�'��1��g߮�'�5�������&�G�`]x��z�U@Θ@/CF��&�d�17/N/20a=�y�������5��i8���%��m�=�t�6��І�դ�s�g�'V��۔ٶ���;P�S�۠8m�?<g�?������,L��Sa�/(��0{*�4��9����o٬�5�6ܸ�����[y=�u�/j����e)R�����+�MP�nh �e�t��Z&M�2 <��gwZ#/�9��?�#{�"�g�V�f6Ec?�����>� �h�������s1�t7TW��IHh��
A��E�Ǎ&+��$�;ޜT-l�p��O��̮�d���_��P�I���~q���n/ӅA��$ͷ�.� KzΝ.:A�mI}B3� J��FI��%KMs={����H�`8g����06r���'������K\�~��r��.X�S���z1���{Z�y�3�"*��}�J����*�N�P)�/��pRИ��n�����`ia���������"Rג�ݺ�(�{�� �Ƞ��d�嬿�R�����#������,)�K�fڟ��z=6���'��x�_�H?��D��� ���9sN#(�q7q�)P��R�j���r�t�l#6��
��?�ic�Sv�����F>��A�����<����O9.Ǡ8�Ğ�q/<D�F���1Մ��f�x=��Y��c�_̑H�8�p��L��VY{1S`���0���׿.?���HV>���]�����O���]���(B�P8���t/R���|}Oyp��߱S�5��e�jReݨ@q���5Pq����J����M�F��C�U|�?����͎^Yi*����k~'$X�Y���U��b�sl��=�;nйf�����b���h�Ah�E�	;��p�7�4��M��G~�_�����-:���Mo�1"�σxy�!�)c�����Ft:z��R��	W�K���M���}�LÞ��̓Iu�P����ӲMe��V,!�I㊙���f���l��#�]�NFI�\ܼ*Y�]_n��؉�z8��4W���M�-��im��uQ�px��1[�0;d�شl�<�o��J��]��ON�8�� �vC9rc23l���<ظv��[��a�G��*�`���vbִW��cx\��������&N���s4x;�Hǆ�E�����Ԯ�a��*����N��~O�t���3��UFZ�jkg��RHc��%��`b���T�E�"(����ep��z	*�|X�0�>��ϸK��?��2A�4�!�a�/5�~9�~J�+��1�~���UJj��/g�&�	�F=�(�s���tw'�0+��ԉ���7�f�],rl�ʸ)C��/�����l�s�[��c_3N�K�(Ȁ~��#79�s�+�և�e�b�"����73k����të��7�1�U�˚U��J)���$���ުcn��Gx����ļ��z����v�0�y,�g
M���.𙱴N�qQY{+l�@�G���oF��]�� +d�`��3�Y�f���g�;�˘�e��Aj�����>��ݦa�V� ���ӣ�蝘(sZF����c�)�}���� j�y�5T *�;av�}�]���� �u�&�Yt�cTJ4�O ��(�V���{/F0Y(]�k����4=ŵ(�):�����JY��{~�쇅P۲���˗q���!�Հ.:X*�M��7�|ݾ�&ҫ�^����(ZwJ*�u}�O���փo�O���f,/u6��X$
8�^��:֓μ����y�t]���oS�l
u#U��?���7�ѫud��ε1�E��,0�&R��q+�#�"=ǅ��=;�kw���釬'8}@{������
��7��;n^/&��Hy2KW�Ɩ���J{�����coϔ��po2��WGx<�����υf���R�\O'Y�.:�<R��y
�	��-7Gfpb08�GP�Y�~Fl^7��G�"�i�fT4��U��x�Z��aҼ�sc�SHS�r�(�s:��l���ٱ3�Td
�y��aFRt]B�+�T�6ҩ�B��J��7�,�7bH��n]XO�@�{��5U�9���"v�em؂��B�Q�i,��*��	��2�R��>�h'1z�dvMҁ����S��w�H�����q�pH�v����σ���ˬ3 ����!��n�:�ヽ�7�~~�s��t"`~NU_��T/=E ��]���+��&=�Cŧ��<u��v�71��+"vm��j6�f���K�q�y,�,�I�7g�i�ZJ��+�Ĳ��m\���r���'��G���s����|>�1�l�(/�,7?��#��|[�[�	G$���j��"�ۦ�dqy:�"��yM���{Q����x�w��則�F(aK-u.�؎.��1���� �t����V!R��.�WP�G�����������y�1Y��Ae���PnE0צ̌tK�kRC��j�z�T=���2���7����yv��*��W4�Oq�D�Ce3�fM|dc{�j����ml����^�U&���;��9�|7�T������=���ZA���G����L���2�_�m����w��"�{~UV�
d}/;���tN*?�c��xl�b�x/�9�7���P�8X�ܠ�}���	� ��{����3�-Zf�c��N2�mzf<>����C�AX�C�N>�:�g<��}PU��w�ƞA�����?M���@���]��Ȧ����� �K���'>?D5O5��O�a$���E���?������Q�6�6������8ii�p���ό���$����s�3�JwO`ye:�P�e�V����c����RHPZN� X���4Q�������uRf?�N4m����$���2ȃ�O'O�4�b��%�g�
H��{2G�(3�E4�QM8&�v�,{�����"�&�E���ڲ�V�k0>܍�.�.7&���mO�c��Y�R(�KA{�mG��3�Ci>G5Y�%a�j�5c),j`�]���}�>�7�,0��>���~=��o�`��
?p��cl��b�l�����,�v�H{s���t%���ٜ.�����%:�/��B���/8�h��8�wn���Mv�r��'%1� ���4�&i�b�H�#�z<����dD7s,0���Su'C�9\�񲗪���>���� '�"��>*�8�!hI�A�%�����(tJD�Z����U�����^��g��s���(kW���ݺ�;�������3K��fw�I�es��1B7�=�aSrv<��A�;+��A6�)�CU�+������7k�p�yo�@�:9�ce�C8�[���~~~�:NU����G#*Ǧ�r8��>�⼪<�l�S6�↊N2,��2 ��f�1�r��<��$�9�S4�P�,���E�L����su�CTJ������a��NX�g�{4�iJu�i��9�M����H� ��]t����$Í���>�r��Vr�B\�+��f^hփ�^�=�GmBNv�AJ&(��������yv�	A��b��ce����B(����.�i��\x�������Х�PGL-%+�(qO�hm:c,��"�R+�iʪ���h0��
�dѧ�����;H���kr��S┡份�k�.b�R�H�s��!��.0Y�e¾o�:{M[>�G46�̢�=�=˦�؃}s?�=�����1�����FS����z��b��%���
P^�(���*�n�) 9�g���
]=(���{I֞��¦f��9G0��8�e�L8�Kn�kY���t�;�(����O�$��ϯ����"K�1Mģ8��x���e����3|�קQ�aK�K	]קYt���i-5�Y\ü��/mo�%ɑ$��G]@����!�-g������a�4n�*���X5��z�o7��BWeFx���������s�[��*P���^clO���
#��3�e.���$�[��1�U��<7��wZF$�i�����s��B͉�x�(�E�R%��2x>�ª��������$��k�R��:xѯSPO���EĜ�dY�V`E�C)+j��WI�y�':텣��M]rf�b����!o�$��_��2j��b�x�k�](]�NC�=�^԰�f�=+�(��@	�� ������ |��±lbj�s?�h6
�q���6�	-=	�e�N;��H\<��sS5��$6T5a�Ƞ��Nec���`�H�mܵi�H�C��N�� �l��Bo%`$Y�������������`��5���ϱ|zlbZfpCQ�i!u�EF m�o7
A뫯�7�~�6,�(���4M,�/cQԾ�xl�'u߽;F�og��n�Rd�AM��ei�k'ꮌ��;+P�<�
Q�|3�Q�y��i�T�~,�K#^y,��w�5i�^+A6+6 ���0���D�T@�e�{��Y���Z�����4Q'�}8�5mf�b���$w��
W�LEL@���}��V�ؘ"�����q�(SO�ȘIQ��@�n�x�Q�#����m�q=�F��
�v�4=oə/GT��6�����/,��r$	>�(ψ=��_?���h�� �A� ��W_�����,����C�V��@gB��1�ĳF��0�:�d��z!����P��o�f#��Y���R0��l�`������ɵ�&�m�E@9�� {	<ԃb��<Hf���u��Ҥ�	6L�K�{&A����Hܹ�R'.�qդ���))���m6�i�^~n�L�Σ��r`P�I�]d�V:�)����h��%}ǩ�`y�xn�gk���̱��#p~�����߾����6�$<���"����t�
*lh;�i�2�m�b��z��K?��w9�����r��_�Fy�����+��߾��0�B(?�r��0�qʖ�C��{��ٮ����g�)����q��I�'A&��B�:�]]�D��ҽ�����>(��D����G���5w��Ð��N���b�"	'�*����O���YoNl���G���>)P9C���ޔ��u&���]X7�	��*�t9�4X�n��/&�~����/|<�R�����"��k.f4m��N?Cs�ۀ`p�[js��\���ƴS�٬��$մ��RT�Q�P��q�!㎲~|�2��l�@��f�H�=d��Hn*�Pۚj�%���^�ЀQ�T���C@{9��!�0�<[/�Q�WQ�!��_�`�F ��]���e�
֘��f�=C��;][z9(��Ǎ���bŉ&�gw��Ͻzyn��*N@����:����x{vqF�a�Xl��V�=O�<Z�>.ґ{��(f&��W�H��6�~�>�#H�?|���[����_b�=`:���c�f̀z�E����z�˱j��g�yMk9?l����&�I&8`:c�w��F�(��X����l��bs�;�#�����l�m*K��w{mJ,�q=�y\Jg�,�p���}�Ld�fJ�Y{V=����4N'2j��� ������Έ�yhF�y���X�̀ץғ�J�<�e
�iL�m�<@��x����3��5�}���yx��8i�W���X��kς�N���Y��áʺY�������^���7����^�{�V��ƻ��$t��xS����Z��RQ�w{K�P��r�Jχ��bܧ�ѱ�����!Uy�6��#�1����E�n��,qlT<䛕��I1��L����r,��<1l�뛄���|��z�ƛ�����.&Nc�P.[�DF:*#����]����ﾓ�{R7{�	��,��!Q �'w>#/�����9�}H���?k��c#��F���������n��׿2C92����E�.2J�u�BN�4 �u��ʦ-�A��tp{w[��Ue�v��C��R�O�U'	!FlXa����^3�K�V? �B�F���E5 �[�aVm��'|��[�Mg�9�K[|�_|�(�dҺ�Oy�.��q`L:��+0�a��<�k���ӟ�k�ￋg^���8���l|���E4T��|��j�@��eUPj�:��z/l�n��9���v�x��X���%��5|��;+������������%��A�XO�7T��Wg�\6��d��5��{|�*CG��
� |����u�q`�3 ��Ž����z:�`���@l���z0�i��V�4�d���.�h&l�©[orl�3f��t[8�7�x�W�l u��
��h�T k�i~rH��I���y��DX���N$:FL��e|y��?1K�)�����v��^�pЄ���t�I=F�yL�
۞E���f�s�p��v?a �����������E�U�9%�~�l�����m�X�R<i;a�{U#��x�; 1X��[Da,�U'��b��*�rF=�a�}{i��B��D����*�^�e�Q�8n\�Q,�;�Ԝ�Ⱥ�sނ;�∺����#(a�%
��:�˼$_��Ui�F��wӚδ�e,�b�Y�o)���/�U0X������4q$��a�I˕I�fB�S�
ĵ��S�ߖ��t��"�]�;
�=�^�Qdh]<,+���Lx{��fa�b��2)tӐp@���_��yVmAPu=��.�,�t�~���=�����,��i�T�[�O��'BR���T�r�|��k��8	�� ٭ȸ�I��'k�,�"���:7���Y���,��'���t�R2FC?����Ć��hb�5�q����C���Q�MN(��^̄q2�b:�J�^��=�u+����:�8Q���qt�c���di+V�x!�I��}d�8���pJ3�l�4M)��������Zό�)~���Ked-���&��s��R�%��T^.P�W\�����"�R5��e���-����t�"Zp[��L�i�=��[Sy6����ZF��u����DB���0��|��C���Zl�&���L��?�#[�鬑%/^+�7�3�~���pJ��0�wI��GzD6�$ӍIc� L�̽��62�4曦@mK�FJ#�������of5F��W���޾�Hy�� �7Ym��{�,�{vH���j?�!�.8���/�|�ow#�\#�_)��.�Yb2��$}��l#*�`BL�J=��لrR�I���!�K[�2�|)�hv�������UȏC��U,1W{�6���������D�$~�(gwi�J�u=vzG���κ��a|�@����GT������b��Cq2Yrƍ� ���$G~�d\4vv����q-������|�X���nh:@����+H�Cl�3l��<�rn˼*|r���������M�و�
YFf��!�M2��S�\��&ס�L�eO�rpw��b�lE��TtO�˒� *p�����~�g��w�E�A�^6z갻�剘)!����ݝޫn��}|<�fюI'4gm;��NVb�6���xֽ�`T���f�^2�j]ྛ~�^A��z�R[���*��@IH
A�>�R��f䴈PSi�Zha2��H$��1&[�5`!�<�i<�b;��Nr��W����k�e�X9��H���y��T�������Źew�Q�i�3c�$Hͦ�@i*\S���43M���f�WA�E�y�|����aT��e/G���ₙcY[���$'F4JE�r�E�� ��䚑��Q
�D�.���ӘW4*����|�M��G�W9K��*�ӹQ��Ԍ�i��,�9�Å
��X?��ctd�	�������j�6��Dq�<�.&�6m�Aq	���N]m��ً�S�@S�[�\��o���[�̬�X�!����ُ�\���
^$P�X���I30���$΋�@|^��_� �y8�q����gqρ��+��r2�qm�t#J̾�No�jH^&~��v�lǇuT[�Wu�kgE������6���1�����nHo��)۬�t:Qm��OT���!f+x���b*�Mœ9�Q�3�[5����Tw�7�/���Z��JJcG��b�9�qh�k�PPT�:����28yև�^�m�I�33P���r�٧��R2R��9E�3�L���Nh�.+�v.�K'�m�T�}�f�L(6g;V���}r_�Jg|��;��J�(�҅��M�/���:'`r�;��o,f�fp4/4R@�D�e�#�
���ݖ�qq�w��1�$��R�i�H�Ji@�Gf?�����l�sI�R�=gY�FE����d���X;.��Ǣ��b˰����2�1ć�C�lCeYO�1?�k��m�ב�"�ޠ���w�\c���ƥo�mf�8p�3c��D�+��d�ēRMr��Y"P"S�ӟ���˿�Kd��m���.O�.D�&�=N�%�#>�ς�NX�af]��⾓4?&�j�[��@����C4v.9n��f� �0M��z��{�m�aJ͊�~�f�FجĨ���tO��Q�k��4O�(�����){�F��<��;g��sv��	�'fJq@��P�JF_� ��oD��NA��KN��!ݲpݞ�6���uY	Ն�N�������2�.�ͯ����Z�M݀.�k߻�gb��NknJ��`[����Mۖ~�_��e)?�t�T�ҡ1�����ڽ����kx	�*}ee�l�󘭢�*nD�GH;��޿��D9�nJ�%i�^����I���3��,��@����+��3o?OW�}j��O9,KC��S�L��96�KJ���Jn�Y���xA/|D!����FfQ7��h���SH?F��I��H�(1�j+�q/̑�E�vaI�qNp���m���Ds�h��pH��I����n��_�5,�br���=:�RY�f��C&�r��.������ ��H���%j	w��aAVɜFɸoab�N�o��L�7{q_� *�B��24�jC�Mr}�lA�Rs.�/_c�ف��[4�1��CL�4͹v�j�yW=��gc%�V-S��ZP�8@LHf@��{�u̺��;���I���%�nfB���y����Gp��+xw�3d��{���%��+^sf&�R��oT?�ҥ/��Wa�q>-���0Y�,�##uB]�ir��]��3*�����4���ë>�8� �|M�2��� q�4m 9��_*<ћ���m���UI�j�s�s�+#5-L���8�d�MbHX��[���"�1��/��es�5N��<+96� M2wpF��-4։^�N�+f:]��a-�4�6z��z�@Kd�������������K����W�J
N��=7є�M�y=�T�՜��>���d�m�7�(W`}�������xV ���P�<����w�4M�tHCeu[y0p��R�H���0&DA����k9@���9�N�e�@CF����J\Qz%o�LW�w���ްm��Ѡk?����e�z7�2) F�&�C�� �5�']T��V���&���IH҅vW������T Պ�倸�����%�k���!_�J���_|)��C<7T !�>rM��%�^�c42��|M4��8� ��<�#�1ӗ�@�r����x*���� tVYǸ^�3͈��"���Wd����3!�JJפ���������*���(H�r�����e����n#kG��7� �W+N΢��I=[}�����M4t�Mn,���v��w�������S/p�PoL��.��3x���:�F�V`Ҳ�42�$b�g�pa-�%7�f1T$xQ�ص���7L���� �cVxש��9I�M��ߏ��[@=ׁTʝ�$�/�d�xϿ��/������őƏٔ�Fu 3���@���SaXn�ҀƎU�E�/��s̉��Uކ�2,ݶ����g��#G��ݣ$�V9�:���ζ7��}�2oպn����A�e\Ot�qH��"x݋PV�͊=�z�gB���%2�+Ǧ�tWդu���̎#�G�i�(>�h;1q��Y~�e<�A����|X�C��D6I����_��w]�Xz�걼_ġ�Mz�l�y_LMv�eyv���x*3��b�cmWUn�&��q��V����v�U�;�kd��>� ��T��Q�������Sڹ�h���LS`�;��J��)����.�Η꿥��א*l����ԫ��>N#Л����=��z����gƍ�f�n���S��7?m%�c�z�$�ԝ�&��(E	dc="�~|`�?��u&��� |�]�_c����TL�X8X�p��R8!m��ak���Y��P��X`PK=�i?�Q������`D5��;�\�H����(^��#o������l�n��/i����+g \���iRb�L8�'^��ɍ1\K41�m�h�^ [��*��48^���C��9�E�� d/ �= ����(l;3�rmωi2�Sz1<>=�&$���\Q)�hޑ�iB:�?�<KV3>���uJLv�n��(�a�̭�����D<&֋�x9��&�R6eO��BvyxN(G	{0�8���(�O+�h.q�5_���d�ltbo��E�t�\f�i�zn&YYׁC�s҆y���FO�v����wU�0%���s�rh�ݤ�v�'�6+�o�wLI��)�eR�E����B�mRƚ.�&h�[.�ϱp�f��l�P(h2�g��y�DBw�t����ܝ���t��άH����Ԛ��`�a�����)Xp���4�">�C?)�]W0�QC�p���%�&)����q̬�e�4�-+2�t�r^i�pT��fe���Yphs�h=��v��$wR��o�J=�)���햍"F`s�<�n���'kʣ��d����
�U3����A�F�A+�B�0�F��lm'Cq@�s����ʃ�MfǨ ß�͙�sֆ_ �}�"�ДLO���r�����1ߩ��h��j�2ˣU7m�b����n�[������P��4�V=a���̊3;��2������i�pJ.��S�
m��'ǐ,�)ް��Y~���;枳�O���V�v����m(c��!Kg�fk�Yp@�EK����*���7����wS�S���П��1C@�8����`���1@[:T%�Y�ˆs.��	3#��8����97�OxS�U�3�wJ�J/�2��KN����.5G��('F���z�'m&�g������\�<7���68�Ҋ���>2��T:�'u;#�u�F)�y���0�X����"�D*�kh�=Y�%$0��&A�뮨GyL��Sc��r�(Z�$��@��}f`��̴� �4pZ5n.9\�^�? `�ؠ��"f�>>�������2q��������X-�5�1����~U�7~��%�k���jp[6�i`rQC�n���slXVFR��EIKD��Y�3��N��qO�%;�k���|WF�D6׀5PH�0�6���/6H>s?{F�K}�{�v��Z�e~���w.�B�w�RPPs4ɜ U���M��koa)͹Y�|��59��Y??�ǌ�;d�]6�@S��,J�J�>U�������r�m�`�KF�R�&�K�3g'![cP����S�����?c���tb7�K��S.��Q�Y�62���4��c�1~�H�X�m[H�{M��E؉�_c�X�6�����<�5n#�nU��̥�G��8]^zzfdx�0E^9���3	�����玁'�I�*�!切���;O�8P
aL�9�����s�2̂��X�-�Q������D���� �88�02x�ψL�R�M���:Kj���`��[L4�����Q��q�q�Y.�|��:$��|uô|{#� ��Ө	+L����ಪbj�Ͼ�l)�:]8(�����4	quHx��Q	M���A沖��]Q3����\�A��?��;%8����\��:Q*%?��%��@���E�t��K6��k���DcpV���[�r�+�V�d��{kM����Ep����p��G�ԕG�j�)�֯� [J���7yA�a1�~�@�`j3| ��	T+�����N�,+yZ���2��Ix��z<����6q|�����ȑ�ƹ��pG.S{=�B�m����`锞�)�<z͓?As]D���he����"��w)_{N��� �I�[�1�qd�n9}��� �gc�jE!qY���(c��N� ��-4|Oݣd��7#�n��g@�q�Q�4�=��d��>X����|`^�.�q끁r��f�\�͉�svs�U6G.t�w���W�o9r^���"[%�=CWi���w�=�0�FM��#���^��$��K� /�B���m*��������6��4�1_zH!��.�_~�eN���8d�us���,���,JIn_�Q��T���#����g��G�_������;b��cjH[V<
��.wͫ��f����\���E�&fZ=+x��6��+OˋL���Ձ4Ae�*���ɂ�ê8�q�:��-����N���^8��Ŗ+2m��)��ۣ!����Ҹ.�EZh��Q+>�5�5u�]}g,(&�T���1�?��!�� ��8T�l��u�m����*l����Y?�M�،����K�8*��נ<0��X��ٚ�m,�'��Xg����%��{w�?~|l�_�}X]��añ������a� 4�(���q�����ǟ�xp��Sf��.Ql����d?ٰ���_g�沺J�N��>U��n�%~�'9[a�̼��SJ�s���no���(q�-����F����.l�ĝ�/����s�)3�h���З�����J�$���9G�3fb�����Ҍag	G,��]w�t��bmc���0L��X�bu�iT�lx��4�ȴ�ݴ�����I������W_4�)����)��~��.pX��x{m�}6$�R���	�iҫ��t㰩����7&�<�F�}x W���
��]���v�|�)�c�+3G �%��7��г�C:����@�,iȌ�;�/��t׍eH9,�jsT�ms�Р��K�,���[�}���
&o�N]�y;)���o�=��+��t�i�̨m��[ß�a�z����{�V�lxJ,i4���g&�Ɗ3�e��V}Fv�R�6}Rsa!�/�7*ooڰ��Ȫ�`np/�$�cr��|���>e��M�e�� �*����܀<�\c���3����a��������Į,�F� �؟bM�x����י`���q��
@��Ph:����և��u	��z��q_�6y��&*5�rT�%����ͻ�-c~���wKc��ujI��ޟ��;�K�{�-�%4���`�/�M�b _�p����՞t%ܑ}Y��=)�w�ްq�>�u��EXm���l�:�������,e�(2P�z^$;�O�p��(�t�4��q#�����N���p��&�����>FT�4��|Q���j��P�M�sc�����1�1�"�M�moZ{�DK�}_�ї*�7�>T��+�eSloQ׵����B�97��z�a�@=�{���mT�س�NZ�����ѯW�s( &0CU����&��-���8n��0�o�,\�䱰ەl�[��`�S��R9�Ҽ���|�j�͍��f�sSSB��vr%��nJ����5{���~W�{ˮ36�4Wt���i�lx��A���������g������Zw�(s��T�:Q���1�ʠD�����i'8����l1i_�/��,���j&�!��|#9��5�ak���*Yn[�)Z��֓�x� �	�M4��'A{s��C$��_�^��=�S�%��Զ�RhC�������ld	n�(;D �2R���r�6���	�f���DB#�����`؊	q������4.8Ci��ҐX�uĀq��wl�7����RT�_����GfT�������P�)��kz٠���C�s�y�|��R�_��;=R�{%��6�uƀ�/������+��`�1K�����Gm��{�L<s��:�{�DV1�3Ͱm��f�"�dT,���22Wx��kUҽ|#k�@�á�%B��A9gn�
[,
-X�1�'#� >���u_�70Py��D~�R��8>�,�X��.���0�d��m���-�$�>aR.�C�Te�ӳ:��8]� �:�%��<�>�}7�J��͈0�ޔ&sm}�D}S,$q�M�2��C�A��}��2���|PvU�j���&3P|1#�l��(���ܼ����<�������]J�J�Ru���L7�C����b�:Z��~
 ͓�ޏp}�����Fu|an���x������@�.�up����1�~ l�:6ö�!��0�0~c�"GZ�Tj�U&5�pJ��涌��i�B]�D6:�`��N���q��_2�H[��?{���-�󂾗��L�삞����O��cÍO�\�Ӑ�52Ͽ�}`y��ϐ��<?W�0���(��}YqOCࠒ7�ޗ8p@c�2P�p�����ͻ���D�S!|����p��qzo�d�nS5<'O��z��D �O�/�M確��&�~��b!vWv������5�1R��{̸��{=(3��(8��?Sz,a����+������>j�wK2yΠ>$��1*��:�����Z��'{�:ؔy\�+��;�����jLm5�[e{-�d�.��u2D�}tW���ܧb����Y}���r��y�&�4M9��%���[��
�j0�������b�n���ԙ�L�0rs	/b�,��б(��`� ۴ 8Acc���p^��ƫp.J��W��
͊�R�M�a��AϽ�A��G�뉛��B�F���,_���u�����L56�v-�N���-�4�<4���{��,�sS��:��)��0��e)2��� ˒2TK��9p�M�q�҅G��>>�K� $���P<��y��2ݗE���E��!���D7ő_���2��܈'q\a�;�^��93�������Vٜ�d��
���>��XT|�������[�-˳�A1�(���r�6¬#���TLpxcnf��Ţ1"8,�o���b%ם<)&��;)�)o���=�zu"��d�{9��Zk8�U]�GK�F6�j��(��WY&�R�Ӆ�Y,˹�8�u�s��徃�C��޴R������ٓ��(�d�kS�&:��lBf���_5e�������'���2�Ln��F*L9k�	X�(#�,��ǌ�v���ƬZ��,~�4�8������F���$wbww��>Ǉ\J�	���=0By��)�m7���#��걳P̓�u� �W ���5���a1�����*��Ә؛ڭ��M]2�L��Ӷ ���:��^�.�<� �N/7>7��l̋ڦ�A��4Gw��@�86uOef5yѮ��0�f���C2,�C��+0���߯g'Y���n��"Sb��#����d����5���ϨƦqMlh^30<�A�>p���X�1��FlPC`�"*3;5z�>mL\��)=u}�v�i��㙙�@��!�_#o^�r�4"�/�41�纕�{��` ��BL�f�7�^���U�YU�]��A}�ϰID���䁽�SB�u�9�nNA�iz�R��:����L��06=	�ROO;�@�	��%}�?���A<c�91�zo��e4E����5%SmMm����H�ԚGF��8�"+@ E���	�p����O,��������_8��&=�}}��ߒ-}�x������6�^���0Ͻ��fm�7�-��F���$�_M�5�]nv�ƽ�=Q�ƍn��i�\`[�7�h��1�d����?���m,k2�*w�Ѭؑ/Y4J/N�8;����8���_ŵ9#9�M\��ک���;ós���!g�tS�f]S��r� �����ր���Cʺ,� :�\�dM\ {��'��(������?���x�~�1~�� �V̆ɚOWј���>W���H,81���3c2�׸�ڷ7t#��6G�)4%52�b]���R�nu��X��3�1�X�?�+�6f��,y�3z���=����F��
�E������N{1,N�bA�@G�g<�Y���GAp���^��p��z���Ax�JE�����U�������|�!�v�c�y��8�XK�0=E������´ƕ]gUΧ9t���+��P���yvٙ6�T����u���%VL�~&N�(���H�ǆ�/N*yZѽ��C;��RWd���r���NI���1��E/������'g��ˉd��X9����4	����4-[�a����z'�Y���:��e�ъ�]5�JJ�]~L�k� �!�]���m�Nnȵ��M�t�r�i�~#`i���A��bq8e/|>�)i�U�&ԃ}L�->_�͵�T��J�'|Q�J�a��,(X��MX�}�k�4��ڰ�^�Td�;gI��n����T/�M�y,r�e�Y|j��Wj���-$����#Fȇ���_��p�x1���g���{b����~�d��P�lb�i���Yn��]i�n�H��ɺ�7L��$��.N@5Um���&qfS�z�~~Nt||VkR���0
��p <)k�,�"-�T�;6��M���T�1��)��aQ��#�ǌh��):5m&����ߨ����5(�����/�Y�ϛ����s�����A�����Cxo���w���8E��Ą�S�r�Y�]fk[�>ϓ�� L��`nY�*�S�������Ʀ'�Xa�pfԛxp��a�	T���*ɁcE:aeG)����>F.��~�/e+J�[e�&�r��Kq~wr���8f�Nd��������D)��uQ��ܬ9u��v���Pe�3��4�Ep�qo��FCI�`jf+&S���;V�q�T��>/mn3
^���������ʺ�kr�~u��ָ���5�VKf'�UN���,���BZ��X��oOm�)x��!��ao�S�Ϊ�F˖D�[��L<�����2J��4�;�s���98�7����X��TT��FD����U|0��ج	��|����$+�S�eC7�i3����I�7{1kl���xP��I�T$�sJ��9m�񰽖�ּ�O�گ��x��4u�Q����rڞ����Y0X'�pX�ᦛ������b��@�}�}`���؂&"tG�S�f��lY��pI4�.�Kb7�xQ0��J�oH��@̊
R�l�\�'�"�p* �OLM��k�gPF>>>G ��6���t�o޼M�2�~~������M+�nw��]���{��K?<�:�#"�h�[2���;�Yc	�>}-��'� ���_4� ��{`�LIg�^[�%`݅	�=9���98āՐbi,)�Q67�3e�y
����"�{�����R<2� j�b6P�T�é;%f��n�d��F�d�T�\�}�ad�^�i�����.����UY���&�|AәŪ�L�1�t��o������Q>M��r���I٨������PJG����!i�3Gw��!�S���kAL�i%*q5P'gnBN�ԊK��Wq`������3���m�at)��|]��� J�X��nڼ����.UinP/�y(qJ���nt[Gp�i���h��,{>�a��}�9�T�0�d0�9~ߘ�%t�B&�ō����`�E��)�~Y8�� x.~3���5y�y�9�|x6fYȓ�c�%o��ˢ<����?��|�Aux�g'���)J�Yۆy&y4�@0�TJ�����{�9@�,��Feea�f$�R��ᛵd��V	�1C2!,C佚��{�n*��mw��ù��g	�$�������([�!�X��9�-��kڙ�i��51��oZ̝e���g����gLh�8��E��c�,�ָ��4B�y��tU:e6��tj��A05�c^4�`
Y蹂]w��P��%��x�$z�%��巌��y���DP�l��Pr�0�=�J_F�d@Ul5Q\Vb����,6���1^sQ��:�����A���eucp5l���iu̓���H�oZ���<�H�ba1v� >?��F�w�)���%� ��C��h�ݦ���>���]�H��)_����=b�&Jh^�I1j�a
��'�N�o��~j<�&��ܯN��4��h�=~�p�8�<��?�1L=�Y�a#8�,�;���y���]wײ���I%�����^��D�iZ+���H��I�.�M*\�(�=ӕ��3��Z{*���.����ŴLX>�
�,	�2���	��EdPZr�k0��� ��:n�MZ�������au������1�n�{%��w��<��{i��d.�3��`J�V�gѦ*'�_U/m�\�yT������R˹��]��πR
 nץdf��W�L�W��3���)��7�:j�GT[��B\۪_p��ppHu耯ej�ِ���⩮\P��7k�1��� w@s�H쬷mϴ��4��]36� 2�@>CH��Q�y ]��"6��;��m������:!��Q8]�KEO�Dn�M�d�Gv�Tq2���a��"c܂��0#q �pG?���6*ֳ,�z�:X������������K�����N� �i5tش& ���d���aP0�,�&%��\�Ў�/6>(�����j��┼�F��7�X����G��O?�������ⱽ}�/�z\�>(�ѥ�����A��%�~�̂"�+����G(?j|G,�˰��#�/� �>+d_fk�P��������)j2��r0y���<>>�̚���U��i%�~O���C��!'�YY�	���s~�o�Pז15I�V�_gY��d>�$a�9�]�'�,,�u���S;���A֒.�|EYT���D��9J�k��Or��V8A\���E�/�st�=�k�;��=g��f�i�-wrXZ�����3x��eBc��c&H|���A��@�З�wa����Nji2���^
�1�CH��"=���h"�s�̋�>��
�w �h�������xsQ��}�>)�@���cD�qB����~<�g�
Q�	K���x~���ũ����nB`�D �F��ہ�!��"���y�5-=��׎����������Ο~"��2ԛ�U�+g�}���q�=�o#�n��<�n��|�IG���ȝ�-�e��o�&��}��7�Ձ� ��$[6\�R���2�&�fTW5r�?g��y����sVW}�3R�0�T�y�l�cd��0�e,Ψ��5��M.OJ�N&0I��̣R��B��G�\d�,�=+9N�k�P��N\�6�[1Ľ��� ��o����$Nko��*�2~�TA.�w�t�Wȴ�Xq���&�v�z&N�C�I{���)�ؤ��wf׬�� ��:�RY���N�꽫��T�2��⻚/��U_M>�%�+Dg���Vu���49#� �:#-1��LF�@ڔ����
ݎ��БG�T�ߍ-����VG���B/�ޙCKG�_?b+U|1�n��F���W�X��$!I���J�b������u������x��aC�}�۝�1L�0`�$��pP8fX�vYo%+��D]��,�?�d���J�5^������Q�"��Bڭ���H佨b��'m�/�S��3�< ���/��N�/ۆ����,Ɠ֤��|�1)[x&����5%'���������+g��(K�u"��F�q��5���|Nbd � g�Ee$��;��im����̦*���D+;��E$���l#��y���I/2���D���hn.A��9��ZΑ��]��9�YI��x?ާ�m�*�y����m���'fK	fיJ��=:��r#C��!7D��}G�*3�i��w܃�T�1��s�#ڶ�/��U�����zN�I
�?ǽW�|.���u)�u�n�^� j�>I�0<� �Ĭ��K2< ���I/�u���/��.�#8�)vk|��N�qN��eе
��4s�J���/�
�r�����H}ّ������7���E/����駟�x��<8i�Mß�=��P2���E=�6H����Wo�����n�P�=G����S�O`%�� Es ׎נ��)� #펍������*c4/����F��b�� �Os���ŉ� �v>gC��Y���x&���L��M8��$�A3��Z�� ��H�?oA����;���D������1 ��}0��'���--�>;!�3�E	��t�#P�@	Li_���H��SR����Ħ%�ƦN��=��`�۪��{Ѻ��m��~'���)��,$��1���[y<p�Oߍ�����l�B	��T��n�u���!
�ag����\S��o'd�ϱq���<���^A�G�W�}�5��0g�4<\?�md;�2�^��|�����J����yev<?_q[���^� 21�t휥��o���d)�2��A#�q�$��
�����p �7VQ��&�7H�	�X�%����M���HX�H�h�C�w�2 /
��������Y`Q�K�["�k�{��ft®��JWS�����a����.r1����.6���p�D>���[��D�;��@�׻��n�~7��d��Ɗ>n7�*�, ���ؠ��NGI]P����;L��.]���x���N�q�+�)DzR��\t��^�>,NF�5�0g����(���p�0E��Rk@���I�m���ta��ȥ��ÓuC�����`����[0�@�uT��^dYr���j��ˢ�޷�J�Ms�c��M#Ck��ڀ{�!�?ws8p� �� ߿���7���6���/?��������ݑ�Fl���(���f+���-dk�M!HrNzN��<�x�@p��/�}�|����~O�7]$F6/dN�z���a��@;Ӿc ŚG��s�o���=F���Ҭ���7p�9�9p�4����f�f億��|���~;>ӽ��Q{���{�͟��&l�f+�O�۵D����眢d�1�`]5�'�%�L�FK���}��7��8���@�q��6�b�L��y|d�q�(��5'K��=W�Mq�*b�Re�:�<�	�onL�_���g�l3�L��t�)m��F��̛>"x��lyҖ��iX0,�E�^�X(� ݨ��iO�����?b��|q$�I3~|�t�6jb�KwR��s}8Vc
��)p9�{�.�X-��ԚF�;o�Ԏ3r�����(�E���P�0V�z��yFZO�$��IC(��%��L�cPf�)ʦs �`�й�/�TwUZ�ع��XfyM����u�{�1Ӫ��\0he�(�o�SG��x�z'Ïm0���嶆c愆�l�ز��b���hH���.q�e�rNyl&5c��j�e\G|�ܦ�:2�(�#���!+6���g�X���S�+e,�=+2n���=B�*+�	��!dm|���(Y��fI���LƳ0�N�F�d?멘|֢1g�x�8�&�L����XmIƮ�kM�+�֪,.x�K�h��s���X+}���]?F�����JW��_�is������--�'���%|%�t����_w����B�n�7�yYx�'��^�R݊Bc�.w=;�zk�,O| �Z�T�1�AJ��KĦ�M��4�?+zp��09�6��%\c�vuIղ�x�v�t(DMµ��o�׊����)ʖV��9� ��o�gv��k�tcbv�9��Hd��,���[��������oqx��͙3���@�y:����:� �N2�54����y��V��M�o۹,F�1�]ݥ�S8��,���أgڶ�� ��aHޯ?���־��}�yL:����`>{I`=�q��ro����q/A�3aj�b?*����M"|��_"X�M�G���NH�5���<�zә
���<�Ij@�g�C��#���_a�"���I�׀o���u�ָKޯ�=�>���U��iK>үb΁A�c��,M��5�rI��{;1�@)�1��yl����ۃ$�Or��l��ķ�`�k�Y�wG�%Mmm
VZ��?�G�2��"�^�Ц�Qzh�@��$;b��ֵ��u�� r�b�f�x��ڮK�Q8׬�t�1��q��.�!D��L7%�p�j.[�W��v�q�|6.nD�D��.�%mſ�C��RG��<[׹c�I�\��ÿX:�ylL�/��+�*���&3�V��օ�]����a��Y3�,R���F��N��ۆ#sM�>����U�/AɄ,�ǭĆ��?� �-�Y���f�`��r�՝hHX#�7�=m�I_鰲
-�O�({��b4��3�l�b��(3/���9>�YA�����M�H�'�=�)*#���3z.�E�P�=�2�ԝ����d���:��Z��1�Q��rfFM�7��0a�I�(�T���=�ۚ�I2����k`6B64͞%�5���;�a95�����I���/<�b�{J{���B2�]'��c�b�Pp�'�)�C��(�	fC�f���T/i�����;�g7��^��j��ŋ������T-�I­2��-K�J��XO��,m��=�nyN��>ưm�\��:&�x�,�Zc�������j5]öa�|����/i���?G@���m����5y*K�VB�� ���P�s�J3���A&�k�K�FiEcj�Ņ�(��В9�^�l/��I��69�wH����"�����G6�os�a�>h;e�ͮI�cL˒��x�d��T.�T����{dg�q#[�����?��i��
�"�rh�GC���nnL=���D+�pHI����Nb�ΰ���~Tkm����l�N��xm�*2�ݠ9a]2Gf�0��º�tд�,��/g�O��@�,
g^5��q?q���1>ײ��ʡɔ\h[�uZ?��������hY.�g89� �jÉ��ɋp�sB��uK'6�;ChC�j6�j��2�!���*�z�Y�Ћ_�*#�"�q�4�~'#m���5��?R�Q���n���q�	�M��2(���y� v�悫\�U�)�p�_������^ȸ&s��k[��{)��"a�"�b���!�>��
�qʽ�3O�#O�M��  Q���v�,��@`�:�0y���,�f�9��-���Jn��3E��	���N:`Κk�9=�����ޤr�c|˜�Ix�����Y�̳�"CG�f����	�*��t�7
�t4Q���*?C��� cMT����6�u��A�ʵ���Z��:8�,�!� �� ����/#��J�׀_���	��v�M��k��NW)�y���Q2SNкS�25�-�](�.E)'����T���J�S$��w���pf9'UR��|`�9��N	��қ�Ik�<��'�9��Mr9+ZT��mIJ�߸'�$���s}���A���:}I���@eZWl�LM8j܄U4xk�|�+��$��h�|�{�;ߺ��5m�E�R���w;��A:��u�)�F>7��7Sb>�؁�q/G~݉���1�<�\o�"�ax�S�6�0�ȲbH�a�s��Ϣ�Pl��I��$�"��T�-6M���}p������,�����
���͑��p���>%l:f�_���tN�f��&y^�*��3=-��F�-b���2\n��@RM���OM#�)�|ʶe&��K�θ,5V�HRI��׹a" ^��&mS�x�0�"�~_e���C�t�?Ŵ����j���f�&u������8c�fj����wsS��<��4��7�gl�s��m�� :��9h�om2�Izo�c�1JЅ��A�mmoWfs����5(�YG��X����-K����KBqe����l�Uc����`Z��1���VAx}���z�����?�6�T��%�$W��j�Ӓ�f����(G3�X$�/��9�iu�_ ���P�͑PCIg��B�D��$�o�0Ң�iub�
Oϻ|�,J u��@�a�(#XV�j����s�lx<������.`¶�r�K�_`��2]s�c^37�>�3V�"礟�"�l�fε��ޱ���|�,�c<[��R6��s���]y��E@��_��u��+�#4��bY|�ή���$|tl�ؔ}�U"��o`|�!🃓����n@�y����=w6�H��#]͓9٘f����"���_�mp9)�El7D����*��,�U��(�×a\3y�X����<)#�Y�B<�p�K��^8{dG��,'�d��]4m�B���V�6��4;�[mSd�1��5�"��t�)ẫYMn
{�#x\�y}����J@3���b�����������_�o���Rx� �۴c[���=�&1�>��f�N����"˙��QQt�Nr��g)vm*�Z��w�&~Cn�bYݵ�H�C:;����3~�,��u�ڬ�Уr���%�������~i5hJG8�C��of����jzj9d�2��-���;���V|�S�lR���]r�S��0�����͍��K�YT(jq3�t:$���~�&q��Ab9_,g\R��g+�*�Nh��נ��1<�.M�Xm5�iG�����8�p��+�Qj�x�᫮�<J�������ܗH�g��.���su+iO�h����`�"��if�ߋ-��;����l��ƥ�hx+�c��{�`d3�L ��~l󹄓�4�~�V<�U�H(�m��k�%�l�ϼN�+�BU�nwJz+�U����m6���X?YǱ&Va���!��B�S5�K��~P?��*�����/VϪ��
�i��UÆ�t�Y�T����cP����ܸ�Յ����Ok��MRVa�ȳD�|㬓�%��d��$��;������D��"���[�c��/��=���p= δ#d�m�V��U�Z�~/����yJŗif�0ծ{�Y9'Y�9�����&��<�!殶��v^����P9<�<�i4��RӾ�����	��z��U	۪�߫l7f�/Kf�cG=����P;DӤ�	E�͒�*+b�#6�F�x@b�YS��>r�{Q|V=��R	;n/muh_x�j�b��3 �9���.�b.9$ig�hvSVD������b"��g�-�-�94��ac!ʓ��Sf�f�Օ+L�<���T�4|��?&ō����t�g(&%�C&Y\�i���͉�\�y�OSʭ�@`}a]��+9eYXWwu)��G�^����]:W)�^c��W�����z,�'Y���d������0�Zƌ���>h^������&%�����2�t�yr�F�A�9�ķ;��?4:Ѭ���ǝXnl<�).�.���"0��,-���ŉWFR�዁tH\�Q=��َ'gR�p�&`=z#����I�ڙ�e�ă?f�
�a`Xˬ�F-�P�|��Y�Ɉ +�^��b-jz���C�
U�I�xַ7T���R�z�C�u�Y��^���vi�m2|/��PVm�)�tx\�����6�X�!�M�N�n�:�K��B�!�
֭a.d��5�a�*y�5�:�]���%��9�nI�:~�gfuP$��R*<����ɽLz��>:����w6}��j9	�A�=�
���ʒ=�ص_�N<�4�Q��Q�8���KY.����'�y2�Y�	+���y���a��?�`��R��1�H����ddĜp��+7�.2]� ��W�Vu:yFэd��-u��*BqY�P9.��׵�01���4G�ϟ~��)�<��$q�(s�&�ӓ<I�H!M#o`~��2cf���M%�8�-3���<��(���h�ݽ��Ha�dV�4#mx��)��=�5*�V�iF��F�4�逫�h(q���ҡBd6r�r��.w��+?1֋�幡M���H�%��Y�0���d0�Ф8�>�d����^�^g����\��HY�D%�lR6K���g�Ua}��)�X��I8 ���F�ޞ�>��C�,�1�Y���8м6����cn����.�5<�sg�l@��!v�fH�����ƣ�{M��p�w�s�ؘ��8��v�n"�N���=	�1���(��u���T&P�)|Iθg�a?n���*~�!���U'ALh֝wW;�=�'ko�G�3R��LFZ���H׵�F�(��61-gFy���߸]�w����N��i+��T֮9��1�S����3��KGW��b,�v��\ۈ^Q@�Q�A�|��7GF��R�cH.��X�%)%48�qY4�b�U��1)��%����ʱ�4i �V4�LkuQ����̾>���xg֗�w7�l�|>�$TA�ԉ�����h(�~�:!����@]��MU�A�]��i�^�t.�쯊�������p=�O(�}ݿzhrw��[:��~p�fW��5qQ�bB7�1��P�g�{�p���ϋ�Di��E��ڐ괬��5A��H#�T���Z�Z�h�?Fè����9L\�xM�o�g�����r"�	"���0ݖ�k��Xi8'_T#�y?y�5��v��|�z��`�{J�E!�]i���ԡn���7��@Azl��'�[j��a,��2V���h	���L�烬J���Hݵ��r��t�@�H�f4.M��W�&�]���z��N���7y��&�͛�G�t���.E��kS����Q��:�TSQ-�t`�h$����ȚsF92/J�zZ�����o2h��ذy��3��9"��@�S�Ȇ�D^b�V�pZg�x�Q��|8c���E�YT�#�7?'��C�h�\^󠮳��w_�`�at'y"���# źa����B	�^0>� �?᱊ �V�/r������J�q�8��ZB$mǉ���4f0S@6�p�s�7{A@�j��p�f��w�4ظ~#
/�=�Q��7�����b;Q��wM�~�#h�n��й)��A�~~����43��:�#��%6����g��,��0K>s�ߢ�vDw���'7��m�-��\q�C}��ۦI�ʢ
�6[$�m2P��6,a,��$Ţg��jf�i�����5��~�?}^��ry��PQC�I�ۋl�I��WY�$l������(�(���5|/ܫȿ���UWC����F4����(�'�t�w9L���f&E�$������ѸG�i���� �����EG]��;)5`,�sSc�膇��+#�����И�ؤm��8�CO-&pw<i,&�����9y�,1	���<�
3S��s������?|����C�8�1o��Ls�Q��1�#�:�$�%�mG�����<���k�߾�1�����q�@#nEU9�]	9�"��C	=��l&����^����;�D�����2e52W�}Urj��)3_�!d��u�ּ��ٸ!b�c���z1R&G���<�rݷ5�N���u��3�j�e���9�$^���l�XJ�U{ъ5�xcf�n0�ss��.��\s۵\J3��Ø�<����@�89����m���q�}����z�������#-s.������S��6
�%��.F�y�n�ǡ�瞢dyN*1��2�Y�k���~?���.O�S��`��U�!6[����[@�
1N��_�x�\Nqŉ\��є2hgvΡ��T�s��}�gp�Ol��]���	�/�ɻ�)֘���Y
�4~Xd��/F`c�@��#�w�ϧ���hr,��P��̚��0�ǁ%�NF���ڥ�g�m�J� �~�9F5;$��]��ҥ�WL76��:\p?(�z[�<���6�a{]��Z��Q��j�b7�X�]���5Ny�;���(�L�k�q��E�2����Y�S��8ֽ�z����J.([}�TݔP��"�RᲚ��g0�T|RE����	���@'��|����a��0f%���TS��YE���$��:�4��$�Fت�Q��_QDbC|߾A��m�N|Xd0�h8�l�MǇ���%�K�����kܰ?��@4U�:%��F+M�R�0y��%q���\��?�>�B���V����>�n���1ҏ�=@ևR+��{n�eN܇#ug��paE�)�U(�D��(�?������{�ͽ��6�7�>Sȸ�t�[��!J��?����/��~�Y�8��,ИXzf�?1��S��	(������P�|O�u]��l�x6V��KV5'���
�_Q�1K�f�mbd=bH�3��:��STcy<�߹�U��NIu׾@5Vi.(8��:�R���D21���m�c��T�����T���-Y��<���Z�W��488.�3�|A8׈ς�2Z��\l��B>�!ACZ����r$HV��*ύRq�Y �??۵���w��e������|����ϥy�ল?��.QZ��I�g��.�ܜ�\jM=8�
�ߠ���J}p�Y�E�8��F�x6_�7��<7=��p������
�� �!���A��g�+Ӡ�X����������}�n���Ǳ���ia{�w�Y���_b��z�@�&��f�w��u���<s|��¹�g��
���r�u���!��o��cR+��ѐ ���>�(�n�ϰ*�=�ߕ���~����O�3+W�a���D���լ�!�����L	�1����g�J��>]���wE��k��xFs�Rlr�L�����X��@R|=�y����X�'�\씕�j�fIO�Ľ��1��hj��C����/	�Ovmܳ���tM*���!���?�k�F�,;����KQGէ�6a�j�J$��_'�y�,c���6R�Ikz�9��`�w$�՛X�.2��n$E Ս��Ba�	0W�� ����G�U�zzv���6e�VH���)êo��!3fw��6�RЖs�8���9e�x]g�����=��x���"c@ Ģx��}\�߾��j��F-7~/ot�줢BP����Ok�EA�d�`������
��qEc��C��b"f��ms������8��S�l��A�8����x,�?��?5?��8$0K甍�c�+B�2�Y�S�N�k����jҽM*�TÍUB �zwc�@.�| ��_B�7��_�n��'^}��h:֕�qy}ג/MV�H��akwwl| ��7���g�����YwI5���|��3�T�;�7[u�EW����%S�,F0�.6���c������W��F��~G�aQ�*F0,ĳDe��#�q�G��{�
�P�M&��X4k#���t�5�d��Ȅ����T�����l��2�G�pH+��*y�D�n��pp�H
��+g9�dGv;�O�@I�����C��Tc�i��yCyHFGUx譺w�ZcSgr����r:���X(8�%}knd������75GL����|Y�`T�z�46~X�_BF,�zTm�6Q۷3/*X��0B�bx�4΋(c,�m��,�!��3��[פRF��	ev�ۙv�=�s�����3�ڬ`ڒmj�2<�#�nW|f���Ʃ���y������9@LA=_�3=H�k�g����wYJ�I��.2�.���GY�iD�F^�����>&�`N\�
�*�d��4}/,�� $�1iQc6��<U�*��N�L9r{Q��� �t��v�g� �S�fH��x����� �ٿ�Z��]��@������ � �a�w�A��̛�q�<G妜�I��h�]�Ls� �W�z����� �2�^�A���w�lZI�i����:���u�>��R:�>,�ǐbC|�ݷ�-`�����L���bEF��Rς-�L�Mՙ;whw��Y6�o���8���� �g��� ��mt��f��u`��S�휵�Q�3��=;��� ��1�9cZ<ὐ��0�A��il�G/6��,==���������o���)�KM-㋱��=|9r��*7#�w��V�D�aq�h����2�����ō	��>|fo��vʵ�o�u�2�1u|ſ;�O1�`�ܜ,�8�3?g��lM����7o"Ƿﵫ&߷���\8\��p*0��u���A��ˑ�t��F��_�=r)o33<W���Y�#���K��&�ۦ�����+B�sc�Z3'���r�eʝ!$�3D:��D�����n FQ�!'>H���=�'=k�ׁ_���cNXH+ɮ�l�\ }�w��H�iE�)|��8#�Ƞ�/�axw`]��UY���Ͷ$�S7qcQ�"+�����w�'���`'*9������q��}R�h��!�Nio���ܺ|E;1�0pZQ|#�DF��tr?�,�Xl�J����3o�m~���tDv�Mh�����ɺ�vlaG��@zHɨ1%c���EC�xe�����Y��T&xw�9��SP�s��R�X|��j����u�:������m\H!��}?��J��>E�,���;S�8���ӡk�/P�G���� Ɵ�����US��A����h<� YA̕��c|�6ȱ�l��]ST~K:�S������{xwwUQ�s^�����d��O�T`9�fُ����v�~��<�,i�9�ye��_��J4�<zP���j?XS�V��tc�
L����>臡���F��w��$���,��H7���o`��Du6��o4&�])�t[�U�%��â�K��̍��B�(�}���\O�@U6�y�����O��D^�=�jŕ�si;��M~��J=Q�ʼ��\���ܘp��t
��Ȧ- ��tJ��R-cD��U�|]<ɰda(�BJ)=3�I�؞2�K�����PAi���Q�$Ϲ���\�>�N8��c�5��g�A�j�t*�YӖ�Q��!���a����>d����+�Cs����쇾��׼g�fY�e�V�a Ҵ)v-R_6��5�q�l�-�N6�I�2�9�
I��iԉ���ƥ3��W�tv�g�5g����Su����*����[���d��u�����a�书�e�H�}EoE�G��]��"9���n�d��4��T5ú[�~3A�U�k-�������k=������i@�������WKҷOvܰ59o���kf;���Rqh�!�Ӝi9=/ݍ��v�Qvb��?��f��L��x�k>�5GU�z� ��ӟ�����.���̔N�ũx<U%�>�;�\�/)ر��o�ʐq�]��1�qId����P�	��.dʖql䜒���c�7�y�>�s8���P��@s�B��]d�Qht��מ�x�6e�)��Ý��WS���
��H�AI�T���qlu�+`����@!��)��ԂL*\�|?:��t�2��R�5�o�<����*<��h\�{�t�9���]1&4�6�+V�>g�Lt0��ᚇB��%��V�fPQֵ%��I�s�Xm`=`�(^f�����V~�3TK}�~t��b��T��R�	����vx[��T�R�b௸ok�D�3Q�u�}���}ԕa��pFZU����w�������pY�N�:�^K���B��M��ۦ����W�ZP1��Ï�@Z��$��� �R��21f5�Ƅ�|��V��7`p�j�Xo�ԸIdB��;�s������ �	av�kL�x�%�4���Eg�����x��x���p�Y_e����f�H7�\��!�G� �30���Y `T���}<�_P�>r�ߗV�eΖ���2��+��3Zn�$�[���^l��n�������}��铍��<Ϗ1����9���ڄ�h ����:u��؄�QΗR���`,�ğ=<Ce�D���	��^���7<����ZW�#6OQ̀1�v�)�Oy�~��9d����|��6*��&�s��c>;|�y�+2��S�K��Wed���h��ˌ��t�@�y��	�\S|���'TQ�M�C޸x8t�qH_&�%qcO� \0�<7�+�����_���0݆�p�{{�N�R�h��w��}�|����m�d,�����sL<I�6�&ڄ��+�uu��H�.��R��̉��o`�?�̙0�r�rY�H8O��s<�i:'�}fz���>&>��T��+`!�(�t�3i�����?څ�e��Kצ�q*+@w��E�C6�Ω��������g؂�g	-K1�5����W�u��/��v�	�AO#+6#T4OO*�Kw�\q�\t�o3 x�0#=�ZLoH|R�=�dZ�!�Δ��"���˹y�ԩ�>�z:K=p�!d�p�tq��V�C�|��93`�Q4"�8\nb���Yd���L����V��B����ߩUx��VP�f5y=��$Ok\�m)�L�z8'+`�/�}<��X�̀�sc�Z���єH?$t�f�]����+0H��\��Y}��@�ۍ�l��Ou8p#�D����s��6%!�M��w�����yF��BJ�J+��n	��5�a���fa~8a4��~֞e���o�~-��&��ɇD6Qxg,_��ùEGv�A��e�xmQCN8)��d��A�9۽�x�A���e hL1��aF��?S�f�\X����:ȸkZ�	��׍��o�s#�7 �gQh��# �Ok\A�Ԯ��39)�k�[����s���1$FxR̌�s�|`X�@�6?s����u`yt�31o����߿�~\d�lqx��������w�b�1l�B�R��,�%1}�ZS}:�wUc��y��&�AⰚ'�A���\7��૔�%_ԍf	����yj�ck����vc��g!ue��vcj|M��%vs�gA͊���4A���k��Dg�<�o�z����$��}��,�ss������͔ں�,u�:��՘p����/�>m6�14����i\�EL�E0���9j06$p"�*�����#��8�+��M������ت�ى��*��+�ill��h���Mtp�w�aL��3������������7�va3�)��s�`����lW���A������[����.�����@���gq������쎂P��z�f|��?��YOfCs���]\=O'P)�N��"��>��؀�ϹY�*(���E��D񷡞����9-#���QLV��@����k�����ϒ�sR�2ci����v�@yZ�vئ��`�2���^|�z�����N4�@K����GO� ��b�����̍g���K� �ذ�Gs���@;WTaN\��)J�IJ*�d�
��~6��
��T#]��zV��A�%���4)a��{�sM:������.Sa4�:���@�+�O��]���`Q��$�<op�����*�	A���'g�2�B(�pb�᫯�d.����aY�k-����B�2�3�xs!)�$�櫚0�΋ȼBN.��C�� ��?D6���,��/�����Y����^�)NamU�z,46Z=���:���>U%�
�s���E%�Ͷp_7_n��a��_~�%��o%ǃ�G,�������h9����Ad�ܩ�r��6N�a m�,�`Қ?/׼JV.�O�|e�L�����Q��Q��F�+���
��o�����k��~���u�^xvo��A�!����U?�j�<U��Z�,zg�a�jm����-�a:~M���)�i�����\6�D�M�*��I��Y�ml޼~��k�����؁��J/��|)M˄a*>){
�VK�iJ���=a�s�����X�'P̙�8Su.�Ԍ��.�/|��_��nV�Q#*�k��Z��d��/�����7_!��{���5ӥ�I��Pu#���o��vZ�G�%g�%�O��4���^w"_6R�:��������j��ʇ2����*�N��]Z����Y
z$ç�}1���,!)�]Ӕ�u���86�L��������#�n��q�Z��k��g�so�Q ���]<��3��nP��Sg�vI*��k��P�����3�M<��1�3��[��9����7�x�2�f�!,Z�-��,�a�}�ЉCF����lVaTU�􊢴��;�Q��\͜��Y�^�u 0��X8��YS�j��ЄG�v!��Y}ч�~\�2����F'ϴ"nU?U��ke�0yv�X���?^ދ��q�T���?�5�C�T�Y���&��JYf%��q��mq��_�޴M��H�<��F7^"�������3ϼ��F�D�諮��273��@Q��T	@wUVfd�����9�*I��2�����3��+=h�,�tf��qx9�
ㆌ�TT����d���\������AjT�(/u�����������s�繜43E˴�&C���1C�{�@���`lE3e�5�Q$l�a3�OY����y�3Tz��CD�� aT��3R�"f �U�lQ�7+1±��J^�_����H�Ya^����e���snTm'{V�QJ�,����q�ㅍ�g|9��^�����ބ���(K��Tx������v����q�_�Y��c����Ȟ=�
��Ғ�2�/,���)�-|�C�y~�Sx�D�D{���-%�F/�3X�@0Wp�7/n�3���d(�s3h�vS�ʼ���Ȼ���f��x����ja�	" 'ϛ��e�fn6�����ȫf~:�����������Q�uqq]S^���$��ݷe�xëP;��=aMk:(S^:�Z$t�a��<�a�\��^��)q4\��^D�
���_օ�<�<��<1��d�ڙ�u]8�������Y����@q.,���&�J��:�+�-yu�w����FF�&ԳHazF��iCp{�Y�$9��-شBB48k��	��ث�1������9�Z<�vb���uB47�ڰj�;t���
5�10��D	5.nvVe:o���O�A�YȤd��& ��!�|!{*�Q�]��9��/̗���Z%�R-�k��N)�,$#�[u�)(��������9���U��l��$��>!w��W���x*�j�XOF!d�f��\�����TI�J���B+k�*��N��a��C��V�9{�.���P;�����-ͧ���kl]jcI&�b���QlӔ�x�=��[;W-{Ѧ������=��ԥ�|枚��T��4���_�ƅa��H�n�f�e�rF�#[V�������u.4�֡�58����W�aX��p��2�N4��jz�1�o�S�����&%��ū�l+�QL	p���˙���غ�m��C���+o��
O���W�%����f⬲���#d �ք�+�!6M�h���?��fC�[ukdOx�!Rr��Fd�*��!
��b�c�����&�����3ϗɱm|v�尗�
�\:��KY���g˭6�[�%����|������ oG�S�|�Mк��{���'���٦�<���z��˄����!ڥ�Y���>�:�A��!E"'���&0n1����! ��9�0�u6�mϋ7�.:ֵV)`�����û�w3��}S�xP#>2G�C�
�zX$ɗ�p����.�(ŵ]���4+�����.��@̮�\�,f߸p�VL�{�B�!p��)C�z�4�MV����X%��WiR2V���N��:l&R�"鴰�[��v Ī�ڵ�0�� �sb!aA���|G�k�3�e6/��aN��;Uuj�	�w��!)lx���L�	z8��^��gс�k�9�*l	��y��c8��L\�?t���úby�H+d\�:6��	�_PJ�~���uL�2�F�$��X��`��`�34Eql
W�g���Gs�:���h.'\6ROg��ս��R��}z����+�4Ա?X��M�愦H֖�X ��s����ً�'�9p%1�Cx�1���ڪk-6lz/����yn�'A�;��{�L��F��ȶ(BN��nY2D��$�hs��*dS9jf�Y�9��S�s��>!�C�S�l]1)�,�1�:>˔`�)Q�B��m���
�۾,�:��sn �<���8�-nv�8�V'.��zuba�4��X��~�Kc��i���x�����~�E	�ޮ�U�xF�m�E/��$u�Cb��1ZHAn�(l-������}Rg��!&bC��V�!0O�|�3ͪa_�'ɏ�%P���sk_��*�c�Q���>tHI�~������'K�O���u,�ZE��?�׺iʧ����ں��&�i8�z�s
���h;�e�6�"�ҖUG�q�N61L{�c͒E�'�$��t�+k�Rv��'&ux6�� �wֆNf��A�~z�}0 r~��ދ��>M�8f��^����6����������F=0<0�o����n�1���P���]SWT��o(�O/RH��m&�ʒcgE��o}�Ǐ�Vp4J�j?&d;1N�a����)y�I�2�@��vR��J6N�����t����Om�5 V#�q���%�g|��2��	�?�^��9�J]BDz����e霱6�)��M�4v��(|�x���3�X=�6��G�ԩ�'�`�5��i�5�����w{`���z��Y���og��E�푾 JP?��˯�� jQ'��<=�PӋt����#B���U~�!��$	x�����TIA*4�����5�{���0�tg��M�R&��m`�~eY��ҫ�
',Rb�wz���Ԁ�:�f8Al�^]*iy(V��B��ob?���x����P����;�c0�-ϗ�I�N�2s[�eNM��d|��n�ǡ�)�@s����t�ӫ�Gj��E��9��l!f��D�h+�{(C=F��C�/��ۤ犱0���?ܪ)E�y��HY�
�Q��!4��p��F�w�#��O�j�ٿ�	;W�A}f��_�:��js>x}�>�97���I�O��u�"|�L�G"m^B�0�s~����tō
/h0�q���懓M]9�a�Xc;IM�y����<��{���$|{��"�Oڙ����ϡ܉-A6�?|��r����|v��M�!b�N�%<����"����C8�rᛱ.����#N�����@R�!��:=;����h�dIP~��
K	)w	�c%[�opPWrԶsz&.�m��2���0;����uL��Ͳ���d��BV�E�7`���t�m�׺�^��!�'���:�Z�+k��q�QR��7\�y0M�[�
a���a�꦳�7��\�Q�M���B��ѥ�Y����c7
c�M��� <y+R��~�ǵ�,��}N>m�5qJČڶ17���y]$��6vsN���B��
�x}��Y�
q#��?�v,]IC5���|x�� �#�?�y`<�n&�;�cͷ�
��hH�r��ܤp��3��p��=�xƙ�l��]��C�-·9ڭx�Z�i(Ð��i,ٕ�6��]��&��4����"'s��*���gA㨶�j̆D��B����*S��U� �VR�5?�<= '%�Y���k��"���TDb�]\�!�c36y��/v$׉[��b3I�wV� �k�F������z",\��:*W�ǒ����{I�$^�I(�H�_���%f'R�ŭ�t#��� �Whª'�0�����7���ز�ay\��-'�BS��c{���p�,�Ɇ�zI���q٘o�$"! &B�[W�jQ��阚��!��a�0t��N�lܣ�֯_�$�4��T�Z��&�B����9�9���}y���|���/J���Fϡ�e��&dU9�S�qE(}�"#~?w:���\�qu�M����?�K	�Y��
lv�VЂ،9�T��⊠F�CN�E�6'�Ӽ�$.�؈�F�a'�¨��Έ����D��F��	��+�=f�Ž��j�qAGؠ,�hŬ�bf�^D��[��d,?��~��?P_�#�\/����CR����{P�}� <���������F��u���1J�v���}�8!w+x�]f����C+��qg���l���>k�h�����j�48ie#��=�~�����x��
�ii/~9��$N61�m! ��F�o"�����������ڐb1�ر��m6������;D�z)����Ƭ(�}҆��{s�p��@�Os�ڑ&MG6�y���l�J�'�����C�=�C��>���X$��Lzα������4�����GxH���`�+���z7�k��O�G|6�~6��Mr�!��.�����U[�V|�8��J��hI�X����am�)���!��3oŶ����K@�}L��F^3��P?�j#��H�w��{�_ڈ^4�!Ǹ�*���! �>���1"�\WL�cӗ���<�Ļazx̸&~<˓ۋ��
�ssK*��E��k��ٷ����F/y��B�R*��7��$CO���$Ey'&�f��ʁ[I�s����",hA*�.��;������G�p{��/{ʘf4湧�}xq0"�e�)� J	�8IԮu��
�E�"��7A�Z:�=�����=���?�9��KB�4���R��4�r+%a<iH���U�8���������ur-<Ү������(o�xF�Bf=��|L�',p�0��RD¸�����a�J�'��,-���ƽW칅g�(;�l���(��MY�{悥�u��c�㧸6<���{��FLx ����󰷇�����K.x�8��M�]r:q_$g6̻�[��4#e��8lwF�%�Gy��H9o�p���ԵC�Z�����^%eɞ�<7�B鵄pD�_^�/�{�x�~��X�Dt�����`%{�}_�\�\��ց��g�������-�c��V��M�\�]�D�z���(�����:|ZjE��^p�{ka����`���t|�}ӟ~ǉ�Y���fV4��H�����<��3~tƬ�_4��b۳͒?%~����P+#�����bW}|���J���I_���}�u��lw�����/����p����Bn0\0NAΎʭ��2n�&W��Q@�#U��� ���_�3�Q��^�w��1�w�U�կr���$ak��x���K�tH���f��;5�;�~'��j�#���}nL�|[舙hOp&�h��ś�S\��^[��:�}��p�Z�^�z�s��8�Ɇu��3�#�����B0��tD�z��q�F��g0�Pu�H�s���|nx��y$,�|���"�����6���
��3[���s��3�p��i��y�}�)kM�ڜ6��Y��J�Ig�C~�xPB����N��M��s�7>�v}�	�(�ё��
�	�k����L���>Wb��p�]��ui�)�gt�DD!X�
\�������ipNx���e��?����S��#K���#)+
�u$����0t��.�,��Y'_�^Pi<]%^L
��T�~l�l��0�_[\X��=��H1���� ��+g���Y]�oC�Y��<PS� �{d4�
��5ٸ~,60��޿̾;���8�}r*��y��Y�ܧ �cr���w�V�_U�����ۑWiO�"�̺�MR�p8:��!e�z�6H.�Ov��s��(�8��A<c\?�@�p�0�Ѹ��N�7������p��y��qk&��>�u�y��q��[7:��pٔ��*Mo9-\t���L(vjW��}��=�e����?f���-E\��m�k$A�
�s7�{c����7�>��t�X��S�xb���Z# ǋkJ�1��O*� ��x���d��T&#�����i;ȟ�j�<��>X8�29zҜ���f���t��t�L�C�S8�O�F߽��Y
0��xi��_�5��B��iH?�%�YW�ᬋ�iR�"2d�@�n�ޛ��^0�l�J��.�/�6���|6T�م���7����ɥ�!�ǈ�@�ʿ�뿖����H��w�zo
���燞'<�*B<�mh`HY�|��(-���v&�s7��s�/�8����?���.�c�,���Yp<k�V��[���Þ�O�
�>EΞې:�7�a-Bǚ���!5P�hV&�;��	�)6��ۘ0>�0���q#ևMx���_"�v�Fa�����T
������%ädU!�^�0��-���0h�!�|c���D��o�(JR�~�m��w4����`٬�x�k�k� �������>K5#d.E])������ex֧Iz���	����B-Cl�Y0�;fy�N�u��W������J��Y�4f�;�:�3��%E���Z�Z�d F�O���gF�Q�J�+q��ݻERSus�h}�,��.g�iHO�4���{�<�_�C�����f�M�n���-3e�wp	+u�Z��풡��n���G5��\m]�=���:P����r���,�v�+���XE�q%S��ј?==�'�ٛ��!1����.R�rxd�'�����>����@!�R4�L��g�o%�8Vs��9�������+����ů��'s�g�R�H*	����4�e���.���R&�o�#~�"�lV8�^�}lf,~X%���a<
qPZ�6ϕ��)u$��γZY�5=�،ѓ���j�0ޞZ���)�'��ߵd��T)�����k$s�@�EGu��n��.�&�w3��Y�kVߊRAd�*�]b��	!W��eC�r��9�ÛH��9�ZxO9��C���$������ؑ=ĂB���f�Y�]���k��?:�i�t}�M���j��bs��wŨ�_[����Z�̒K���ͼ5_G�9w؍A��Kd4���J��^�?���p�����N�VIQbjOV�ƌ8�V7�<��BɢPY��k��Hz��~{#�T��>����#�2�O��p�mL$�S1T��Xôf�9Fx^��k�n+��6GiJ�Au��7��U�8��]>�r�x�m�6�΂�"���-���ׯc��0��.���`H��ѕYg\�FtYx����]�04�p��GUU��&�����#��E.��Ԧa�ƀ�Vv ���[���Y��Uy�6�}�i�pe�BS��1>_�1Ⱦv��N�\�Qt���Oɓ���AB��C�z���8>j�����<��HkC
j`(��Q�Wz3e_�57G9�O�xZ�Kb[N�I-s��u�Jgx���6�I�`�x#�dk�:�(R ������{�Y��Y�4���y��]�Ǉ��E��zld���b���8��8���0}Av߻��a���'�hX����� w�=3��)C��<9\�C�׀�~�؄3�!X�]:	���Cx�H
�8ؔh�q^x��_�ބ�|���Kb�y�E(O����>>�H�\�K:>M�؋D)+6( a��wxn�;�㐆Tp�F�W��s���j=���W=�y��Pa����*:�J���uL)��18��G��w��}��> �"[m���3���9������x$^ѽ��e�>��"TuB0���
�Ϛxl�L�n�x�^	ZYe�?W3�V��s⩧�����UHC�7�j1�5�������b� Opb�ھߗ,�h�7ʀ��#9%6��3��-Pw��4'%�R����;ʐҋ��#�P�@ϯ�J�ׂ�V븁Dq�iD�}n�Q ��ĵ�(���������}��Ҩ�U_����v�	�Z����qK<���ڒ�S	M�!����/�M�{L.jY2tv��:7sy$^Ȱ�C�,�y���ق�����G������TF�u�ᑞ���'�`cpx���pzw�H��[� %�u�S�1�������S��IM���)[�Pq�}�F�^��|E��L.\����j�	:��A�<Ր������%��?i�U��'9�,��i��+�f��5i:�� lT�/��^���:��e�L��ފ�{wR��O���u��M��{x�a�T����I��XZU�Y"��ͺV5��4w�E�vA�W��a���6��m���ʢ:�1�K�Q�|��v=p|���H̬�1�����u�n�HbEj����0y�� �
�M�Q����k���%%�,W�W-��s�7��N�NԿ��8^v�G�4e���e�S��吶I�6�?�V���Ϥ?�hN2�j��R��(\[�vN���ߊ�K!Ȕ#����5$�vl�l�+��K�$�f�h�BayQ���6���~�m����j����
s0�Za@۫�e��9�'MP1p��1���'���vL��(��+��r���4���3�X�5����&�N'�mc!	�
a�j�&(����:���MlŽ��v-mB��O������_��Q��S$jH��(Q������e�&���$ի:�43�}&����8�C2"K
��-K�u�'�H΁alLp>$��+��	�Q|S^'�w=����!��Ƙq��gG���g{ޘ��Jؠ7�����7��>_�/1n���u�#�j�={�A�R+h�=���G����>$w�7obְfD���&�_���Y�	B��S�#��;e���Ny��qp��jdwS� �����UHy�=ϸҰ6�i�觎�H�Z�̈������J�h'�C��^)xB�|Y�*/��Q��Jmy�څ�$i;F��N���	��N�=����Q�6V!����ݜ����.��@�p&q�O/��M��t)��O���ł�F��� cf��D���|N�uqia/��j�R��k��ժ�)��������*�ɞE������Sd�7�,ܐ�^���8w4������ ��b!�e���MUו	�ƻ	��H�&,̱�@ϋ�4�)a��rx��^1O��٫2성b�8z���%��(|<G<�,��L��v�+�]0|�bH<ֲ�0�6��D*Y�غ�8��"�l�Ĩ|h^8��0�N���0P#A��Y�F�ȣ��(����{�a��Ο�q�7Y[�����W��P%����%��!�����Y�f�Q����vS�U���D���))N�M0Ֆ6A���D�f���"�vYj{��!����i�@b:V#ڥ�l�#&�� ��{���-L	��m��T��+_d���Ζ�,�"cy���9]�y���6����I�QwJw�ă =ɭ]�W�M��l\��r;Ff4�qېz��l��������0�`Hc-K�S*���;>�	��K������m��SLث�N
N�!������|�<����:�(��F=�ߖ_�%ƚe��u��jH��}80ׯ��*
~��m<;?��6&�~R����n�
�0O��������"׻G+�ǧ�.tF�z��H�ʻ�:�+�(,}�ถu��3�1�eI��G]�e�x~�N��W݋���T���W�?'x�_��B'y�e�G74
��MF�A�M�����Z�;�%1v�"#�S�1�*\�  ��IDAT�#|T��4<+��_[\y͒W�p:�N����b-����<��y�'���>i>c,\�����,K�d(c#:/<R�����#e�ܗ��Q�z
OUw��F/��=�0��6�ւZ�T��E���h��܁�	�� 5a�6�E�uYc$X���{��M��d��<�m�����2[�!�!��UM�.N�6��S��(Ʉ�r�I�;d�6��������$���;6�,)�+ZI82�Y{_��t�fi��@���O���W}�v�Gy�6J~lb1Z�!����̎�S� _�W���X����e�xƥK�<�ua�Ӱ�D�t�!b�W5�h�cx�������^�&�$�l1��$yF
>�+�p�.ѨP���7Z/j��0rY�=�<iE�w��/�������j,n��띗ZU��Zk~�*��ߍ�&5�2���.K^�8r��u��$����2*�kDv=_�[Fc@�i��s��49��x�Mh�MᬌL�S�S�ޙ�Ec�h�k����kz���.�e���~�;�kQ�ep�Â�@����1�s�ȝff�fo��Y.�;.P�������Z�ϐ/kh*���g���Վn:�:/U@b����+F�/mc7L(B��ɲd��j�9�ٓG����>Cu|tY-�=w�u����{��<��1�n
��?x롶1������I�	Oq���
*G�!rB2����>F�ޠ9��6.fɍ�Z��V������ўm1���Ќ�������h1���K��kR;�Y��'{G$m��ɶ������C@�w���ï�c��9�Q��"�/�|Y^�=A$�0�U��$���R=$'���ê�>�~�8�LC8�n���p�y^���? �d�����"�^��<e	�F����'�	N��?�ujS@d��׫���"�Y�]UeƭV�Xg;m��h!���N8�N�U��.�=	�*/�5g6r#{3�'G����������6�ɡ�fxN�,�4Fq<VQ�")8��b����}_�wm�ZN�)<J�'��W������r��ަ`�_�5��N!���Jf��6~k����NaP۲L{eX4nǲ>f�Y�x��^��rEQ���n�ʄZ	
T����~'�VÐF�z�a!�rȅن�T���И�ziT��K-`܎����lWV���}��!�B5����,~<��s39-�aoƙ����)r��֙@���1��S��o8DS^F;����+�j��",3�Ė�w�%�x��1���M���/���u�3;9����S���1��x�==H���JT/)�s��ج߫·y���D�������1����؜8�NX�y��}��J�eͱv1�O�vjn9;V|-j�E ��P�vP�L�(�e����?��Y�ȕ�7�ƈ�����[��:[Q��(f�	6�k��߅��O�'�������x�wu���E8n6�����bń^��\�J>��x<{ gån����M���A|����㨕9��[q��V��D��i�;"��W���&j��m�b���A0�[P�־S���=���&���pʼ[O ^M��+t�(ٻT�
�.p�_~��E�$4"L�G�ؐ.)H-֛0�7���m��1��q�&f���y� T�m���&ww�d��*�
/g���OE��H��X8�
x�G7_S՛���[8����o���÷�r7���Y��::���g���S>�AIU+tv�,�����^��l�����p6�>���2��S��-�=��p�����M���^�Zwj��SSAl�ߤ 8˯{)��>c�\�s��T��Gm��h��LVA	�9v�H0�P�������V
b�E��'�qH��W���Ԉ�j�@��8��b��\��F�0����g����1����1�=Y���0�cN��y��>�hJ �|GNx#n�Pq�)@_,ĖZ���[����𐱣�/]RS��D��#
I	5�3�������~�L`�r�Ȉ��	���Q���̥g�Z�Q�h�{o��7gbI��FK؄]{y��.��,� �e���Xi�`�1����0�-�߯r�p�sxH��{Q��$�QY%��Js�Df�|�~�8������u��m���!?��[wq.|�5^�h��E�j�K��C̛��l|�W��z{6�f8D��Se��Ð�yo޼JJY��n�L�M��Bf�	�E��:ot��P�A�,�8J�f9����q�ដb�w�6������&������^��Ý�ga�9���K�2ꤡ�7�$�I�9�b?6b@(+o��r +9,�� ����D"|m�}h����� \8��_c����-�$�+:4N���L�j#��1m����G{H$�爨�R���ܠ��!���]\�J�W��h�Ti���{���x)���vN|����G��jw���]mGڄ�b��Е�����/�oc�-ὓ��k���z� �-ͅ���ED�$�����(&�[	lDE�L�4{ۭb��H�fޞ��� �H�F=z,�f%xf�+3<]�ӖI��^7
ZS�5([��zm����$�&oj�D{��5�n�xL�%UM�ON��tX�(�Uxn��'6¡�K��c	R�3� �ީ�5�C��v{��aH7*���}O�lH������ta7g�Y;ǂ�^l��4)=���׆��g�T[����������^eE9B�c�R�ׅ��wGO��:�+�z]d�#k}w/j[~�gI��MR�T��T�੧c�
�Oz��ӄ9t:f�,�n43=ϣt}O�a�G͕ʕ���#�y�N���>��]kA3�� 1�Y�)ְ)bv H�B��ӺT"Rς���<�rD������{���e�nb����=#�V��<��}l +m�ﶎ��͢��=�Ih��Z��q�/�⬽���ih	J�/xqWal����� <H��\f���I ���7�D�s�2h�oq�K>�e��<��φ�ݯ��#J'��]����/�F�t�Z�ͷ���(�S�7x7m��:�xO������x{}6lq���!l�Hx��=�p��Ja6��؞����&<I&WN�}p������[��0�!*�wՉ��L�mE��B
C
oH����I���c��?��H]�����
�N8^�_"�q>���/I�:A�b#|?|lc��p���U3= �$y�;$����O�^�Rj�`�5<�ׯh\#4�R�}΁��6��B	b����1�����J��z!��	9����H�T�q�k���k�:= ���w2js<P�&%�NMa=!yd��KL�t��q���HO߷Y�@��������Y&����]Ipg,)�ͅg�n�8��Xv1��agC���iO�<�k*ʕ��֨�9�!#\+���{�}b�޾
|�p��eAh�Y�G�𮧽).���3�Y�"����s���;���_6�'c�a�N,w[z��W,BX�*�4��׻�w����p ���~�79gX:��^���N���9CTa"v�l�p��j�M���Q!z��W���A}�3�����5�>V�������B��ߵ��ko��ʹ�$�G/�/K�\1U��g�)p�&�Imp-�+��
����J��I����X�T��0�I���TQ�Q��UO�}��ە�*[�Ӡ
1^;9ʆ̿$�Uk�-�����^+�K�6¹��	JV0U,7*b���{z����<`-+���ی��}3W_]�x�A�7����s�>�a�s�)GS:5���I�%7Y������W�{z�-���h^9,V��^4w�\ys�s���!�m�mg'�mEe8&M0�R�J&�;���Z^S4zJH��˸�g�o;U����F�S�=j��3�ȯJ:W/�΢�T2~c��x!��˗��N�"��<�����}����QC�i�\r��0Z__�4^���Z��AF�����9L���S��D�MC��4�ßib]��9�w6�Q�¹i���W2����%JH�<�$��A*0�̬�+��$�a�	0��+U'�����)��l4f_�/���g5�vJX��2�A�JB���$������N��ǆa����> xmG��z����E�J���b�����]�o»��E�OlN�1�Saˉ����]�C�1h�T�I��]�U}��<�	Qa��[K��V�3���kh�[\��1��+��.>gXƟ�3`, ����9.�ʫ��fo�j��9���ڃ��=�����%�c����t� �.�l����yc��oazw�]�����,xbE���H:ME�5��s�,�_�ò�������Z��??�g�c|,�ec�z�ܪ\2f����H@�E�&oq/�����^�Տ�t�y�}���
z0�hP%A�]y�E�p�IJ
�[]E2��UTX#��K%=��m��ڿw%���������s�*%�5�\4R��{��2�L�u�����Y!��
��]��=dE��_����taHݣ�5��Ɏ����=����z����n��>�b� �y��U�����	È�8^I	��,���s%6�V���N,�jo,�R�viǟ�^�~�&�^?�Ա˞R��=Hպ�������G)�՚}y����{B=���)�C�f��Y�,�xА��'��b���7�!;EL�̆x,"�'r]�e62�W�*�h"�S�	���I8;me"�JO�nDd[F0�Nb����ؗJ_�N�#)�7:�'��W�O/Z#�c4�ѧ!�bsws�h�x�}��A_{6�d�-X)�u8gN�9:y���[�����ː޲]A���4������ ��#= Jˁ�y�1OO����r"���|
=��ߩmn����q��2��D���gA	��r��Ԣ�����?M$�pf�C�˪�Z���+��n+o��*�)�u`򀒴��m(���7a\p�H�g↳�� ��W��*V�f�:�?{�meӤ�k�ժ�|.7ě�)iR�Ԯ�.�mȽņ����/�f��,�<KB�3q��Nm���y���]�fs������Ɯ�@�Ø���@�����G@d��e��.��wL<�,�gJ#���v���G4��׫vQ%�6G5�c��5�wV=6�ۆ'��8QG֟qT6T6~2cf�ɘ�z#-[&�!�RXB4�Ԟ�'=������F�B
�l4��4�Ϲ�srq�ui��-\��x���)a.b�N�	H	��t_�r^��-X&�G�A��������֘~�0\�w|�gS�f#|iփ7Qgv�;��xK�2<웋�␺ �t�:똸%���~�	��AA��\Ðx��hO`���)�����Fa�v�s���2���x�i2&y���+u�r^�eNo���W�\�%��ߩ��	��{U�P��2h�%VJ��c�	�_�8	*3�P&n*�m��7&�2��D�seuǈ���R�k���c���;q�8���?�
Uj]
�HC^�y`P���?������a�&n�o��{l��D��\��\�׬E�WBԪ���흈��D#a��k,�A����3���ae�6g��z���n�����*�@(̽�J~߾ߧGm��k��5�B�)�xR�P��6�V\r,�[ZJ��3L��t��q�Z'�`�n�)"����L�a��[m:q��~���Ԉ�o2W�k����Y�]�Q�F�+A����z�X�]�(v�x��)ۆ�Nb0�̲�^�� ٢�"�PsS]�!��V3�Q�p�J�V�yjTV������Y;sW}m��))�6��n�㞽����:ra��j����J1�~���^�8V�g��僾lU�Tg\e��DlS�[��u�a���Uj�����a�w�Y2�$�R�����t.>�d*r8�S��Fh��:ذq�#�~ ?rTr�%���X�U�K��?�;$?��x��AX�A&I��~��&����-a�Pܯ����1|h^D��[I�H,{� ��z(��+$6��1�BX�[� ��j,�f%�v����h�`�vsu��Ҩ���T�����е�u�����u%J[x��ǅ׾<tKB`�w�� ��$�А���Q��^�e�x)�f��{^=e�)oSHi-=�9�	C Q�)� �����u�^��FR�,?�~ʈ�}������1�?aF/iQ��L�Pۍ�wq8d�8为�J��!�f5%R����6pV� ����CL�t�� �uJ�]�*�G|��`!`�ms6��B�ºU�i���h����܃�=��Jڟ�I�9WV�?�����08�X\ ���:�����7�������J�"�u�Q����OC�L=VnJ����i����\��v�(�q��U�=7���!u���aCꌆւ�H���{�Q9�og���r'P���00���"<F���$�*�Y<?%�`,�%x߻��v���nH�}�M	O;.��66ni!��n�#"%u�E��iO�s�߁���O?�����(\������u9��G۞�6����raQC9Idz ��E|ǩ#%u�Z��5o�6,���w���ĵ���u)�l��{-6�1DV�q=+�T=O��q�wmD�ɺ���?�So����PȿTL�G8�1���b�ن,2p�"MD���1)�N˹��M=E���bu ÏʲZ�
�xH��O�^Xd.���je �xw]���iǝ�u���#���ޒrR��j�Љ�B�7����
���1靭v���!��4�C}�
y<��%&(�D�~S�94^'���cq�PЧ�(=�`91�g"�Ԫ�4A*^���p�JDo��ÆP���(O,td�^p�����	�M��=��-7s[C�ß�:#N��xA/���+���=#F:0�����@j�����T"jQ��u��"W�ƀ���y�߅��5w������2��z��?�JYt��?��tkAN�4<Zܳj�h�3/1T�)
W�>�1�����3���T�N�j�\Ga[:u
h��}N��s�G�"����!����ɠ�aχ�b�*Aw^o��4UN���{aJu��.��W_h~�"1�������� 	�2e�2��+«����ċ����i������K4e���a�%��jA�+x@��}��mϵڬ{�_Lrx1�$r&t6X?|�cx~~��d�Ub|���㝌�cY߹b;���=&D#���UJ�n�����	���%B-C�1�uC ���X���Rc�M�O�8rGV�=7��mFW�����3?��S�ن�F�P#K~�Q��B��P
�!H�iι�bR>
4���J�>i_gX���]_��"��A�w���lz�����>Y��lr�69 
��2��)��R��gEa�L��d�萅0��@☞�U
��;C�T�P�;�[�؅Wy<d�u`�á��7U�s�c�Q�BB3���x��X\,�chì\jU{��~p��cG�m+I-%��1�����O��S�~~���M��`�4DU���ou�"+Cٖk�Þ�[2`���}Ho����#TB��X 0L/ϓ��o�_��/!�*�_�=��۳�6U���D�;y��^�̰�*8G�D0i>d����\jH����s�� ��U*���8�7j�^B�d_���sx�_��Z~�����/�J�X|�8����h*�T��[��ܪ^�ի7g��FE��e��!��Qy��N8D5�X<l �7�$Q�f=��'�&N���f��sa7X�	��z��eN]�ˉo=Tl,���Y|S��=�y#�i����x2�D��/�=�Â����'6�����0�0��}WWM&d�,"�X��h�(m���\=|>��ꈾ�Q��g�09&W�B�rr�qu�_@�p�I���A��f�ͪߚ{��xV�?=��:UN�Z9�(ȗ�)^��=�G�J�L��z�k�Π4��.����|���"����:6���f,�?� hs4ϓM������-��Y�Fk�掰��vc<4�٪{;���8� �-��&כ���ӟ������(�q����&��	���R�wP���*!O�
(�_˜'*u�қ��Ğ�)O�J�h��SU��y������˯�~p�,�J���?�!�=�V|]X�6�!�U�lo�=��{�����P�w�(j/'�����.��v�%�^��p��,�wYj��j8��j(H���kzb�a�����⋒�����Bs�	c�^��*3��*QF�P�е�^�'�S���Jd���#\�(J��}?�ǚ�o��N��y������%����}`�����Od���&�r��7�����@�UĢ��ŒS�hJt5V|��I�����0k���
��êO�B�xHƁ:���XK'hq;d��H����e����PW`�	�8b����6����n��#*/:\at.9z��Kבk �6ڧ-���u��co��������1��ͻ˒ڤ��E&�S��+���#v�S���tl��G		D���0Qs��΂+�a �dT�C�)x��6��p]�_\�3���:H�xR�zj2J2���Ҁk)S���F�jN!4�ݑ;/{R���)N�P�7���(���%<=SU�{��.R���N�X�>K�I�̳�o��g������gV��$v��/+}x�x^�.x�~/%=Y��F(�D���+���B�8n2�>Ӷ-1$�W=C-ЪV-˒���P	���Jn�}@�����}�z�i�ʠZl���g����k3LЋd�g4��u=|@<�k�WH�`�㑡1��OU<�fp��=��K�H|�h
R���O��3�����ؿ��)�n�8!�t:RM?��?f% �hb�Ɋ�	���z��;�*:��d�^��wj�'��&XC:R�-�<U��G��ڕ,,
oX	U�x����?{t�	}�1ӵ��}��rQ�խaY>�^9R���,w\��%�յ�{���t>��8��˕BAh?�?2��8E��{�i�1��B"��)�c&Ƌ��*5K,$�p�4���7�R�)�a��ٮ7i��Y���"S�'�W|p�)~�\�gQ	*���0K���>�Y�0��*(��b��҆�<������`D�k5�^�Crc�Ɉ�k�%�h�⅊4RwWXH=�p���~�-Zͱ��%_�z#��?��+y��>�0�]b���Aߒ�6��wL����dV�ͺ.�fw��køU���+җ=Sc����(rs�P�=�a��?U|��~W;9Z�*��ȕR�GzL��j�&��{SݘD;%�MK�g-J�zw���:�%(������J7�D��f&�"��:f��v�vPu���:�� ѐ���8|ɋ�<�,��x��
�����طj��ğ��E���A�v��S��}����4�Y� ����AȐ�/i����Q�<R�BaJ8�I�_r��.CZJ��孄��nČ{��~�wUm>��¨Vj}%��C&T��6'aH;?X�tSb�6���	q���A'��D��uŤ��B�^6�d�A�k�"n�!����% ���	�LM��j�.Ѥ��O<t��C�a$6��i� ���ÏaHq�֗�^�jl�	ho/�=�[@М�+ M�U������!�`;Q�6���:<��Xy��z�QJ*�)l��:�[X��LR����DH?�.�Wm�Z�JR�Ϫ��z����mt����z���gjUFG��#���9���_5,�h��jۍ �Kb���lq�h�B��b.����u3B%-��V�V�U�}:;l�qG."���yL�u͛�Yۋ;��bq���)�#��52�g_���sU�|iغdYl�ѻ�Y����8��r>�ի��\Ҡ.<��7@ՖU��J3�N���>e�(tb259��IV'W���@��M�l�YB��Wz�MB$��WמRo� �ը���cw�'x�I^{!����wl���;j��IƦ@�`q��jm��T�$R���ך��mP\�	l�ݴ,�k��/Ta�W�E��H�D�<�����.i�f*'��������Э� ��8Z��Y�V �dXUi+m�'5js�N�"ʉ��&N�1v�O�Ns��i����4pc�5�gO�m4���.u>c��[k��qs�LY������_-�go޲W��{�r��U8VQ��{瘙RD��j j�4_�0�!V���R�T?U5,G�lO稗A��?�@;�<+��OT��ss��E��f�	�2��B<��wh��>3�%�j)õR1m-v����/��˄�?����_��$T�M�d�n��-i�����b�|���͝����lY��fi��c��P��+��`����	�?pX�$ȓ��"0��f���RK�ξ� �튻.�)�{v�^�-t���	cm]4/���wV(c����>G�����fN��]`�F�7�o@2���< j����^����ȋd#�	B�	�N��1��mx�䫂�c�d�����Z�w��܆���n��nj���ޟ�E/��ۓ������Ǭ����]���}��#F�<U<]s�2~nx7J���+��]�MH�/9.������@ev�3�ctr�5��hP�������J7Jn������0�!C��P�T"f�ip�u�
Ǿ�q��09�}�37�=ΆÀ�}R�0A�k����e�_����g+�b�c���3��]�麓q����/�ѕ:��x��:?��s�5���������S��<	*^x$ލ����d�(#4�z��O=�uKf�X$�F_��X,*Ró)���!�g��mkHC}�<���ؔ'-�Nٵ1&ZYJ��);�+_~�%��KV�����Ґ��aR;�9H�Z�>�$& D�q��)�r�>J7af���k��6ɡulf�o�S���t2`�?��s�����!�� j�	,Ӝ0aM�!f�<�Bڮ�w�F�D�p� ��1Rh�H�<�)0ޢyG�@ߧ1u/=��_�^L�����
V,�vXLL�z\d��ac������%���ۮ���2�hpna4����+AmB�S؞�����L��C�Y�ǭ�p�w������P+�0�'�`�u<�6*�(ƛ�=K\�%nCR�b�T���2��X��H�F���� �m����ƕ]YG��Q�yP[��i��&��X��a9ϓ�z�n.�(9������s���c�JT��{��$���G*�k�.քqL&�٩<�I/~���d�&��b��	�F�u���8v�ISJ���W�r������Z�*��+�J�i�P/6���L�y��P��k�M���Ťps��o0\��=>��8��wY��hQ<*Q�!u?�Y�?����] ޸e[�mo���!�p�&�.�-���p����5�۵�=�>)>��������8C\�l�V
Y�&N�&���u�
���5����k�]�9�%������a�c^`�Y+)HZ�-:�̚��1w��b� '���v&0��]p�b��̚^��j��/Ƅ7e����ɪ��˵�QX1Z���bݸnY�����:�~���7���qxNm�9D��I�,4j�B��{�ӄ�vZ��O�c��F-�T��1�%�z|�z��(۞M8b<{ZϷ�/M5��]S��Ŧ�n����-|������ր������%v�נ��ؗ�q�2 ��^ ��{69�Â}{^�V��FWȌ+���g�6�&8��i�,�((I�~�^<�c$>����q=��2��p�e�ɐI��L,d�
����b�k�^���F=�4� 2�0��n�|h1�j�aD<�]��K��G�7q &�t_�a��9�ڂ��n�.юE���]���3�^هl�WڊB(�m���]��`6l����	I�~h��Z&�{TLysa ��e�e��"x��䢂S<�h�|������
g���a��?W�@���unzl��.=� q~g���ܨͧ��;i&t�^�d�A-�Ik�,�����veу�:0��/l���@ ���J@T�¡S!������8��D^8�� J���{]zf!6��D���*b��X.�Z��T-mq��V�]���Z�*��f��+5��>�]&}Qn]*�9�Կ7^�9|鑦�O-�m.���"�&���^�]���ʣL�|C�6�!&1fCWJ���?��5�/��>�iý�!}�6�W�'���rt��#*>6��1�`̉_|�D��	I.������$�*M�υ`�����:͒�P�u^_3��%���F��ޑ����&��	�����<)`Ha\.�р��]a��$f��dޥ1�i}�K	���A��u�s��:%��V��Q��SŊIzw
�&.���� �S�����w�}�{y��:H|��h���"Ď��ń�Qz��7��ECU������:��3Q�U����<!�׵������v
�Ǳv�!_��b*�.=�w.�鬀��٫4� ���\I��l�,�(��z��N�̂Ȩ��OCJ~rm����(�r�z�Pdg3Q��sB�]QݰnJX.��.7�e��H��la�y�3���\b���Y�*�j�>��(�����@h�؝����DH����yW~���^F�/�?���"�K�6b?���!(C�O�%"GB�mf�¨���(�0G��:��\{o��U�H��aD�6PM��W	���a�!��]�=���U��<��8����=��u�^�������<f��a����9�C`c-^\]䤋���"NLxӬ5ˮ�c�̗���w�V4��v�1&�8n�=�QO���0;#��ڱ�~��ʟ����/�����ߟ����%j�D��-��ya._ebf�9��687�mO��W���7�kH~Y�X�9'<��:T�B��X�qj�Ԑ窱�6i�(+ׇ��?yУ��E�k�cw"�Џ_��C�ψ&X߿.�Qg�#K3K|�N�-Rji�Q� ���!�?h�j�QUB{̜��-�5�;��X��s����pi�z�v�@�ȱ��'�~˘ڑĿ��xn�iHm,kVIF�|��c��Y80j�;y�s�9I�ng>(5YN<kTH?K���_��؋��]�.�;ӫux:��P���,l~�
6�-��p8
;�'d̀�锕@�-��Φ���c�x1�l[H��|�S11܀����*<������ۼ�mtZ#\�ï=)-��q�>�GW1&�z�6��R[cL�x>��&�&��Z��;�9�$u�T������ ޤKR׫J-�r�qx\#6��~$mM��FԼM#w��w�1g7�u���d�1`��lI��S&jB�wm���Z���0��0dnC~{�u>��1�����8gx[� �4���5d���DQ'��T���rׄ�t\��a9�+
B�e���i�ޚ����z���\�0iL�3g�m��cj(16��ѝ7ݒƽ��I�����fz�u��j�����9#<m���w�G���I7�X ����Tt�Ĝ�9,UV�J��MOJ �Yx����Z;��$�-��`�Vg\I5�e��x`7L'�Ԗē���ڄF����]0Bal�^QG�l;��C��<�NG�2���6t��á&S<Y\mj�CM��Q���>�cA#���~��5���9�4P-�����<`D��@��Ľ*�XŜ�.<_z�OO�������!q&uJW����d��5n؊WT����&y���2$��>>=�����My�S.F㌭�8�}�L�ʬ�7ShlD)&��U���û���%���@��Rb���MR�t_7��s���)N-�cQJn
�Tɏ���V�Hr��c���� kh�荺?(�D��]#����\F�tvl�F�,ʹ�R�L��
z�u�5�^�,�3Ų�Z��5v�1�=���Ο-�8���G�Cy�������/�!59��@o��3��%�kV�`p\�B����c*t�}I���䬊0L�G�H�7łR��4R��؈�	�,4Z;�p��c��Oj�<w��s�-ʱ�l|đGz��&�צ⚵�o����S!���s$[�\���}
�.�"��s�q�΍�]AYx6P��Y>0�	d~�"얆Ø���hS8��|�a�e�M�m�}�0�51����cR}���"	ջXO�L6���P���.� �'�yK�!h��ύ)�Cͥ��(LI��x�M���v%��N��`�IX�4m�Kr�������P�W[�͈��&>g�P�H���4E�Պad���3��K���N�l��f׆��MF7�w�JG*��<���:[�x�Ш^�~��+���B��g쀾���{[��)C�)c��7�l>J6�*'[��R��8ln�U���n��s	����Q;4��м�p�T
� Y�\x�7��c}������ L�$)/�ΞH2���#�0�q�P��Li"p���^�d�eV�t��Ŀwݓ@C���>~�@ӱ�cK�7O0�)�{1��az}��0�I�P;�O|�S�k�,�j�%�[��wݳ!o�mi\К����5n�w�Ħ'Po���eN�]9[>�P���8�����P)�g�89�[_TY�8��·M�B3��)�}�=��s.~|���cvZp�i�Cw*�e�͹u3���$˨IۧQ�<h�]��߻���a��������yΖ���jIcc��I����N�#�m�`Za�Jw��h���f�KfP˚�gZ�;\��0`.i��
8MtL'�tݳ��L��kD�Aȏ����S������E>���t����槉�����b�NY���+�H^wC�X\'�����Ʈa��[ɼ�㸻{�J�&�d��V(0NXP�
�7��Nl��#�d�S'n��WL$��A+j���h-�����k��n>����g!�$�9<�q]�����*���>���������RJ����k%%#���<�ΕB9c���'�ŕ)4�g�>U~��3���B����	*� �dfx�l}vYq��8�S�\؄����8Ϥ��s�w��{��c�=�K'�~�)!"�NDW�n��!�A��rb�������>NI;k���^�!�!�k[�Do��N�� s�4!\4Hv��!�ә���^�6l�1�`r�EM��ԧ`UݦX��etNl6J�	m�Ĉ��ƚ[��]UI$��!!3��֟�%;���jO�y���[�:~a�筗�b��1��.x��9�&)`:�'v�����U�Y:�!r��u����d��T<:�E�?��hMA��jCi0��B��u�y��� ��"t/�Eą������cx.m�����5АSOs�x�v�
����XO����U��%�����i8�%�V��[�Tȷpnbbh[|6��AõP�������4�NT7�;ȣ��$�T����(W%��)$�,TL�k-����C�c`ڛ�=�>cc��<6�s��Mm��h�Rv��gV�{��\���抱a�����w)F�4�ږ�C�[�����6�e��.V���5�W;��	={{�^S6��v-�c��?��� ��:����R�xļ&�3�)ӐVV����ۂLUK��e�JW1kϝ`H��m?�Dx�R�7���B:�$ �?ƒ�+a�}��R0Ț�Mɧ��Z�2���EP&wO4�p`x?}&�ξ4�S&���e}iħ*7�܀�8�7�6��QF߆���
�l���l��4j�B���q	�7EX�hO�!<x`z�-��f2��`�1����>�w���x	�&w:L(���G��̷��F]�_�믬��f	jx�3CkÚ���c��j����hX��&,L|�>�)h7xe��U[i�N�8�s�_�����ĳ|��#�������4&,$4.����g��C\� �
��Uo�?߮(�a��8� 	,!L\D���i e�4��6�g��B",s�w�i�Gj�%�N��W�9 �Պ��d�E���P�(����F�����՗���<>?�\ņ�{�Gj���0�/>%�I������=:{�Չ�^�;�:i�*//Jl�P���Y��d�a�h���[�pVՖf�������C�.��J�7iY�S@��_��+�P(�lOl�����s��K83�A��X��>f��J�R-����=6Et}���<�\d$9)��D�&�K,�&%1u��~5�4њi�-��O�i#Y�S·v��d�1�g4Tъ�v"᳢�\x�np5��y�Þ��o\q-ò��Wp+�Ns��8��Yn$tb�ܞ�c�&�`�/&�"��n7Ys^/�哕F�^Zks�UL��J�dZ��Eo-���W%��s� ڸL�����5Uy9f������ɞDr���I���	1���Z�.=agB�0%���z�V(CB�ٙ"Y�H�I����}[����X�)�I�<�?׉n��,�,���l�k�4^����}ɤԣ���ƍW�NDm��Rlڰ�1=ρZ�nj]���R;@��!p�=2����2�OZWmrG������^�|6���5�(I�E�\��o'��'͋��	��oRs26=�ٰƔ��
q�V��ܐ�F�sc�i�%��r$PΝaH�)bϳ��#�O�KD��H6�՞��+��B�+=�������f�:�Jt(Y_��XZ�]Q�!�t�~�͵X#����'j��*�%��o7ۜ������#C�٤Ҹ7��9<G�w��E��J����g��]���$T��pت��T[��<ܠ|�kj#�q���Q��u��8:|�A�C��-�*=�넦��&;�z�r(gwj2���]���8�G�r]n��C���������'�D�����A��V�L`{��m��K�>P�̂=����d��@S���OY��d	�x'�j�)��ߺ�ƔF�%�W#�$�d��/�z�+��.	Wd�>?�iJL��6G����z8�$,6ɞ�-���ܐ����!���}ØE6�6�Q��+��j���0��n�ס�V�����@bh�oklS�P����>a�`�`}�3?G��}�6�2�s�jU4
�M����?{4��K��v�Ն1]X1��7a�5�޵��c8�"t��[�ͽ�1	Ri;��zюꅷO�x��Hg2��Fa9�QԦ�3��7EX�������s�2�ky����)D�Z=e"L�V�?�%ӊK'�*��h7�k�V���aJ�'�3���x���?�|p���>1�.�k�ö�=�����9�����|����0`�J�kӤ��E��p��}��Y>��>�_m�c����zn��-5�GT�ŔΟ�S��7{��Is��:No����cR����0w���"4��N�e�A�3I�U�qt���⇀��;�Ic��
ٸ�	��&���V�a�Y��L�+�vx���8�?X���E��so�Rc��}-63����h�2�u����l���vO���xu�D4]��_l )��2���#�ǧn-	'�?Ҹ��%�r"��+��Y[��4�V����L�;\\I�Ek�/w��X����vCM�[����Y���R2���i�;�K�R��4��&�ۉ�� Wٚj���P\ؒ�aJ�I���j��,�o퍆!�Q{偍���5��ԭC��m��fL[O����D2/�_�sLd�]�f�d��će��cۆ�ٳKx��>Ss8G.���6	��Y��j���T�ۛ�?�b�"����ʉ2\<B`�B�ŭ}+�~^��z��G��:4�K󻶅t�w'8�@~у�J-]^.֌3�����5>/�4�udϽR�H9�I�vw��R�d���G*�
	�h���@z�6"#�`NA�,9���a��ب_8���1������.ʴ�?���c���w�����r�bH�͍?;>��3�X�Bkh�%EI$g��
���|��>4q�O�Ĩ�'�-(�c�^e�'}'�7�{��P�ڬ�m��~�:�K�����B%*��/�]t�k�>)�:7�j�� ��[3���h��ᢗ={q�䡚�`|�����¼�m�8�z� ~�I�a�n�-�a�KY2n��{i�\H�G02�*+�0�KÉ�=}��;s�	�}�̀d�6�u��vW��s{b'C�?$�`�����-�^��?U�����e�}�wr5����=c�E��X*]K��^V��	�Y�:-��&�:-B���0�J�yCB�m�L� �]�Aޗde�����%ǒ��ߚ9	'u����JnE�.��c�\�Y��1�#��t�A�zڦ��Sn�|pT"��1J"�R��_~M��9C�<��t:V'iY�ʬu"�?�_��\X�&�R��zm6��<4&��O����P$��j968�z�L�;�'UR����oO�أ]*Qג���~PT��d��X*4M��<<�L��>�+X�O���5)��mJR�K<W�7��{��v*�@g��+!_���p�VV�>_��\G��r:���$0�.!��ʢ$��I=��JQ�mfg�G,P��!�>��(�C�I
я�̭t����:�Df-8ˌ�8Cq��&	\��L0͙h �p�@�ԟ1OO�}-͹9�}�p�c�䕽GG��D��9���ËԢ��rb}�"�&O;���1��]k�>�Xd�l*o�!� ȋ�Έd���P;8D�4�jϿi>;$�!j���xմ�a�\�u�."lօu�֮[�L'��^9�꣇(�èdߨ��Rۍks��,�[T*>=�w�4�+���b8K����v:VC�?y���3.�7���'�WL$Њ�`�2���c���1����g><�Ա.�*]f`S��U�A%��_P����<�p�׵\�a.���~��ߣ���؏,,��}z�Y8=R�+�ӄ����6�*��6��f�~�u���Q��Ami0Lt�rG��rU�ɩ����V��8�K$��i��Z� }H���s������t/�k���#U�����H�EZW�/p���00��Ə�i�ᑺxW*-�<�j��d(0�Yu!�Z�5z�M��TKm��T).Di����4���҈�5���KE��'v���c����oYN0��YRh/,}8�*���v�굧Ę3RS}{&���x$q�9
&y�Ĵ�x	
5�P�Sl0%��p��[��Ð���0���^�y.xܜge�}o��>`�ḧ���������|�*��pS�/(��Q�P��M�ki���z�ckG���kr߄�"��v��z���;+_��kl�wY  J	�ZԠ������;@kZSM�$��ةK뼛�Ђ�ɨۖ0B$�NS���=�����XrQSL�A��}~6��=���<�j�;��N��C�X{������b��n�PIlR�\M�Y�NgƝ�6���#���r<ڶ��>f,ϛ�#
}�9p-���(��ņ�zv6���y��l�l��>6Q��zM�p��7z��ڴqGd
�y`�2��<€�\��ax��x�!;qa{!�]U]Q]�Q|`g+��1O�������D�=g������ M��]T"���&��<���q�P`d���hq��Z�;td���MǴ��W�lQ���g�NI�Fx�}���S���9�	<߹ψ�s8��ߢ<�������;��R�Yf)E�>�J������lU$(��"z������0 �dzg��X��(%��+)Ҙ��dM�fWĘ{�_2����Ō��v�m�v���j��>wk��ɂkA�;*���'1�5��@G��k�SI���c��A�o1�9���6#��9�B��:z��Hx��׏1@&��26LiIC�$O���"�� 1ZQ��Cp�����3M-���O�9�_��*d͔ͬ\�W{e!�!/�c���LI�����%���C���rzOcN�<�1���>ƀ�dW���4M�dO,�[�����\�<đE�_��y$�d@]d`ʞY)U��C�z�Z���Y��\�Viar��!��9����z��I��0Be�XG�+�\&\� 9E׉����u`ua�Sץ��1������Y�^����%��߻�',��L]��-OaHƧ�+'\��	cI9, �D]�8�{c��b���	��Ѵ���PY�|TJ������S��VMG�=Z��b�-���h��>5�Ƞ��!��9��	o�c�8�g�����&v�H1v/T:
��ٞ2Ѳ�Z���v+Tq���P*�*�˓F�l�M�a@��a0�n�N�}Ub�m�M�ǽf�xb���<�"�k�ǡcL�q̍�] �d���5À",Cś[�X�����4�T�YCF���r��-O���m�m�s������Z�,b*=������ʐ�f�^�xޥT� �j>{t�Ӷ�B�W���IZ8s)��)ф�tٮY4��k��Z}�&��i�l?��uz��Ǥ�!"�<il��SW���d������F~���'1iH/5��n�Z5��z��8a��2I�Ĥ�aD�׍�I=ۡ�����^�o%���6���t"�|�U���T!"��At�ͮ�u�8�^�>e%�e"ϭ�t� n3,�����"�;��h-��	�SS��Dɾ�P���x��Č��=t�W�1���?�����J@OY��ɓD��5}9�Y�g�92أs�k�b�Xe><2H��lD�}M-,a�7�b�R����'�
 �5#��PiZ�~�<�3u�����=Z7��
�-1
&�g��Uc����&X���1�*T����S
U�2l��n���^��mH��)�>���"#� �x\YV���OqXN6B����L��}^��c�p�.�����h!ɸ�jZ�Y1l�^Vn<�w�غࢤr�RrZ�+p��E����׶
���P�ŷd"�X��ڪ��̅bG���Ӑ°G�c�$1nBx�������n	9dc�F��~�����?�=C��8��X�!����u�Jb�@��oܺ�֢,��8���c�H�{�G��f�6JM��vZ�yڱ���]����(�P���f����W/㦂�DI��I�"dΎ���"��E�M{0���o���5����b�b�vʕ>O+�[�] ld��M�P�x�K(%�օ�c�g�&s��(���u6q����`��#��w�WQm[�T����eJ\���՘�cV�g��Y�o�T��'�Z�ܐ쀷}�g��{�{��a��<�B�*>R
1eg�����!���5 �8e*��B��vR��:���"����$Wi9N�y>H"�x_5���=�}EU��.�	jm.-�fѼ?H����UM��_�/��KۛhIn$I�f ���L&�LU�]=�o���d�fgg����x�yD��-TUDU�Ar��:_0"#�p�z��H� c�-�Y,^�-P'ఙ<�9n���
�C��!��F0���F�2gY�;���
őI�'�^���ŠtL�8�;�1fC�0/d�-<'x���%�g�ὲ�����0���3AVÓ. [Ԋ5'��#��'��qf&���,+�X�u{�%9/)V�6�;�����`{��J���7,taJN�s���9�F�b�K��XyD`j[��~�V��ƲN�%�W,+=�~,檎����*��ǇE(�� ��$���Eƺr3�;�x�l�p�v##����c�z6M݆��HU�۷�csZ�M�	��h�\�?<��9���h�~��{��s�J���-��� #A��~���EAC��l���h	��2�s�..0��/A���JLWc����|taʲaos̰z`����PL(6C�r�VU�áB���'�5� ����.s)!H�HQh`�iX0BA*p�Px��� ��o�����gx���$s���P���]�;;��O>��F0Ut�������X�V�$��h��jޝ{A��`���\�HJkݿ[�L�k'݀���e5��e3�%�"e�ʜ{�T?{�[�����Ơ��5���&z��4���� M%w2{j�6k�K�
#`�H\ͤ�['���	�j���#?���wa���"H�$�kI�`ֵ3�����V��;}�����7>����=Hh��z$dD�a+��β� ��<���{���Ԣ�|�}v�ms�VɫW����:OG�� �,w�N�˒�Ŵʴ��z���J�������_����FC������=�w�X�������2Z[Dh��#w�$ԇ�Bo�#�'�9,OW�k�N�Z��B��������[�����%!!�w�>z�_>;B'$��FV�ћ���ͪ��Y$Ĉp��b�G���)>˵'�}�F:-��JH�<Ú��D�u��yB���/�
x������3@ѺS<Ql�=�����r_2�T�FQHO�X��)��8S�&B������	�l�f;�ҙ�M&G,�� 38C�����VI���K͸�����U�?���O�U��L��z ��֨���4�,�,@��c���.��Z�����r4F�2Ff��KN�ΏYЖM~�n(/�%~�����F�q��"��Υ�q�k�U\/<n���{���ƌ��N���rdǒ�ws#�.��i�'d[Wv�G` N�1n��ͅ}�_���U���ug���Q)�I�uBbg�{k���ap����A�Q��{��`�!\(���z�����a�L�@2�& L�,�^��ك�y�0���ғk_�Z��o��@5�>Y��iã�u3��`b}2���!�k&�!�ҲX�Iaq�`��8�dT�߰9j�>d>ڂs�Pĥ!|e^�2GͿvG������G(о�A��aߊ8�o6�r�L2�)}B������-{_�8T*�b(����%��U!y��k�s��r������K�|��>d�:{�ó�;$Z2�_}��
G	�u�q����[L�L����n��a$����,��j�I�����m��b��p��l��
{�Jz%[G��+b�&���ȧ5� ������wB�?�����v����*����MkBF�v$n<�u'���h��{=��Q ����][��h�&h�5��Tm���M�_eװ����2O����R��o֗������HY���-GKDЛ+�ݬ���M"&I-��o犕	5q�"a��H��=v�,x�*=F����}��o#�`T��Y�Mt�#�g�I%9����^R,��3���ֿ֢:�{�2���<T�jJ^<6)����|�����VJU{^�*�Ɖ�:y�p�G�l ����`b��ڸF�� B�ģ���<���`�rl��4�TCG�A�����L��Y����_��omS�˿ڗ�-�;m���{26���;]��DK�S����
Ɵ~�IaK���ɻ!�tg��[�7߁2�Ww�\����˟��'=t"�=p?~4�$XP�7F`�\��FID�̢�?�`���{��PJz>�}L�,��q'I����T,P��m^\�i�R�;�B	g��=�A7�T���#�R��1hJC0�:MH�D\Pvu�J�p��DC������d#ʆ�t������sI"L{1I�-�"�N�eiĜПK?�� G'a�A��%�hF.#.��g��ޒRl�3�|դ�,�s��;�
���(��]wy�������^�'�<����e�=!��n}������0��(˴rYvL��4�����h��dY�h7�ϞA��k5 ��T2lA�<���t�9��@�X"�}�R��K4�<"6:��ϓ��^�J�a���z6�M��4OΔ����}���^z|0�ިxi���&c���X��ͣE���A�Ma*F��A���?�Q���o��\�A!Qf���G��z�>�`�WK�mS&�l�M��f�nZZ	��9���zXXz�0f具�֬�����`1���7�}����}#��\��,5}�Aҫh������0��\c�C���#ɫ�z�s��}@��Sr�f6�0�LN\�;+�T���,�rO9�����&/#��xm�	26\��Br��tĳ�=��*���^���̫O�w�UA4G������g�B=؋�{��;iZ+�{MY���T�H҉0
P�p�;kX�����Q�?��N�&V�0�5�UE_T!Þv;4 �v#�����{���׹�W���{Of0)ֽ�-Kj�\3�?�O->Z
ɷ-�`�y��YA�|97�1� [�x6�z��}�	b����L��A����ȧ�$W�џ~�E�����[9�!
c[Xzk���հAo]A'��Īo@|����Ĭ�g�&�н��#�l����m��~�
���:B�b�ko��h1*d��q�&>hC�TV6�h�����Ou�K6�%0n=�C���va�Z��.�n�a�-x.����wj���^�a@}�$�8	�+>����H�P����9x�^G�"�T3�u��+M��b�R��dB��W�l֧Ÿb�G�	T��`�rH��8�F���O6Y\�쭐-����R9 ��x�$�b)E�������xWX�c^j��~U|��Q졋!�yh_��B��B`��X��L��zz�L;�����?֊�8A>���D
�RBI����;�c_���*qL�2~��qo��!K�:i����C1e�o�p!��ք��(]���B�h�̵�a�H�AE�W���y���G�;m--�Co��M���'5��SΌA��Z�b���,�#p>�.O8��&�5����y��b��č  =����4X�D�+G��G7��?]{X�� �{�������VɑJ�լ���+��ēy�X��Ԣ����1O�G�4Zyƅ���������}<��0"�	F�]����:ks�V�Κ�����/�Ю]=A� B� dURBZu�{��$D"ݑ�3�,�l�(Y\�sl���hTp���mJ�����i����ŉ�p���������ʶ����,����$H�ZEVE3�@�;ͯ36�Xu^�<F�56i��+�(��8y��9ؽ�w�Dr�7��m&hX���U)9[<����/q�3̆�֖�y�Z�'���5� Ʉ�Q� �H*6�L eKY&�r?�A?�axI)��<{
�ц�#��%+�����$L�wc�j2d�<,#�<3�� *�s�-҈�.>v��Bc\Yh3���dq�������'����軛u�ǩ�.&T	��^/�/���f�>K�sQ����k�/bŶ_o�p[���C���\s-��.��� eN �S����7a��Y�����f�}	GځK] &A:�t���lG�����1���2|��b��'R���~��>�J#���#F%���%����b���_~�I���\��Ɲ�I���(JDE��_����ʵ�|��33ky�]��Pq��g��!�EW�Jل�`$�T����Ųn��c|�j[��JP�:������϶����;�� �Q��p����CD+9ן��؆��ƚ5.E��z��2���7H.E��XEUѼ쵶C�3Y��=|| ����4�=�L�ޢ���F����\��2r�l��$��d�K \^*xau�Ⱦ+��*jd���Y�f��)R'���<��E�X�gO.��U6�"�	[q,�(�Fu�u�_-�����@Q�k�zP�#�c0�ת�ޡ��G�i�Y���N�{ؙUJ�m����5����q�a�5+\����5?u��y�_�{V��uO?�9�	e/��u��V��yX��{cθ��k�s�m�t+0����^S�4eڡIݔ����*D��f؅u2�3�{����O�i��*��T6���"�Q�Niٱn��TLQ:
�l6�h�����s���a`��V?<Z�MBs���D�YZY�h�*��^jP��z Ѳq+�7�r����d=jp���v2����dC}��ԧ&Z���r��NYZV��Fgj� ��ϫ���̀m˒V�h+�����$Ðl}r�������D,�x�\Y7m�}CaC8EH@�ȋ�~� ~�Љ�� ��ג�	#0����,�*jJ{^ѹMH���BZ8�.9���#F��n����������[aa(c^ܘ���!�n��'�N~�[�P�g�v?�e��(*��u�}Tc� %��� �c탊�+���R��D��9�W�@8�2e�O=�dY%��Ic!-���Xn�Sĳ�C=Px��d{��V��kr�4�	��H1QE��J=	�Ń�:u����6���ѳk,��t��^���KT��`ت��|τN�dd#�� .�|���V�L��(�(`q�<��3ar����V2g�$&~�j#�_���"O����8�|����h�G����ߠb
�A2>&��g��g!���b^;�v�do$@�P����9�a}��Y�Bd�p���UŨ0�b7Uh�{���%�L��n(��zh��N���y5��L��Y�ރ��t��g�,��dGʓZ;����:���0�F6�d�!zDwzUTd��3��}V�H��uJ��hYt�b���ո?��O�;�u�rR�EH������9~vog��U^Z�Ғ|���e�/���1]&���i�_��%/�ڔd܇��f��<>N6�#��2����a�G n�D�s�uB��>���G���q�ބ�I[�?3,�������C-��>�3Y��io2ϰk+�B5��Jrj3v��R-'/���E��dC������oz����/	H�o̥�fr�-�j$���v"�R&+fꃈ$��-h�j���b��
s�BaV����������w��6�']\Zf*��� �\�)a��~��Z�O�X\;R��p�X��-��D���?�Y�+�"�=x���(_���	;
RyI�K��[L������������Obo��j��!+����*��1�L3V��rv�5���ʄ��B�_Ą2��*�Z���T� �-BT�	�8�%���4Y/'=;pi����B�#I���c��ڊ:c�Ζ�4�EQ:��w�*!�Eq�B&���H+_n��Ð����y�D�[���{��2�B<���`�=�.�O�GZ
	D~6����,�:@ߙώ�t�.h ��9;��)d����)�BTz�W�&\����]��y��	�R'�k������;8J�g���]VM,Y��	�͹J�@���9�{�����}�|~��K�{'@��Dh�UKMZ�~DUC���V��������z��[�ݠF�w�����U9Y���G�H׸B�4�XI��tm>�@�bq���BDsߑ��1z,�ӕ<{E��p�G��ev&5�7P�����I
T&q���"T�V�%�,,8��ꮣ��������+�Й}���mtv����[��ǜ%ƚy\u��p:���	,O��Q�����U5q���Y�Bܨ�Ž+V�ӳ�ʏ.�8�ږ��*��� �A4>�`κGX�̛7/T��P��[y�X��R�L�TP��s�	K��KaR��	Y3g��`_.��Zb�D���Z�S��ꨒR��������1�8�I�m~�3�j��=�V�9y¨�.����8N�+������@�hr6v+S�K�Z9�t��SŅ�|�4@��l�{l�W>Rr��P�~���&[f�o���j�=�~�L�d�Q��/V�=������v��r�e��0 �&3+k,������%��F�6M-�Z ��0�ota�W�|m����" �ĢءJ렚ٛ���t˾�A���&��y��*�`/=�ֱܯ���Ջ���׊H�l<�\/�YL00�d�ф�+�lo�oQ�
�u<��d�@Zf�-j�F]5����#�������h�v���
-�+;�Cc;#29h�[�n��݌�5#И�b��r����,0qr�������#�uPP(���a���F��y�0g@<�P�FT�=�b��� �k�$bł4�����TXQF�1#��� _,�-�]��I���E���V��N�:�T[9Xυ�J{�c�6ﲍK��Vj�7S�D_����49/�)g��Z{6k�B|�`���zP�=�1w�p��Ͳx[���So��s�53�ß��̣R75C�:(��! �⺪�t&�z����r�<Y�!?��YJ�P�$"�ƀTY
w�����䬭l0y�|��ni��je~��7�!&��\���a�,�ʺ�*H_i�_>O�z� �,�-��%�G�9yTK�Y}R��䕺'J�/�O?���̬(�^ܘаB��������Zg�)KE��l x)Z��Zo	-H)�@�~\	�M��F����ϕ<F�/yN��",��`�Q�m��I�=�f�%���ă쓧u��Tx����0��{��V�K���
�'��ܡ�� ����\��l����E�p�b��2��k��=���*Z�N�T����a$_A$��}�oad����=,'���!%�� d�҄��"��1���3�� 2�p*�Koeί���4�[��b�&VPr�����u�0��`E���C��ߏZ�vꬿ�������SBBܫR�lT�V�,�V�ٹL��
(�wN�#��,֐����B^�D_���4��p4V�q,S>�!L�{YҋT;@�(d@��
ȝW qR�]�;3����>�e%3-'	�=�����O�@���'�x�,���Y��I�j��߿�b����OWJ�Arz����j�K���nIW��Y�֞��H����9e(g�˗�l�WNֲ�>(���~T+�ɓ=�8ِ���Ma�)1�j��'���YX�E���jUӢ������i�����E��۷�0}����fX-�G�"=ƪ��ԪF
�M�.�5CZ�+�iu��;�Z�"HE�$�!�@%��Qh� }\��*�,YW��}"��X�tDa� � +M�Cg�I�Ғ|7F���+l��	V����
G��<��'�b�,���	�b�7�<ҫ2��}1����xNƮ�� 觰�̼�?zW�մ�;K���!�yr�;�a�P��bg�l���L`} ��Z��g/	�5*1n���,�]b�������$� Hz�G�ĬSnb��gX����Bm���Ls2�^���</����Z^Y�f�t@@{[������vU�Cb��.Td?#(L��j��yLP]�eh�8i��Z(�{Pk���}��$]o�K���7� {��8�O#CpL�Y"��"�#��m��Q��8�I+�}��tj�p�O������Ζ�V�p8���'�*Y��� ����4kN��=���%�U�rL��F��9|ڷ�%�c	����``���_�E��ב���3[�<��m-F�Ԡ��a��i<�Eݫ������v�	$�Da@j��#� Q0�	h� 3����/�0�Ue����P���y�����5�^'���Ei�RN�����T?�3찎��Aޤ̫x�浡>�L����hY|�`�,��	,�e�;K޶��q|S���V'�0���d����'���YĲ�Tϯ{�!{��wu�aE�r#Hj�J�AY�xv�ʼ�ⶵ�Dn2x� ų��R5�����v>��I��C���T�*d^�p'$0Sfo#ǳ��cL�*s�IY�'�5`aU�>6"/mK�5k�K�gf�\p�O`���2Q�q�y��Y��|B\m�Z��R�/�b�3�7fuSU�[���2�2nc7yFLʨ���?�5E��(����i�
�VWQ�b�C���^�ҽ[4�cƕ��.�:G��R �[�B�M�Ig#�xB����=����Ě����O��8Ҋ;v��B*��u=�TY�ü��<��K��#s%����=<�X}B5#���@h�X������ƦwTD{��4��̯̏(�Br���}����i�H/&�� #�Z�׍		��e�o?[���?���?�����{��aU�& wч��:;�g(��mL�і�=ښ����Y��#���Iy�hunULmI`��� ,�:��b�
D"m����u�v�<�=��F�\�
�����޹��/>��(���YX�p	�c�1|)��m�M[2�m��sYae��Hr�����w�)��&H��d*�I6����w��.��{R!	�������r �-��7��_-hV�ui�-a�
IDb�.�nr ����2��8�7�{��в��wr��A>[�3�~���K����JY,�LK2��g'�s1����h�n`�J|�]�41j��$)/�*QXr`�M=���*�����zP���,y���@nTÈZ�+�Ti���Y�����*Y�>8�R�$$�˅>�8�~���Y.w�{S�6O:�fn֤�Lw��%`S���,�����5L�����>��?�L����ɞ��`�4��T+��	�C�%������k�����_�����r��.������V!+�+灠R�A%H��l�qk2�ZMBjP2�xn��kѳ]9|Eɼ~���L���:�d8č��MdV�	�u��~���F���,��!�$>%�5Y{Ih���ū�k���s�������-�����E/}��QRN"v1Dd��^?G�Os|��ެU���O	�1xٌ�ς�7�Fzݵ6W�*H7@��Ҋ�+E�7��e���Ԁm<8#Q�[�	-Ж���ߔ:�T�8 �vk<�2�ĉQKE����'h
FuG�8���~���\R��Z)���:�@j������-���@�>, ���u��p�(�3���H�4�����B��~>c��Gk�_��J޲d��K
 ̥	���3�l�!2�����Tb�POS���;Kܦf�W�Z�J��R]�f�ǌw�K1������Dc8�rn�sT&�ׂ:�����'��L�O_��R�:@�@[�ir{X^śj��sb�O;*_�~��$��&�Z�l����4C<��'������\�6��6�v.Ժ;F��%��)��`�C4��U�]��uO���/�?T�QJh��.��0�]0?-��Hq���f/n�������� �	�/~�Dd����5Tv�C�Q	U�+	uXTB!�c��]�*�$}�T�<���m� t��f�	�2 M�,v�,�ͬ�Z`�^	⎃7�B�$�_�l,Y kdqX����)�sAO��l�=��O`��R_�$2CD;-���Gj�e#Y<l�k%�|V�ǳe����+���	�m�������B#T�ЂXH�Y�G�:����T3di�v��N��\�ܯp�� �=����~��!!J\Q����	K^��������	������'�s��|��0�*��߁��	i�十��%�� �HƪɅ�fzJ�i��?x�19������ot>>��F���^���	�,*5|%Ș��tv<�6j\����V�8cYzP/@�6��0�����'3\����YY�X�j=�s��A�70�{��L�f��gI�Y��6��e,D�����Q�B��:%z/��x��hB��9�b��#�<�Y4�b�k�(!��|��z��.Y��>�:6��"��qc��%-$b2.�L+Ӻ"�9ۂ2&$�'tm���?���,�n�k���y�E"e���AFh���ZcM"<?)�K���Q;�/����`��̢�H�;�0+%k8$�����h�T��[two��n"����O}�w��S U"|<����/�.��U�BT��|SǷ4_
*E7��h�_�i����1�f-'���<���b�/c��a�Y�V[� ^�ĉo?H��$xW�&\Ɋ��%���Vw�|�4o��V�gз�k���6�%�Oel�dԟ~jk����_vȎpI-̰��.��`@*0�`)����nҘ���#PR�*��3�ǲ��5	N���ʆ� ���d�B�UΌ�Gl��]q�*�o��O��s+r�Xt�g�E��B�,�d�d��:�]<�PJW��'~Y��R
�{�3�;W���A&�<����Q7.���2�����i�El��ؼT�tD��ܦr)�1d���pݙPe>��£���Vv�^f�ס�����	�at8�U	X��y�k�rK�ļ��-������TC���w��bN��8��h�=bb" Ξ�4��)#;&&�����CJ���_�V޼7*5��5�� ����t�g8��^�
�Q�<�1�fQr�:$�Xt#[PT�p��<�G0؛er���-TH�0��n*�����n{?htS4�PͲ�q��?�O^�Ę%�I���V2N�3#oE	��Q�(�Gt��"�0�{����!]3K��"��y6�x�������~��s�b��z���X�ۃ2~U��3Q���c���؅Ejkw�J&�/"�IS";��Q�`�[���U@�:�+lƨ��ep�ek�9�f����jz�ʂB���l���H��ݒ���Mv���+i���]V�T�d��W.Ku�;�k�0�"5A����i��,�_�%�x
�8a� #��s�~Ql+��
���0����"9�"��I�y�t����a�{�D�ڣ!�ջ��u��K�J�En9����K�2����!�晾R��g�ɉ�#As2ws���G ���Ѧ�V?J1��oTK� h����Ы��H,�w��s�AeJP��5tPGY�J�Ȩ����rZ�Pn��-Qc*���n@%�>]�X6�^�&��HΜ��B5�O�q/և� ��~��X��{���%%�;����(� ga�%xX3��?��0��G(���Ǆ���n��دG���f�XU�q��9�*�h�F&-��Y��c�]����̏�d��X��FR�	q�\٦�؋D�|2��u%/��q�&�)��&�d��I>�X�ռ�[/B�	#+ ֻM�.u8��*s�Ks\%ٛ̽�s���ѽ�x(*�����b�}s�nq����a��rGh%�	��HV_,�^^s�3�W�Ԁ��f�𴴕�]1,j�4:π�=���H����A1��@����wr�&���z��>h�ݽ!T��hH´$�1�sri�V��Jez@B���<P����o���3覑��/���b�2��n
�^��xĦ�/f]_ί��Մ��#�XX8L?��o����ަ%.�nX82&[}sZpY����(0"�Ț��)h����V�q�֬|��C ��D,K:�T�o��]f�XQ��)^Ԫ�ȶ.Q�Y2���Q�-���us[���:/��{���R�) �6��[ēiQU���./��ƣ�qߢwc��}qq��N	�_ {^fk;R�
�;��	���ppK��<��t�>�2���݋�η��d�I�v�U���Q!����x����$��L��=c��X�u���*a��O��MY�PuD�zf�Y����݁�������Tt�QK��n��pH�(�_�zR�c�Ϸ�(o5д��\/g썶=�ƒrv�rxBo-�[����N�<��~Y��5))�����'�=0��ރB�����I�D�0�~/ D������e��N�+x�dmIkB4�F�s�k�~�g���{���6���5�@5	-P��h�e��E�7�̜��X*ndҵtV�u�|W~Y��L����J[�9��[ڌ�{�0Fς�ӎ�(,L@A���Eq�倸c;z�`KR��u�m���&5�ӣ�)���o}C�yH�X�B|��a�,!.�x�՛����^�������>��G�Ӓ���?�����J�L�Z�J�;lljd9x�b���7t���Tw\�3O�@E�[;�OWwZ�i�� BF�(�%��Z(h�lɪ�;�j,h���3/�R0���&L&+�e����#�_�.H�2\�/��$l�쫯��À=o�����A���{u)պ/�5|�u4;J�S�Y�L��9c��="/�e-��ZC�{�ҠK��#`�чޚ�ɗ�#nQ�eBX�*V��s���,ހ��Q��p�F����w�6e��`1��#>�24"�^0L�<��ܵ�>DX�����N{�YL$�w@�<�6R��()�.����}$�l�d���ߕ,�,i�3�H�O�"���^�Ze�n��T��tBك��� �HA�l�b]����$A&@��I� ��KҊ��F�p��ks;��Ć���A7!S|s��*�H�`n$N"p�Z=p�p �E�m"F�D6�d#��>M0ka�
!X$҃PL���Q���V�s�
���T<�B����B������u��
����ߛ�#�M�x"`b�[�l��|-��Z��Nk�͵�����0K�m����/é�B�x���7f�����S(��6�Ξ��݁��%�{��;�{��>���J��R%Hx�\��B$x�9{6�S��������~V5�,8ם�*�;C�6����Ř��"Q:{�	�/-h⻙@��~ډA[�<X>�@x�۝{g�V�����}G�6��k��9�;m����v���3�P�s&Z�a�h�nR�����e���U�P��=DxĔId֥��g�|�;7?ڮ��!2�-
�J�&�9�ɠ 5�^�*d#p!�Y�uT�2->A/�MPA�Y����
�D��b����~7k=�Z��߾��K��%q�.�N���ɿ�WȑXdgQ0Э1��Z�w��Z jѭ�P���=?w�ś�'��VC<X��U/��%�#����|x���r��
5٬2/��ن�H��a� 2�Jx��� B�gi8&ց�1�*��bm��X-�#*�e%Ze��pԄ��,/%
�FxaB���gp���`�:����,�/
��Y;��!
�n����KWe���uʹX`�s�11�J�	g��hئ^�7���Jf0��֬�q� ��1���o4d4N�̤��R���Y(�Z᪒�%��ueB�!�?W��D�S���>R� ����X�e���+k��!�@o�֘�J�E����[\Y�42�3�ع w2ժ*a;E�!/
��d��PK$��uc��V��g��]��zx͠�[�\��8s6�GFB�hWK��2� �!Ft*V��4*.+/C�-YM8��C&��b��:��|VX^��f�t�m#���c�a�~_�q%�75CvP+��<�`"�Q6��* >>x�D&S�c$��z���5�b�ˢ)�=��XC<�[v��
&!uw�I���8ʃk�YI��3�.����+�H�M1)��/�(���Y4��ޟd�ZW���؈��m�ЋIY,LPB�Ï?�@�a���ʦ�X1yB^���X�ujfS:;(J���Ϻ1Ņ��RF��:B&yn�	U��x$�r�$q�?@I�|� d&�ӳ�^�5}�̲|'�XP֗)\q��Fd�e�h��:+~M�ݼI�X�;!��&yi��f�JI���?"�y��8۳F�����v�� ��H GA�%����gX�zn�������L�3���Q��Έ�����ep���Ef��`)c~B�U����(��i.HY�nݰ���\
s�����[����W3�c��&o'KYI�Y�&�ѱԕIS7h�f���D����#b�̑h���qP?�KI�T�!9^ٞ�rk�'��(]5Y�4g�]������j��k �5�tY�L����ĳ�`ƀm����RR'=eԊ��������W_~��̤��������/��(]��j������L�Ӄ�׿�M�.�=�tvS������$��V�b���1��b>\���,�2��ɘ����
������Y"tۊ��h3d��[�ʸnJ@�u�S������ʿ��O�?��/�T!q>A��S(� �Y�պ,�����^2G{�CZ|�	�`�;-��Ib��W�N񒂘�$k�����-R�'�T��B2�q��{k8�X�倾�KRaK`�r�y^]�]�nqxi5�ݯ�v�V�|�"�����g����|�ͭ	Pُ����ٱm�ģe\Qef �\�wo�`���F�#k:!�&n�4���x\��L�����c�n��Yc��Q=��l��r��۷V�W���Y���'?�T�'X��l�H~ =���P�|T�閛�rB��5<d�ŋOTl< ��1��˺���k ϳP���V��s/2_�'SjR��ȭR}D�7�u���:T�SJ�%����$H��-ʈ���y��2KC�eA��L�Q=Cn�l�$XŐŕFџ�M�͝������Z{�ŗ_@�[�P2��5�:��b� wИ�!O �%��1H���/�P��.`�HR�y�]�ip��6zɬ���n�7Գ�V6!���*Dr�A[�5�;�99�Y#��X�>�^��>�����:/_�%B��=(�2�L��/���)�D��:ˬ���(�kl98_fbb�-ɀ��M��T��|B[B,V;�ʜHi�h�<f��8��v��i�Ͼ�[�@��2a��C�ϻV~�|���$���A��/�|�o� T���;g&;�;:��Ԭ�s��Y'W���d��6a���M���`��{�:Y�܃0<9�3�?����=��?Q<�|�}E�턎�X��H��lu������p͊Qp�_`0��k�[mgJN��ϫ�)��P,�=VG4�����{nb�<��<�X�����v83��G��#k5��������ɧ^��D:ˣ/�q�P$����d;b��,h�¸O�������fF�ENH9Ϭ�%�:.+P���)��j9�#n��4ެB���Q7����]`)b7k�`:7f-k��BP�U���C�P�^7���i�#dn���CӮ�̍H ��W����X��v&I�.v��4�̹2� ��J��^5%%�o�ӯ������Z�(P'�7Y���MM�(�@VQc����O 濽A;�Ul�Eߧ�{�>��+,�q�)���f��&E����{�[�MJ���H3���+��z=����]�^������+3�k��M���5����bu	W.TB|���A��13�Vf<˂˿٘P1�ɝg,p������p�^��ɕ��%V����L�	����4P~���5B�=�j��PX��lց��+�ȹ���e��
�a�]f���XJ�|c�'{��r\�Pv�J�S�O�2�|�
e�K.J�����K��p�Vi�28���*H���"����K�s]J_ɇA���V�uN��x)6E#$�?���Ad ��]�X���q�e��ز���1��V��*n�T~�5���X]��U�I㹗�����k��u)�1�ԤҒ�N	�w�)~T;2Ni�F���{��_b7hLL��6{\S�y�9\��8���?��������V��<����7��'맘?D�o��)���������o:G����Z��NNj�hx��H�w;�CM{�rI{��3�+��h.�o5+y ?�HA�����@�cW��u�1>��T��l
㔌C���}��^���߮n��k���ȟ�^а�szx2rn�ɲ�b�ҢȢ֬R�I(B���^��XV-�F�^�ú�>i�I��|#b~�g�]cB��ʿU��X���²�`��݄ɽ��XF�o4_�~R�	0�UxJ�JHX�u~BՓ�{Բ�������i!{R�u����;;J��3BK
�q�Ӯg��@���,K��w֕W�{��u��h�x���d_
��
A�h.@8���|�'$��h᪌o��"�وW4�2Vv�e�����l|2⤔��aXs:m���	�H�&a�L�V�ŉR�����j�+>�F��>/�;ь�6w�%EZ�h|���A�`%k,qeVRƧ5��8e�������a�M��1����|$�5�}���F���`~XF+��)-ԮƤ�Zm[��٨���
���Z�e0��-���Y[r؍hמI	DX�� �9�UG̈u��gnƦYcp�@{����l��Ү��b��0/%�X,ƽ�5�"IC@��'*�Bv�@��u��H��mHƴ���|6-�X��2�X����-����Ck�΃���(��=��흹+�6�v�i�a�'�K�C���9�T�TN	|nM�3��H�w#��G������x�u�P,S���@'�cU��aT!)�f�OfE8�F�W(��s�=C�rR�����=E��90(Yk���>w�Y�hPˌca 2J���v��ن��Ͻ�	�hx�����i�`+�>���/>)�[�Wu��.������N�dec�Ĉ�! �
a)v�h5�(�=��S�Y��4���������Q��e|�);���/�d��D���]�B�gްYd�|�bR�8Fu%�;�� ��(0�/��F��M�q�G�G�M�����H�����"dw�=�=Íň�p���a< (oqM�-���.��j�g�S/�&����x*�=�ɗ�!@�� �!_�%��\-Huɠa�k�jX������B{��
�bG�\oΙ@ԇvŚ��̩�R��
�|��<G��x����&�Ș��ڼ�L~��k����; �5�	��;�����َΈRlbJ�b�A�4˜[`p.��p�+��S�����f�E����-�蕊�[-k���n��|�ֻ�b���rU�B���`���npV�M2�J�qL^�T�l�L&4�q���ͭ���kr��n
��-DC�!
&�),)�2�#�����O�9�V]\����&$S�L�X7R	"�d�z+H���s�V�~�ړ~o�]\�6��apl2g����O� ̪�����b7�X�V��Dٛ|)�e�E��*
��:�{Vc�`�v����:�z���&��]%��6eqx�'-�nn��G��������������cJ�.{c�gu��m�pб<M�W��M�����a͚r⊩ U0j\K�Ssw�ղ��?dϕ�\�Z�D`�ߧ�OP�nJ�3�%�*G4�[p�>��m� 6���R�p��AF�9���� -�����(��-d�'�Rn�krAK��.��m-���k�k�d�y;��b2w�3R�l�*q�iVAO�AA+��K<=	�#�h��"��;��E�F��Y���4
�_V򢰅���Ln�OaDb��^1�BMa�(2k?C�	�����h4��"P�����w;XG�@/��P��}�yfAJ+�?�Ӑ:6�r�b�K�7����� hAZݞ���\U�#�L��A3>+�$vz T�,3,�܊��lu`i(��}�Vc{F�yA���R�=�z��V*�B�z/�w}��F�4]�	��R��E�����_��#���Wak[��J\42�'lOM+w�~��J�I8��*�3����T��dr��2�K�at�dg5��0�����WR��z1��
Kĭ� �f\O��,��l��ϣ����?�l{8)Y�D��Β�dvz��@"G[A#���-^�3G�UM&�M�1�"���3i��؇u,����jB��T\�Y���u?5';'֓�������1�.�2֛��9I�e�
q��M� ��yr��B4Z.۹d�s�ZIǎ��� `\����F����3B;3�6GY�� �2Έ���8K�	60$��G��G����ix��IJ*-���$0a�ig��û8���2�u�[a��lxI
bR���x�j�ea"�Y�(����)���pH�>���� ������j�*�d�n�zD��Es<=X�e���0�97Mm\�����6!kD��3���T�
�|E
��:w���+��� �̩\�P��.!Lf�D�ԟc�zpi�����,lP��ն+;w�8h��i�]����`O��Il3z��%�4�+8�ꦡ��Yc�6�m.�j�*�uk��3ѨE�޲Ҽ���5��8�}�QgG�O�b� vw;�#A'�X��?/5N�A�ȏ�/��6����b����5.�+</�+��п�~�Z��h��]W�H)��+��Y!�<�d��2g�� �l-ޘݨ	,��K2Y�/�8%
<kOm���hk�*d9�)�#�RJF���p���z.�%5�R�L���f�F0�O>�T0!8���S#��V�e-�� �!�l�2��}��'�q�53�A{�Da����$��d����s��(�/`ot{��Xˑ��xU�,�Z�'�,��D�''���G�8�]���#�꤄�L {�Lo���v ���;+f&%�@L�2몙M�adeiʨh�!,�
x�w[\~��2�O@�"�ǧ�j#|6+��|���9e�A�\��b�wt��h&�D�#-V*�n������ŐH:�D�8[Hh4H��|v�e�kل*�[�ė�mA�)��Q��!*�ܵ���N��gzH����g��.=�ù�\�=*�&E������,Hgߗq����*������{2�c�/���;�؆A��N�2<�3����IA*<���G��E�,H8��p�I�X��	�l!������X�ZD�'~c򑷠5M�;�G�W�D�s��%�m%����{�Z� 5��/R��
ϟ4Q�Є�4�:?��['YkA
�%����͑Z��8�D(53�̒3I���(�f��jGs���BMۍ��� �b2Q�u����>x�|T.�p{��d�hѼ7�E+�<
����U�����gW6&����ǋ
�B ���պ��vv�f�I,�k�ĄEa�m7�#���-�����D���3���q��vc��AK�k]J(��Z��J:+�0א���Ikb������K�ٳ�(��/m9���uM�z��Ƀ�!_�gX��V��a̝3��?�!��et+D����=w|͡��1�Ӫ�j����H�>	Z/1#Db��iK��\h�D���r�LF�I�m��-��[+܀VΖ�����{<!F:$4�52<���݃�l�x�c�]k�&
���f;'p��S�)F,H��� Z��(]��ap@���!��-�Z��+��Al�@�7�%�6�`[��!��%�Yנ�g�b��*�:�o�`4<���Ye揙����$��4i���R��pB�b�
B�YZZ����	��jь�bt��B{#�C�������#�L>ǜ��Pc��Y/&�'$:HPc���x�!AN����u�Y��?�bY�%�W((hMRIx�
��05k8�l�@��߶\&/��T����.pS����"��P^���y��:��p8y'Z�k荒Q;z���{_�������Y2�Q!�[�5A�ѣ���.&l��ͳ�빓� k����M�z�i�l����`��~��5��b(�:�6!��F}�s#��#�?<��x�-qyэ�%ҚTeo�d�1ob�O��2b�����1}����/��/�/�������?�q�%����Ҝ�����`���"%��ڣ��8����Ԫ��C�ԯ.�6�jmM�x��]G`��v-�j�6�ט���#K*�0��\59�)��4f
E-��i�&�^�&@)�(���s����y�gGV���U��1�΋�-	��B�P7=CZ;Ʒ��!���e&���`a�h���n�������>R�{H�Z���n{�.XTqH͵���MFG�bm�;a�:ަ���d�	�.|��ܽV�����z"�##�l$|6�Ґ�ɞ$�sVg=d�b���U�%.�v1
�7��bVii��f�<����sT�Q�f�Ʌ���~����W�G)�%���oj`���u6�4�7�XlE1����|�����GŘ6�����5D�i������M���	3�T����+qϿ����e�-��ߴ$Q(Ȟ�M.6)O-�xV��'ب?`q8�f���n?��9"Nf���%7�-ښv�����R�u���-l�/܂�poL0�e�n���t ��_�\[��O�⬚t���"!B!���P�DC(�f%!�V����9�=y�Ň�2�[�OK��z����Z���(p�������R��7X�YM�hk��S�B!sֺx+&�x�}�R�?�� �h��&�U�3�Ë�x�Y��tA������g*��)S�����ka�4����`��Vl���[�q#@=��� υ�l��gB�-ƭ��E���B�*�k B����n���D��K�4��8G� l�Ҥ4��Έ�z{p��,�s(D�o�[��A�4���
�mH�����S��5���j�Jl����QZ	����������)}��	X^^d�і�s��W#�˪��pA3�	c����ƴp(0;׋^"p.�D�Iv��t����P6�M7a/�K7Y�C䥿�� �[]�^M�������h�%ǋ¤���/i�y�
C�����BEh7\����ܨ��5��h��ka腡fԏs��K*j&�5�c�\��'���ҽ�<>� L��a�H
S�JE,s�T4H3�Q#:�����'�d�<Ȱ��$iaR x|��1N*9�NJ(osvrl�0�I����;����߆?�kL2lB!��łZ8��>"��j4B��$	����]H�E�\���d�u8��/�a�DW�a8P��^U�HuN�E��e4�İB�G�D_��U^��/����"�C�Di��7��m����,ز ���������Qa�8^q�il��W���]�KƋ�TgP�g.ġ���+]�E�����E��G:+�Rh���F0o�뉣+
�� �x����������BL+.�����������j	��wZ��
o�����zR��K�"ׂC���w�[8�����Au_C\^���Y��H��p�	h��M����mU��}�"ͅ��9����� �6�S�2f���g>7�е�� �Qa	$�GuIC齿��_�65�����<o��3B]����<Z�˳�zM9���䜼��^,²n�&�S
'[��A�-��u��M�vmDW͡<����$M�WL���]{��v����55���"P�A���pp�āV�c(���b���@�q�ԝ���͵qLTS?'Q�����ʵ!]����ڞ�ϼ�<�|��5z���&r���{C:0�����t���a��°� ��j���L���*"�=���mT�Đk�����_/���}w{���e,�n��h���:b-��-:Go��\��xN���Fk�kT�FW�3y���e)1������Z6cʹ'�9��M�J53�\YNjw}f�*��5`�[W�p,~r���औ���VpvV��o~G�����k{��['u�#�3�"F����� A�?����,�(L����m�ľ��I��LK )�I�;]��e΃��_���o�����7���0����$z{*�M�D|�po�˻�j ��F�лu��~�������^�r�V�P�����Y������!�������G����E���h*�qAZ	=Bɥx�"u��Cd\6)���M���:�k�C<��{�ֱ�}�ѯ)��TP:�C�U��%<�8C&��IǓ%� �)2�f���iaqt����
��l'D���*P/H�@|On}2,���n��ˤ���W^����U\wZ�����ji��a'�,y��͡OkB���~�ן�J�R�l��p���u�1ǪS&)t�ަ�јy\�$�b�9�^���g|iKR$��P�"ݷ���d�;��o��V]i�_�\����r��fp�
d���#�:o� z��
FU\K�+��JRD����^.#Ӟ�*�n?����O�Y
�\����{^S�l`wE�	��zb&(�|�������b�"�&�-�0d��Pf�$���Y7�[Ʉo�q����f�?g!���	���`!<+��exV��u)i3$I}խw+�����{ŚY����Ą��F|-7�	�-m�9��,08�W��vG�u;C�e���ee�wo���k�?y�� �T�ҽ����a��
k��ΊϞGKmB)�E�-��O ���<���o�}8۝!�>#?K���(�;Oo���z�� �g���	F{�q�8��n��z�M�u~\zCC�b�i�u_ ��\_;��"l������2�}��% ڹ�c� �3��V�0�(��Yr�Gx�G� �%�n��$�P���W3��=W�E��� ̖B�����Z|����ul+��#*�w9�85��i�n%=+H[w��?Y�n:?�BT���p���c��q�YP�|r�㙻���0/����6���愡���n��k�[�Ʈ��
�Y���������]���Bp�{W����#�E���<g�!A��I�V���f5�;�h�Z�=���%�P�.+2f�ՓJ��m��n�!P-m�4�U���wo���7�J���{��䁻2n y*�&���k#�~�U:�F���V)�(KT�X%�M�}�6��#�@��(��ý��{1���L;�4	Y���n��K����Իn�������=��q��(ka�tx����o$�[Z�e�K~�Ί+�~![��}��#&i�e����Xi�����-��<���Q���F |�{*�th�ƹ+�����7[+�&w7)�k���[��8�# ļ���F��ϰ�d�1��_n!�u�`=��&Ɓq�ｵI�C��M�����}�Br�i}����s����"aI�_�<��A�Y�n�XN��m����PX��`hK�0kz�v!7��5��]����]���Ш����6��@��ȉ(c4ɣvw��R�.p�Hs nH�<km���jz>_0
Q�3Iݜ|��S�!�Zߵ��%ָ�[Q�}%[�I�*�t���z�C�L��m�	#į�qRu��%�$	0fηI���~1X#��6����cw�@	K�>�Pά[��8JaX�ST��/e�����""`��17sۖ���Os�U؛���8H���x���5���[B9��֩uQA�=#=�O����τ�6��=��E�dM��"?��VJ���S�?a�]����S�
�{�r�[\ؽ�����-���%�a��n�(�)�bѼ�P%Ƭ���m�r��e�[g v�}p�:S(o,���[�|���TZ1-��t3���eK._h�^�V��*绤�8�K���߿u�ʏ�ٸ�	�Ą_�/J����,��O���F�iK���ª)�[KDh����,&6��|v<��I԰�<�g;[Q��Ԓ��[I �bU�����u�(�+��oXLi_z��a����h��}������JV[Δ�}͐���J"%IJ���!�yj<Zu�&[�4��^<�<�`L��q7ɽ��'��y�>�S�Ҧ��8%Y�Ș���9TNK�}�6QP�y��Ԓ��	������ٜ�Eʉ(%V%=@~%�l'b~��Á��bf����7[�=�$���!Y����S�|�3+�kWX�y ^ؼ:˙�[�@��C����^� ����:��"�_1|@���}ٝ�ˇ�-R$4p�D�u�cx��T�	*)G���=殭�ln��N
��#yF���������=���������S;u+�a�t���1�e�?��.l[2*Z���g����a8��K֥�k[��E"A�V�R��wI�v���מ�?F>(��+V�!����+�钖�7|��R��
�Y�N Ş�O���5<�~�f�%1�_tw��Bcm��?�nO�^��Atޯ���x���>]�a�,����B�٦,\�k��8]']�nB�6��V�w�bz.҅�9�6�-n}S��aUl�� ���y"í����?'��"�ԆVNZ��v�1�!���'��Ei��FK_~�4��B4�-d�f��[�Y��s�c�v{���SR����ׯiX�����b+Lu���^���B����<j��z+��_�kӴ�au4�t��Z���g�S5�h�j��$�`@ޘ��/q������B��"��-]�Y���O�vV��պ�Z�r�jٔ�f��%�uV1�!oȬ��X�^r9����v\!����O�����rfrc��E[��v��n�������X�k����twsś,�3YM:�3\�\Vm�tqQ�܃cI��\�4(�K��X?>��m�D
��|~��X�$Q�G�ĵ�v.�W�Q�aV�PH����y,�_�D+=)u[GVp���\;s���1P�w�PW*�0�J兩����;�i�H�Uu�8�qi'���&Bi��ȃUR��8��LI��d�1$�~��Ы��<,f���)9��C�O���l�h��V��w�����R���5��p�ݚ��fhy�b����`�)��S��lx�A�K�C��h�{Av�����/�ä���w*�du������-	(ZE)��Y��~�qZ^<������6�@ݘ��ܧuǓ�r��_�=�!�脸o~]��h��w*��F��6�qʘ�s�Dh��fܤ.����;�|=�|qo`�0)h-���K��LI�۹��5����)����S��u´��u�qEjr���td��K�6�y�R��Ya$��kSh������o��#������կNBw����3N�gW�����!�qmV��8��U'm��SJ�t��@�M�qA:�c$�'�E�Ԫ�'�$B:�-٦פ��/-S^ޯM��UhӺ�+�!ֱ?9���~��`�'�����r��N�qi����͊y0\��*��?S�4a���t?Gۧ��	RdZ�ɂLe��pBh��+.?hf���A����;�(0�4B�ҿ��cU���|{Jr��ݔ>e�<�R�'j�=�\(�)�)�f�m��jnEWO
Ty�`M�K���&���l͛ݙ3����?V/��f�NA��ʳ?�rvk��W ����p�@�,\��[P6ٞt�8PZ�<��[<�Y�w
��5�Y�!԰��T8Q�otK�o�=]"���-�޾��пek<�X����-���ow%C�sI�PI�%K�VV2�x��!���Y�u�.���4(�m���_->���|�=��Ŗ�B4�Ҟ�V�u�ֲ���I��H�z9��ݷ��l��Y=�E�� ���/-n�g�c�����ڸ�u�x��Z��w^�k1�xM�n�����~�N�EK�ژ�4���}���ܧ��\�(!D)H��u���2�����u����Iy�������2����5&�F��I~MB���[z�J�	V4[?D9���qP�K����u���kSS/>��(!{L��(M�J��3�sZ�nusZL8l��U�����a���"5��� w���'�\����qa��Ǫq��İ>1#��I�m{w�����CQ��7���I�n_&�m�<��pqm��vi�a�Cދy��l�$v%T������ۥRF�Yq��˽�<�e���U��NqУO<��3��[��D�*(���t�vm����u��ͬ�|�� wQ�Cw��p�M�pZɋ',�����:����Rx�\��sa�Z�E���+��e!�E���smQg��Ù�M��r�/j���b��	���A�ܒ�$�/[,mޥ��g��O�H��,S��"�����E�J$���,{�j��5�9�DFE�"��ܵo�l^T|�����%%[m/DC��c07�ZaI�R2�2B`�����L>6>;溃m�٦c�L�ﳡ0�S�������\,��j���i����I`�DKqX�������z;Dꎉ7�bF��n�-%<n����;���c2���e�!-������N���u�?�W^���;~Q�O��ȷ�����c���,�z�=�ikN���:K"[ afY,���A�qE$Tx�)ȓl����r9�ܷ���}��ձ$�b�f��k�7N`�q;�<a�,���K=r��;��K���++y\<\�����i��|mEN�)>���~ug����}�B�_���k	�Z�1�lV���k�0�||�n	���!I`Z���gi�2]�[��pkj�xfH�NM�ckbg��,T��R:>k��6r���I��~���}��ڟ���C?&]�ӅRz��1�X9��38[v�N��\�h��y�#�J��m�,��ǥ��L��-�<�W�f����]9��w>kkݒTH����,�Ycc�VS�'�5&���b�].:7
��vM�-h*���+yM�^�i��qc��e�Q�ogE��r���>Y�or<�s3c�Q��V��b�箬8,�Du�^��Ỿ��R�ӗџ��I��{�ſE���C}������;})W�������DQ"u%���Ȑ�d�*)tIl��tV�v`�1��	v�K!z�:ޮ�ż���0�v���9��z�R�O���qq.S�T�f�Iıq�X;w�2$@��#FW_aq|���%�����������"m����,/�l�/���[���+�\�Z?�5</((��:�F@��Յ�t�zi�1����`Y�X�pH´nƷ�Ʀ�J�҃��u!ƹn` ��ir��]���q���:���j,Z�1��㷛��jZU���tm���L%K4�-I��:TXyqk��B���Ic��ֹ��0�Y��Ć���p�A}:(;Ko�lg�m�}�N��&�u��u_�X����Ւ5��3˗,�N�]�<������v���j≬}�3�V��~c�C%w���~����i[v��d���0�/w��0�	�,L��	�NX�$H7{�ZLۓ:i�n-Ү��!�^���u1�����__���V�W���4Ǽ��˂8�B� '�(~��%�����E�}m�[o�ør��r8�^�m�)��|����|Y�&��J����
��kI{B�:ۈhr�P
�cI-ea)�bK	�5KEL����r-�Х��Wo�_�o[��IB�2S\p
��j��[q~W*EQ�ll�^�0>3�Eg��Ǳ�
������h����+[&&ٺ�eC���a��s31���o��k���M�����Z��&�j�Lŷ�zX��m:� �����}��6��Xp�I����k���T̽��b/Ș5Q�J��J,e�[��[Ӆg����!>���!9��2��[oT��Uf�E�>ځ3[�I�of�?'���a�9��L�����J������g����k�:1� ���{6��q��\yI�1^r�;L\QfIK�Mփ��65^��ݮ��~x"�����f����zw+���?�彳`��P�za/D�s�s����������!�_�����VO]�G��ʢ�m�P��j�+��H]�B�v���*�!����6��5����^l��i����ic$��^v]���t��\Q���V�@ɦ�%7İ���v[�XZ�8]@�9�GJ�A˓k��](�˳���Y��ޜ�팴M(D�H�Y-�r!L��U�q.�3y�r��a��M����^�	<h��B}���5I�����{�dAJ!�f~����r���B��P��O�����f����6�m��b�C�ܪ`�J����.6$�z��ݿ�m��{�x��т���'g(�7F�6����6?��__�6B�ʥF��S>9և&
�L(�p'�3�_ 䨿/[�����̷d���u+H�)��x�n�%k����Y-��%�&��a��ܤt)DH�+E-e���*n�&�`�:�	>9��D�5V0�D�Ō������N~?��0�s5�\p�D�/&z��ox�Ͻ<��~���O.[%�s�I�/m�p��t���+�l����[����Ȓ��;�8�����ZZ��/�ŵ�ۡ���3�L
p�H
���7Xt�j	\��M�ʍ��Au!J�(���\���.!_C�ۜfM�{�N��R���B�Sم��-ǔ9�[!��$��nt'hZqNLޏV\ý�P{�Y'^������P�;&pMh�a��9W�ׁ�K������3Յv����9�4�y��B0Ϸ�Gz6��?k��<Oc��t��p����A���ds�^&t�T��
�笵2(���/�D7��Ğ�9�'�}�5h������4�k-��59���g���|ie���v#`�5o�w}��R��H^�� �n陂�2u:A	��������/{��¼�ul������][�t#w7d�C����.m�.f�l% ��\���� <����۹�J0Lm-8�ݵ��F��8:���*Y��r�����y�e"b�C�R�_�I� S\�;��3t- `}n��z�����s��P6��gb~��K_W��X%�z����♙�c�_����Tz���.ν�b��m���ykj���6@����q�S}��M@���Ak=��W�aN���8�s���E���k��:�{�:�\��,̻�l�B����ac�O1�R����|?�Q�1�yp}?P1˾� ex�|��b�4������RP��Li̍�F�׌)i/HC����aQhL*L����M��i��?
jZ�҈���$�пG����7�~㤂a*s=�r6��$��k��GO�kL�iO�%�qު:%u�N�Q��T�&�{K&���-�S�z#�
J�^K_=H��/-�x1(�& 0}�L��p��X�9�u*�bB�2���'߭@]||o�bW��/�W�9�fA{�.Zy��k�� R�%!��讏��<�_!X��L�(�f�\���w]g����i��#t�����wm)���7�Y;�0,X�hlX�ǔc����|D�C����ެ�|��]�~^������M��Ú�$���6B�Z��?��F��l�~�*�����1Hդ��b�q�)݈���-j����4{;z��˽��m���,Rlt��"�ԛ���H�J�i�0�p�p����&>�K��<iF԰F���0��w�a��#�:l�j�X3�~�E��q7M�KyN[*ڣa��ɉox��p[bc�U7-*��l<9�#���a]��"�`�iU�8.b09Ⓗw�BR���^�k���7>)�R��:/w� ]g���ѐ�Б�ϫR�8j-	r������}�DV
�iA���	���=� �j�Ε��>-��=t��B+>�\ׂ��i��ZW��т%����<;l~>�]�=��^����%������b�&<0�����P��g0�C�W-Q0b�t8g|�E�'����9�=���ޑϟU	��w���2�U�2�Ie��1=��ߛ���!� �4��f2��Q��b�L���B3��H��dS�����v.���P$X��6�bjrs=c\JG.l+�����@�T7�Xn�P Bi%+�DN��o��IK��،/X�� ZH�T�,���N�����, q��g�5Y�ys�o���b{�G���f=)4�dt�U&nּ5j��<�)3 3�����g(��roʩ���q��Ly�r̹��J�A�����x~U������rx��xx�?��
� �B�;�I
O�cd��{�����l��@��)��֝��!|�J�s��R����y,N�>S���6��(I�3iz�nQ6D '�g��d�*�΄��k��ܢ��9�H�WV�n�|ћ��a����N����-��$*,&"Jb��0���C��j��0�S��$�ݗe��bN�d|�d����~��|pC����Ĥ�6b�ɡ����#�N�IU:��QK�W��)�%*�B���!⳨�ƹ�{�J��a>�Ε;��ٞx��ђ�1�T�q�m�����[i�!�m�dj~0��W��V�rN�>�sţ���[e�9��zc�J�/vó�o�,�.g�k�F���Q�a/ip7sR|�B!�1G5a���YvM�خ�@���اW<�{���
 ���|�!Lq���M�6��p���+�a�u�v?\�����V+y4�FK֫�u������y���n,����is$I�,h�GD�̣���fEFd������ٞ�#�q��=W 
��YU=-��"�p�(
s������R���hǞø���up�^�&Q�f�+y#��а���l1��W�I������@�{���!���Y�x��O��&v�Wl�h���t�3-����FŒI�dz�\�az�p�Ս5��j�j��*��5��h�޲������έ�w�z��E�.<Vz�������7C��rO�Ets���{}�l�Q�t���5^<M����\?_`{�w��_�����r[:.���K��X���6,�&Ԑ�;�Զ��/2oM5���<�ͨ���
=�>����hܣ��m0�j��u\{�`]����P��)8���'��=�
�U����h��T����`�r�u���}����mY�xT���P������M~�d>�rD�v
i�)oO�6�����Qjr�c3%���b�������x��;C��G�e�X[?��'�>[ܛ�j�稗�IXH�̇��k���-	W�s��^fw ��`ה�M�t��+���"��"a��"灇[bY|���I�=��A����8���o].�d���Ȳ��iƷ�T�w�U��U����[���9�y�{�ĿG��Z���o�q��t#eߝVV,�X�r.n�w�%��-�L�?2�����}*}�L�m%���Ɗ�s�Դg�0���l�IR{�m�=Ri��KG�&j��{����3Ȩj�������$_8�������2E����"Ch�N��	��NM�Ƙ���o�N�k՛�	%0ѥ�S��x��I��J�c.�j	�V� �]����Rx�p�k������gb[O�h0>��ǛP�׼ 	_���'�y�Wc8�s�j�)�*���p�z8Fp_Ǐ�"��6a>����^W��C���W0�Ϻ�҄�a��f�L���u��1�����H~����㗚9��nz#��p�<.����4��a����_�r9�y��dcd��ƺ}����H�u3���Ҽ/��dQ�0��
�
`I�hF�!���k�<��g6n���`���:Qa����9��~��x�)`:y�I��}d>��J��wb�;���=1Û��W'0���9iHڦ0��H�R�Vq3LLd�5�[�h;{g����Bǎ����݆�'#'��t�jo��x��N�f4�5]���7�X����P��U#�d�q͎V����J���z�FF���������Ch� �f����ލ��s^,�c;��Z>�yN{�S��mc��ĴZC���C����#��5t�V�(�H"Ft���0O��(����Gnj��θe����U9�y<�'?������a��~�scw�A-��㭅cza�l��Q�=�ŝ'�e��&�cz�;iZ���,_kJ~�-��U'���ϓRH�ǁd{�n;��;[��R�U�8�>�|�v^k�4����u��ۊ�>M������27?%Swm��!*�5	��E����K?A~�����\'~g�����������V�<�G3<pH�_�d])ah(�~dѭj��� ִ�J�����'�<�f`;3���/å�y�`l����-zb���f�O�|pѦо�WSk�M�ළ��ɆԎ �Ӝ1֪�o�y���\�T�c28#"��ݫ�mi��ܰ���C5~���>�a>�k��<�H+���t�3e��Q�i�	��d��
�ǐ���y�@Ư����T���׶j����T��dL����� 
�j��>�86˜�Q{X�^�b�"�z4U� ��K�����N���qW�g�R��ww�+0���kyy=ˀ�ܮ5��;��2�pBj���x*����+����/(��x:V��8�����/2�([	q��yNѲ�m�=�&cYo�p���Y��q�^��&UCf]�8ݝ�����;o��D�-n���Pŋ�����k��R�R5�=Y`��h�݈��߹S��VPQYXaT��ZhW������bE���t�z)w�q�'���{���}ib)�Y�^��I�M�;~l��^�/c��`�D�#0{�`	0�f;�y�H+�i-���F�v�z$�ء�m%A��N�ӂ�8������+9'�����<��Ś7�k�j2�y�Ѡ;c�h�Afw����G:p��b�1�Q��Y�[9�/���7Y�>�� ���C��V_|�v�]��P�f�����,ľw�׭1�䍲e���1)݀صv�8MX�ًI\�z1JТ�{0��N��ha�$7���=P߽�̣,o�j)^J��>r_0��a����� ϯ��i��#è�(h���P��`n��(�x_�x�~͌B6;t�w�Ig�E�+Ƕ���=�\ڗ�������&�TcX� '��6km�[x�o�����0��}y�}1�SZ���8���%ъ��;�����ی�~��z���%:hMG�=�5��_ܰ��D�ƙ��\�<L~/kw���d�~f��ܯ��<�"p�A�;��`�yBRP���3-�<�����|>�o����v��E�ԐN>e11�RJ���>��j��^� ����H���G*���A��d�Rո�ܒ�qf|GU��X��q��}�N�&)m�!��R�E>on�#�@)���f���Is��*=�|�;Ν�H�!�]T!:6��M�573�BV�?�#,�a�E��+���7D���;K7�7�a	o"��z��nz�/o�LM��ae�5�B?>�4Σy�摒�>K��������tާT���~���2��1���.�F�օ�lcU:�?������#8hr8��^.�r�^�7Y�R�m����d��ì	�:{gL$Ҹ�"~�c�(��Z�i���Bb��lD��&����GzΓ%s8�z�~&�+7Ӄ��g���4<�ͽc<��nv��1��@���p+A����nz��HI^71g޽��%rc�Q��/ylQ���?^�]R�~`���4�ؼ����uP�X���Y�-Y�dh�d!����2�֒w�)����1y��a8�[d/���ƞ�9����%R��wx�ك�7�ȳ�q�J󱩴,<He3��4ݓ�WR`����y��Y��&*?����g4��8���Lj��� @7.\��#s�BN��\S�zDX�V�o�2)<X��H���?��J<yJ+��Y}C/�������aWLN�{�Ѓ$�	�p���=�E<�)�@�=Zۛ����Mi����l�� �k-���P��2Y�{�����B�h'/@�ƛ�]�����5�����Ʊ;��o�L�E.o=��PLp���=.r��sՊ��T�--<���z��5G4>��9�98I���7��d��H���pU%���"c�wo:P:1��O�ӜS&C��j��Ox@�9��{
�Ժ$�[�&u�kl�L�Q�J�u��*rĈl��d6ݘ�1��W␠A��ܢH#<��g��z+Xn�b����8/j�K��,���Ui��kڄ�>߀7��:o����o�7s��z��Jr�Vh3�B�K���fQ�x���l޶�������	�P�}K��������c�헭+̹}��߅8u�����[T��[C�F�����.�g(�n��5�nHØ��F�V�7u��`}G��A�8Yt�	�)wS*3uO�C]D[5����ڝ>�~6u,��"'B�6X�`�.�A}�8H�	��ͷ�8���v/�U%q�0��ǘ�'��F���`0 �e�6VH�q�ym���p'̪�����$�3����H�\���%iJd��Qb%�H:�:E�&�6�HhrR%djHk6�QeC�ϷЫ5�k�Ʉƹ��t馓R���D��rc��1]k7��!�0�о��q����m��r��xj��Λt��zc�9��go�d��6�����{Cnr�
$�Z�ļ�AE����N�Tɭf���qJ4ɁND�����1�s�kU+�v~�G(��7r��t%ɵ�`�R��"��L��V�1->�tq�JO�'��:,� �1���ry�څ�#=J�Җ6���?}�W�T�l���&]��<���n%�u�|���H6��sTC�
�&�������'�	�L�=8�c
�~��-p�tU�1XU1�|O�w1`������q
;Bi���wg�5�wa�m�4
�$�u��j��,���&�N����W9P�6�.SF�x3.d
�=3�Z6���lC�|�1�H+���f�Z�c����hq3��M/�jl=������Glt�v5N���i2B_5�I�%���ޛ��ȇd������'�e����~}�X�C;�;ʪp�;Ҷ�gq��"���%�b{!{eY�P�'�-"��X8����J��ݵ� _��:3vH$Cl�L��ր��<0���E&�浓~r����E@3�wS����C����\�"��h�7n��0�dd���Y�<���(�Z[tb�b7Ő��'4�ܦ���`�@�I^��p]���ɯI��YP��I�Z
3�h�����1(�
��*2&5�8��HqAf-6c��bx*����Q޴�ދ�{x�)t�����
�7x����5���}�Z����m~��qv�e޷{�o�¿%OH�1U=�n=��u4�3%Ⴑ0r=�OR9�5C��ᑾY��+퓌"b\�=��9�g�L���ҭ:*�J_�����x	cB�f�9�!�AU��u��t)��bʊ���%��@�b�c5왏kp��X�)´�K\�i.|>�0�q�17Cr�a��e$�S� h�[�t��.P=�U,Pή6)�G��!�U�Q�U�v��z"s�<5.��,�u������[EGe����z�P�м�����4�w%�?��z��k�HxKf�0jY��OI$E�3�PaHn�m�s%����PNB�^��ol����c��u�rX'*)$j,7�<O��o�	�j�9?���w�'�/|�Ͻ����2���[_��8vy��n�)B��2T�4h 6���!L�p���p��dl�|j܂M�_s�g�1[��|��}O���Z1�01p��5AHE��"2���['�4n��B�x��[��>�rO��C�����#�7�P��*�o&>Ұ�%@]��!��Uj�등��KBGX�i�y���<RN$���$�w��>כ�Иxn �J�/xx(���؉Q~4�\��4����)C,�T�hf���8@SO"�1�vJE�ND�(�-4� ����c9���u.7�\g��F���,��c�O�I8-(��\M�K��j	��O�b�y����m.n>>�Jݿ��8�{P�1N� 6���o<]0�Zx�#�DSa���z�>�{��*{�\�������8�`�Y�R|ml��.c9�a��������1������e�I��k��g-�%�G�=o��b��7��A���p
�TC�M�z9_��`��PU,P�~=�-��i!s2����pf�X�m��u�{��5��)m�����*��^������g�qX�|=E`�6G^D��S\S����,EEџ�n��7}ǐ�Ɣ:I6�VȻ�����i����M���!17�P
3}��I�_|v���Q|j��Z:������	5i��a�/������V�� �}�n�T�W'�y�X��C!_�)����*k��yo#���m%yڴ7��2��޸nK�;CԦ���jrЉ:�ag3�H�Z��c��m��i�R���i+�ޗ=����!������[���|�3���ւd���Wu����e��T�l�E+h*-�{4��C��.����������x�#����Z:`���*c�E�q��1���"048��L&��9��C�ܟ>����$7��'0~��s�ڝl�٠m����G��\�Ԯ�Q�Tf-����0������y���m>���!�C?E�i��(	MM)��	B>�OR(b���۶D�/���S�T�eqT�	�t32Ђy��#�n}L���l^��M����	�V��O+���$�4q�����j-�:F������'�}�|����kzH�0J�Zk3����ń�n:Q����Jx�@6�:�]���W�Y�p�$	G};m��(�MC:��9��S��}=uV.>���iM���X[�Y;�l��M6o���Ynn�B�B-ئE'�q�)�5醻�"!|-[�:r.�2HZ�wj����e%���B���	�s8L�U[��][���F�����W�qwh`�B�dd^����Z�F������{/f�E��eI{���Ң#��\]BѬ��w�6�j��uɞ��.�I��f����:�mҍs6��i�	c��������g�c�ݔpIg��p������mT6�]k�!p���&M<��~������s<���h�F�"�(A�H�s.}!�P"d��+���[�ߘ �o��Q��#W��,c)�m��u�F
[��a4V鸯��Y�1�Q��״H�����h�g��G
��u�ʵ.Q�UM�l����-=oFFEľ�7#���Fm�)��v]�aY1���L �[��7�%/�<�:��c�Qϖ�=�X3��q�m���O�y�6���\�l�ч:0�0��!��O^dA���k�YBWx���?=<�ǇG1�Z�t���ÿ֋z�X�K��'*�N���71��Ċ�~�������)j]��6�)Y�k�&���"���1撠�� ������u������T��Q���/p����Y]M7us�I��~]���z_��Mx(R����o�4�sS�����W�@)yD�}�A_�<(��W%qrh\�)�e�w�V솊Ey*�h��U'�
��S![%s~S�D�>�w�<t�����V�o~A��N�DR�Ę��o��v��l ���"�h�d]���'Ch �s�pz-50g���j2l�8���(y�׽�͍�!����(̀I������ox5�7E5d��։&��1��\9��Pq�Y��C�����LOQ�n1�-`�*e�V�����9f���\�4n-y�=v�]�l3r#�������y>���nH�$�G��g��.9���t:����EئhS<�ٸ7�?w|Y:�}׭0<��ë�)��H�u��:�a�'yL��^6�	��{B���ɫ�l	����)Zm�!];�?��Ѵ���j6m)l��:P�n��M�`v	t��08������o�u,Dnx9rN"��kv��Z�a��/�K���\�wߞrb�	p�D���͡n����L���4x|,�?��Fy*1�4���ކ�<�O'�Xs�{�i�_�h	2ҿԫX=�u��Ĥl�/�,-ص����?�<t��ɹ!}lH�C�_��Z�9���[��L���ǋ�=NɅ�#"�2�V����6�蠟��=l��W��z�gO����D"�?�BӬ�Pi[��G"�Gx��ON3�Dq;���í�vÄ��1�W��%r��^+����`y����=�o��������[5�Ֆ�PWp��J]{���i?Dp�2��LʻwO�0�����(��h!}���A�Ks���~NQ��tYR翪T��I��Q�z�ɒ�5	��m���}�:�B�(�1X��h�n�!��<���t�:��$lc����?/�.ɵmq�ژi����^0�%�򊐫w�}+�8�8��݂�ZKN��S��i"(>'���11��Z�jFv��C:F�αɎf��5h��m%nv����r��6Y�Rh��A�xX-^�4��@�v��*R��Sϰ��[K�wx�6V��>�C=<��tٴ	�7���go��1O�ؠ�jIj�[��қԝ��� ͞,�3�3_1���z棆泊�݈�o���b�Z�p�Ί���|PĘ�w]c���*���0�`��'�$Kn4@����� ><e������\^ϯrZm�wUq�pH�)Q��=X�Vɕ��0~�yO�$<Xї��;����Y\hH���<�Y�xuP$�/q*�r7��b��ςk.s�;U*s�&3
�]6[ t�����T���v?�n���*�� ��/f�.G�q�����r)����^bb��E� ��� \~u�h"����)������� ��'>8\���Ky}}�n�Ѕ�Un��{����]v�w�qc8�U���ls�%0�[?Q���ϼ����U�k[;cPn�*k�{L;��t��*N������+�@�u�4��Wk��mo��޳T�}s|8��X)�!���S���S�98��f��u]5��#��p�D C��/�C�=X�x4���Eݯ\o��R�	�c���6��{�6�Q���Z��`��Q�߇�Q����_�hJ�==�ǧw�Ib���|��y~ѽp�:l�kWC� F�TK8�Y�$D�SV��XGeg�J=r��ޖN�K��Ѕ-Ns��v��ƴ$�I+��9�)%&%y"v�$8q[��ٓ,��>4RX�I�ٵ��g3̫W)�7�gcS(�xG�d���-<�������3l�&�d��A���nt��C�\ݱ�dZA�1kzeOO��d��.�$}��Zܐ�"e�e�d�mkγ�LC6�\����q�!�Rb,�œz�*�!NwB���E�0
a?cc���H��0�!��҈F��p9G>D�){��N��-4��A4rJ�jQ������F�!V��%'S�f�0�����W�A��(I�ꡋk9��bL��S狀q��$]v�H'��a�!&s<z�?�Q�b��j�N�����Hk�������q���MUClN�x����`ى����;M��8��{�u^���~/���L�Z�f�iH�C��'�!����dУ8�i���A�|��x<�$
��BaL���t��K\ļSV�IW���(��А
=����U�Adr%�D?n3����&��&�8�B��և^Y�0�0x�R��M~
4rT�h�?���U<��݋TC��1X��G/����-|r�iT��%+�U�A�I�aBY!W��A�����Ɍ���$�!o_���Q7R�/��׵q��P��N�����R7��L-aM���ᘻ�:~�b^ø�G�����6��+Ly��y��<�A�.'{�}��,�j�{�!'O�;z���1��6���a��n\/��`��7�������;y�˾>��A�Yts8�-�I܇�5��I0|vvbdm""�(�бT1�e��9=�v�q3�_2X�d5(AԬ|]�>�(���_�e���
�����>��-G�.`�bF"mo�^��3bqb >}����?1h�V�����<~�=�0�������}(�?|�A{y~1
�R�a��)���BL��ӹ�	I����mnɐbR�*�O��w[nI`��KlDCBٻE��p���U嫄�� $���E�0�O�w���������^���˳�%�3�ٸ~Ś��c>}��U�c4#�58T��iEq����|^��F��?㤪N�!%6�B�}s��8��z��6����Q�s�`�o,6-H�vx�H���b<}�G�}R����m�,v0h�U ��24){p�+;֝rS��@��	.�W��bv�dQ�L�G��G��_�e�Z~۟0,�������d���^����*c��O?���姿�$k�����|����vu� ���[e�æ#�Ӈ���ֽ����k�Y�f��}b�;�{x�N��k��k{���������lZ:��8�:�s�v��~����b��#->G>g-B���} �z�	l���?���~�������ʏ?*xm2�lO���O?�(#���r��<�{ŀ��|T,�h,ojݙ�!h͊2�v�Ԟ�}�#eA��&���� $7r��s�Q3��}��ޞ�����o�ʷ�����lsߔ޾	���'K��O�>��O̛(����i��wb�_6����b��C�oz���p���y^��l�{)��SO��z�0j�lph�@��+��5��??�:U�b�sz8������w!�����G�أ�֞�A��"��{��`�8`73^HhH��oV?Y�S����Ō�Ѱ�l,e-,#=��*!�a{R�&�ڮ��s�1ߎ=����G��3��Z\���ע����c�����������|��ɮ?}��B8O���dH�PgF\��;��!�l :o<<?�"x0���@D���"�I������U��{���2R�_�G���2�He��4.����c��V�I"����#c$UtR�2N.6���]=�OHÞ[y��,�m��������ᓉ-t�LT6���jwxf��]��X��^)FoUѲ:>祥�:
D��.*X2�G���!8g�X�3��aS_�
�`��A��$Ԥa��ћ�:̂'�x�%ޝan�v��V5R�/�R���H={r�
7Rº��M�4�^��7@5�kZX��9�`qÃ'hF�l�2�Ԓc̩
M�����`쿻�F���AhH�`��s�#S���4�LFn�mrLp��-�Gy��p�/q/>�C�@։ϛ���e*��"[�ZsBb�H(�����U���c���
�~4x^����u��gK\\�>� u�������r�R4��!�F�"Z��c��%AŽDF�x���*s�j2�N�t����ԦUpឍ����=T*��UǠ�a���M�Ի�3���Ih�Ϟ���!���?5���:�<U�.�S����<������������+p���\r��:Tz0C:	cݗ�S���.�-e2�|
>ʤ�]�)�u�[bߑ=D|��R�9�r<�e=��NQ�G�b'j��3�a��$`O,P	���w"�y|��8h��Ռ؋Q���r�=V�(���\��)��*�ϖ0*�F]"�J�_��t��p����]�ȵ�3��y`(�&^Z�nHcQ��x�����E�Xly�]�BJrjRc�愣��-�_�rDMa,�,fx�:d5��n���7j�����9�[Gwn��G޼�f���ݷ���T�������<��E�ȋ997�b~�T��5����8@��m�9���!�i�Q>��aH/J]�=v!�9N�e�ZU|Em�;&y��J�E�๪NK��Mvג�;J$L���%�]��{�?1�A���ΒC�p�|���똹�T�U���u�_^�5�b� �(�
���!E-q2���g�h�S�yO�*L!8^b	8md�ODl]Y^K�a�/���`6��'�F2-k��O:|�p�C=��&�&�N^����F0�݀b|x��]��_������>��J�b��RbV�*���!�iqc��?��m���(���qS�_������ �������|�E��Fr+�/q�th�#e#��5&���:�����7)�I<(=��(i�<��+Q�Jg��lГk�g�Yb#�Ԩd�ݥ!]Yqe�ˆq���נF���H�,f��+ƪkkp�e3C~�7�c!I�@o_�}-�y���kt��=�Ed�5����񮁙ʠV3�e�>��'P�0��9hԛ����z8=zv&�/��Y~'���8����_#I�'�	�O�R�CS���s�J�=��dG��l��Q���N%H
��/)a�
���'���̗�(_�K��b$N��n�?�e��c�Q@�$�d�*߮��?�MM�d���XӶ�)\e9+{��*�=ı�hW�H,vꍗɿO.��XV�dց�	�&	>p���z�������P7��G��Ȯ�m�n�R���)Q� �J�_öJ����9����n497��3�{xx�J�^�Qw��9�lw��I��}����9n��W.�u��dΩq��6c0�S#�E�݌��ǝ����b�r2)�O��m5�{�l�l���b��>:�c��+�����*�����E�&*m3���=�,������/��
a��/e5���E�A4����[U��ƍ|Z|Da����a��sX�pp:<��iV\y�<���c�3�,ɻ�������_��:��\�DL���~~�#m�O���67��w<�7i��G��۽�ڂ��fx�U.�Nh؅�篂���b!�bL�=�t2;9�.dbD�au�!q� �U>�L^�nY��I�S��D����I����F�F���c7i���MZO��J�������sx"�E>�ܷ!�T�),���i�!T�b]LX�Nr�~�^���BX��_�xtWgxʦ%�D|�m�`��Hn�]q�n*���լ�x���#�K&��A�Xj��f��<@�\Z����u���d��v���TIB���&LpЈWvVO���>g���S}����7�MiDy�I�q�z��-2/8�����I�FAK������j��8������G��j61���4z�I"7!ѻP�y��,��97����e������^4���If�x��ι	�#�P~�&:D����H��<�֭�d�����7�z���d�5.�$#�i-4��]�x��i��Ž*�d��=��@��F�P�[�|�O�|���q�M09�M�{�a,6!L��Ⱥc���7�-o�L�r�y���r(��x�-YiZ�������ӧ�f�aV�|�r��h@�4M��`¾Bl�1��y�-��U�V	�$�k�C�d�?~�Pϯj���F�Ϙ��ō䇌�E>G<=;X�y���0�k�9ε���!MۡX�Or���,�=$�F���o4��Ҏ�&_�	���v��y8�a�
����'r&mb-m����pzsMMf݈J�
<=�=b�#K�1ڿ���"����4����� ��7��6���2O]�L+*�"J[�(Q�?F,ǣ��T����T\��/�3We8M�mƞ��B)E��<8�z�NL.�$^�{�k"�>h�j2�F�  ��IDAT(�aQ���#�!������H��rL�p��\F�L1|���T��U�q�-N�%Q������1����Rb�F�q�s�&�z��04�ѱ���y�Y؃O�
�0mf��\I��]�=�v�l��Žϩ�"?�;L�_�;���/��ɸ�g�J�!��T�G�G�S�FL>�F��W�tU�ep5��0���q�ظ-㎃I����q ��^@),�����Y���Q�\��BGA�m`I�����l`1��u���V�UÛb�P�ƑBgH��� �g��5���9�R��2��ݶÔ49`��A��t:(F�q8��܍�վOp���Y����n�%��͍>d���Ðխ��rb&�nr��ƙ&�	5��>A�-���{gd�0�e���d\Y٨����OX����I�~�a��-�DƋ��\N���k]����S���P��L"؊�!=4�j�7v��Ho4;��5�#M��w��?N6�"���la[VDl���C	�b(��ms-KO`,���*�?}*����S�O�0�!����I��O�5��6�]u{��n���y��}���ӫ&v�0��l��92A�;�:<��s��u�
��d.�� o�J���\O�E�\FjP�7uUM��#�<*�G#�8h�A��ɥ�X�"47��}�0����I>�+¸�_?�������`����p7��vik�Ս-������������7$����s�+~����XIfj�Kc�;���<t{�D�Èk��sN\�<���5T;�q�/��}�9�p��|G%��
���$en�1�	mK�HBN|�R���d~����Zx�x/H�R׾�7�*Q"��
%����Za�j�bo B¾�'
c-9�w����4y�#Bv�l��B�ª��~�m_K_���OO��8��� [�KC��
�������|Pxg��xs���4Ҁ�K���5�Ӭ���W�w���b��?#B�\�����?�s�ր���������2���f���M���d��.�ѝ�/w�=ޕ��M�l��%{.Y�W3�f������p����q�-�Q�adH#Vc���j/z�P�/�X3��4�G���ٱPO�䲬�ү4�/6<�Փ��Pl�]�c�da?I(�y�>��,?��6��_�(��L~�hFH�����LmL�_�s:��Yq�bz�c1>�@�b�������_ZoD�v,y�qW�8j��g��zY|8��ϳ6;��%x�0x�V���V�&W%�@Ė��;i>�(�{���t;� �����7�}����zR�m�T��~���y_��0�r ��Df[��h$�f�����X��
皑��d����vu�'�>TQ}��rgA+�(b�'>�
n��$��'ג��>&W��`aJ���@&�)�N��'����E�Tk���j��چ�Q)5Q���H]{���֖������c��ݐ���G��U�^��?ݳ��j%�����g駏�7S�@�������q��7*���mS����3�s
�O÷?��Η��R<%udu�e���)4*����^����g�����>_d�iS!�K��܈��?}�h/�{�4⯬�ޯS��}��#uQ+�ݪ^�E����]�����wØ~e�������I5�;)	��U�	�S�CP9�7�-�G��D�R�Q`�f�!顶n�f�b�ɀ�]���deV�>sd��-���FeN�F�{�Rا'�`�P�bt9� |qD��IAX�����xW���?�u��g��RR$�=Fy+[��d�GoU=��~��za8�+|2.2�M����<�sk҉X<�ZH��}� \�1nl�E4��w�Ϗ�[&V��kP����!�=��n����K^����'O/I��Bt�@i)�^,2����[��@�B�y�����$���#���Ӎ�!�	'���7������O팧:�g��j�#^�>��8�f��!<M�Dm:��ƶV*w��WJ<2��9����t{,T�"��D��!n�9�u�'8�������a�F�����E|�8�Խ�b<�f5�v xv��(�*�*�*u���fI�Cx���R<H�����i�V�yS��n��c"���嶣	
J(�u�C7r&aD?��Qx����(��i޽)�|�����U��%���&�Q9�jH7����.a�x���%�O�u��\�Z���i��)Ҋe���~�\/J�y|2q���֮ςJ�r���G�N�������ua����t|V��,���eJ"��L�R��T��X�,�(�L��I\��M֩e����[<	����V�͞�А��(�9��E�M�d���a�Ae�>��^��l�G8�,�F%ԇ�zh�~�)������͇�����{������=��Y8�?�?��*��ɒ5*ް�������s��b�%iY�Z��C��x���Ԑ6�cB�N�3k�'%��q*������"��SH0aS���ּ�3�_��<[�':N�&�p�_>�*���P�=sêR�R��+�QN�Q�s��K����a�7j�0��$�?j��%8&��{��^��V*��&C�,Y� ՛��س�4����Ud�?��IgdPђ����>X�IK�:�嵑��qL�s턈�s<�\�*'�a�5��=I�u�p�
�7�ֿ7�5����d8�0 w����I�����ɒ�����<�ށ�U��I��ε���0Rή�tͥ�X�29�j����E���+������s重A'XCGK:$2$�����k�p��Um��������`D�s����ũN�vv@�b8Ǿ�CT��̠�4'���,�ɉ�Z����#����d�}^��E�N��T���먅�~3E!�Q�t� �nH�R�*1�~�R�>��1�$(�p��f̬�*ݤ3�����R�
!����\��"��'_H�WE�y�[Nf�����?��_>�2NM�֭t�qzO^�#����&f�dQe��/?�"#�P�Z��c�a����@�PZP��0�2��U�_�TeId=� �ֵ�ٓ	�"� ��5��ʁ�������8f��F�h]��.]�L0#ſ��/��P��Ƥfu�����ϟ�U�����Ce8Ǩ�^p�g�7j�z��˷��7���@�	�A�Z��M������f-7h@��m�oI��\J�e=�`f�X�v��y�p�G/l�l�(��J��S2�z}��g�ޱ���F���!�E��M����܇���������!�R��s-��CR��%앟����ix�rt��(��֍�p�)�߱��5��m��$�9u��8�۳!�)s����1�[#�{��i�]y�u���I	)���m 1�F�Pu��gkU�]�췔e��^�)���'�X�:/U1�(�PK$;`p������^�U<2�"|���er�dz�T��=�	���'x�P���G�}�����`�jD�������OfKz<�l,"�"t��Z2��h
_(���O�)k�W!�_�n��]��a��c@̳*�� �⬙j<O�	��c��ƨaH_L�t �3�-B����\b���#f��XT�9�ƽEϮh照����=��L��X��d�[5��m�St��N��Ʃ����c��Eqf�-y�ԕ@� �]�%�E�\����h�&��]�L���9O�g>
c�E�uMH��Gx����mo-yÕ̍�Rp���32���6m>W��dFݒ&�����$k��k���B�u���Oz��ʆ9�B�p���yZ�uw�O*h��B�u=�����{��rk,
iN��u�Y�P���o�Ye��@�|44Q�vR��8�I�t���/j9�Si�ߍ�Y�ߑz9�C|\�ׯ_$)�m7N�߽>��Y>�W��:���e��dNVBY0�i0�K���J�Qx��H��h�VJ�kٱu�.�0|��gfE�_A�bC�u4��Gz�%��Be9"Ssz�m��)�	~�"
M�qp���k�BX���US���
�l	h{e���i�Ģ�w0^��[�ډf�إ��_S��Zo+��I���fFP�mR�����wL�9�@��&t7هK��л��R6��J���;�>�á
F�e���&#��{��G��6k�-�ĎD��TY��_�*׃�KR�����6NO�G�\2�ץj�
%��p/���U�C,�?0����O��@��T[��kp��5?M�Q�c���d��dڶ�B�M[Q<i��Rj�������Ré��$����Ɠp�{�È���{�\�|��Ѐ���e_�ʣѾp_���aKT��b�Q��X�Ij�.��{Ql��PI�.Z�c/26�s�T��Z{��]t�Naf�1/�%�0'ӱ!�i����z�(x�ŧ��PxCd��� =��J[�o[ŏ�Nso�c4IB<��h��h`���m�n �S��X-)��}v�9����q>�~Jv���f�B��m ��*�}7�-�q-��5�V2�T0I2F�)v��o=Pi6stn0�l��m0O��Du<TpdQ�e1-U���`��:E<���m�����.BWk�)զ��#��f�iS�#:'���ܨ�Nt~Uj�� �ѓ�����ɸ��`��C�2��L<�0KI:`���aSO�7�J����=_:�U�
R��g�?4�>���`�}q΀c���U��&��U�y�Gg�2�����AoFg��j��a�5�p���(+r]X���e2����QzLE�.I����"�Uct��	HlOjܧ����U��h$
N���ő��D�5�A��{�hK���篠 A�D՝@������ڷdSE����8B���<*%�F!W���qEpS4�!���/hOtfu��кB�r����5 �
`<V�T[�i�c]͘�G�%��>|f0z�� 	��)?�f�Kz�R�j�S��r�A~63"��P	0�(˵�t��$�TŐ��)�����Zy=E�Kg�|kt�b��U b�#�G���<t��₯j�oBkB/<�P*�=�I���{r,���;��R�E�*FL [��a�7srD(����x�4�3J`�O&��ywN�q<#�!�ed�������jT���U���.I�޻*��tk�A��R�̺��X*:��}Cٽ��j��q���S����yk�9����e[aj�@y�|@�4}Kf�J�|�m"�#��2�A%Ho��R��;zULP�~���^Y��S��B's�Z<7�GR�Q�X��+����jNx���{+N����~M�e��ɿ5֐7o�M�ʆ�:[$�(3T���wjZz�Y+����g҃ƍ}��`�rX����U*�t�	�ޖ�{3H���ZJ�����>D�k٠�d���P���b<b
���QHjm�5�o^�!�;��ټi �!Q��x�E'Ka��>���(���1q^sӡ�<�x��ڇh���z����zc�1�f���+�3Z�O���OW�Ru�K(nZ��J߫	&����+��&�\��Q�kkߞ��H���7���n�}�lָN����q��s�,�,3�Ÿ\p�߽S�(6�l�)�m���������o��vF�a�z>��Vv״�mz'�7���GO�I�#��������8�[�K�u����\��U���M	��j5Ȟm��Mۙ��#�`�(+X8�4�d��G7mӪ*�<0X���>��@�&n��^����}Υ����*@S`of4�����zS�[5�����G�K�Q]���iꌌ|F�L�=�7�o��Y���U�"�roվ[J��ci�=Ɖ-vrW��D�����"�
b�jݵ��X9ׂ�i=���M�ܢ��`Lp��lO��O�Ol��uc$J�c7R�o���n^���]�������6ڰ��T�t��*Uj��Sz�,�&��B��՘8 �#��y����
�g�X�}�l�LN���yeӦ� �]�[��݌�x��M)�˦z<F�1����
�"~�ԗ��Z���}UHk*��p��vN��Z�H����γ�d)�N��C�����+����:�x���@���*��Fw��pc����\�1��#94�6��Q��D)i3G����P�d�#b��э���D筳sPA��a��,��q�6L�P1�Q=X�e��N���EI̚��^ǌSJ��Xo�L�ζIyBx�-%��5B�،Ψ<�D]���@P����'zyLv�CaHs�?�!�Ù�Wcr�= �3�?G�����j��MW�V�kS<l���U�Ӥ�ެb1_�*��<�IOi'n���b�,���Z��(`��ex���e6��bD��u㝏&�	�
�@S���A��4B�0��SN[b,����	��zF�Y{/1Q��׆�����������<�R�D���K�b�o��}1L��h	@���oE(\�l�Ų5�V�34!b�آdq.O�i��SR�Mw��,x�!�q�s<���ä�NNp�/3�O'>�ҳ��U1�V�EJ)2�e$��j8�r�Ǟ^�@��5�Ѵv1sp�G�׺����}7���ܪ���4�u����	1�>V�4�s��e8��ʹ�!�u*�D�1U��6��6�m|�GHơɎ��G�%aX͍9I�j2�E�w��NQL�, �5��9�l�z���k�@���u=ߗ�^K���2d���ςh�h	92"<�������z�k�y�#�g�Q����)UL���C��UK1|YjH�"m�Ӌ����CI����T��{���l$�JZC�?~��hI�A��68�N�+C�@=|��k�ڊ�7SVk�+vZѺ�`����g�m�`bI����FCB�H�8��	X�4S~zg��RvH/ъ���� q�����${ T'[K���갉��I\��z��RG������>{K��)��frKy�A��{���!�^U�m�Tn4����R��R~h�y.��S�ECv�uæq��d��z�kִ�����0zľ�WJ�;6F���H^N~0�Ţ�&,)�2^Z�eݺ��$�b��1��53��q5��)�^�:�����}W�'��l-�4����Yᔢ��2���T�,�%}����ZUܙ������giqc�5�;U�� Ts[M��(���y��0�%5aH�n��©n�ڣ�@FT��YP�eޤ\��_��币��a��1���ō�K���;,:q��7܄����1� Qɉ����G5��U����1�d\����Vh�x<�0N��4�E�F=W���a�dJ?P���О�B�@gC�������gk�Cs,|Rz����]�Q��~�1���I�1;Ob��Y�sSR®ʄW)��,�?P9���%Ww�F��q���4k�� �l�d�B�o��������Y5͆�m�����&���U̬3�a"���t@���08�c�,�s�u���J���_�K%�-�5�\3F����Z`t]�*�'��V� (.���e�F��>*vX6�9	�+�:e�KY,܈�����p�0kv���h�+�)�=KXԾQ0���f�͜0�M���by�6�li��F�R����sc�/�c��]�$M)��g�&6�͞�FOim�U�r?;���$�<�o<'[��p�XJ�����p1�w�M:�Wt�B������^��R��dH���5������΁R$uC}�>>�h�PJ�������5�.{����8qPUoJ᪇o�cB�
��ɠ6�1�%BzϲZ�!�j������Z�,Īz��E����%�X��%�xX��V�^�U���i�k!Kߣi嬲p$�@�Gj	>�ҪSn��41BaiN�J;����W(J�|��[�R䟹:L��qn��Q��_{����B1|���kr�D���FT&M�U��>���	�J;��������8�Exs/{V�Ұ����~���	�WmϬT̃Q�L�js�����=���%�!��#%ĉ�`��d��Nޏ�)�|a��Uh Ӡ�}�?!]?��s�Y�h:�a��X�á<=<ɀ_��ȶ���b1��4Ŗ��·��}�<>8A����=���§��
�b����2�'��g��w&��*��s�@��.�Ҵ�8���P��Q~oSVo=�ߞL��h�� 	a����$+����e_@Z.���*�#�}fM^��m��r�+Ġ�f�0���,M���`:��W�C{ETe������!?<j�$8�����j�R-m�jg�T��Rs���C��9��[1��X]#i�:�����ۊqF3������mD���״��z�x���ׂ��,a���d-�g��j"@����"齚T䐔�6��|h�Q��FO/Č��R��y)��l��҃9͠��4�#�1`r^o�*���Y��{��.�;�j���j����Щ���L%����jnp	�)�v��1�P�K��y�.ë�]M�C��$��Ӥ᥮��Y>Q��ܖ7_���7)
������(k{�+B�0���I�����f:Z�#'"��M����9�(�i���n� B���J�ߍ���Z�o���M�6dP^���GA�a�h�c�q2E(-��bSa^��yz,�s��x�C�FO�ه��*T{T1�&ɯ�GzWKNmV�µ}P��є�1�l�9O�a�ч�M������o�ä���Q%�mhDGr�"\�V�G�z	A��Z>��Q]A9�a�Z$Yv��}5���xTc	[��V��������I�����D�P�1�����dSxV�zc|���Qc���ۚ{F`�5i�2���m4^H��w��C�l�����,��`���SU�c�tX��L����K��-�3a�j�+ 5�#�MOĐZ)�"�����hkEZ�X?��4�H�2J>��jҪ� ��d�*= ���^n�|�4�E����
8`�וЊ�g��o���E��U
y�pް���������óR�o�9�ժ������	����X�m�^eFu"�3\�+�MQ���`�T�f��q�t��G+�<״�)���3d�L$�ʖ+��So��nH�=/�Q~�Y~f�T:7�«�Q]̨�PĦ*>j�Լ���{� �Z�G���!-~�����(�s�� ��J�I�ʤ���]';(����� 	.SWp��Swj��ah��}���˾��^Η�x<h��~ߨbD}JB��E��Z���
������,�s��I��}\�l��/�'�zY����B��*Ǉ�X��-75.bH�>��4"wJ%~m扎fL�P?�Ʈ�;�T�]�O��@��
I��6nY�\��.1�ܓ���N���X��Z������õ�߬�vh��Z��71��eσ���p��D����R����[x,I�M�OK�!i���rLi�����F��MǶ��!�1Yl]g�(�K�]���]QL��4�i�=��v���ֵ���8J:��`9֨x��Zh ��W���n���C��}�њ���E�2ȑ����B��5��m럛{��mt� .�qp�V�\�EJ�0�1��8P��0Ŕ2�hb�x=��*�Do�*��#��ʦ�.��Dn�8�j*A�탏��`*G�&z�.��ƞ0��x��S�q�k6������z����_z��'�Nţ?$�g�eMH}1Ly2>�������Y��R3@jd��sk��P���`)���H)� �E��^K2�&�i��a���-�\�	����W-�[�ӝGZj2zz}���A�j����!<Yō)��u���[�7Z�lpΫ�d	�#�!�Ca�������xh�M��h[���*�`��,�m+��T�Jb�����W+J�Aov5Lu��|Uᝫ�d�;�Fd�8��E��{�G`�U��mm�a��hQ,0�0M��U��]J��ɭ>��	5���դ_D���ZG�A#����m�A�|˝�Vh��
i�bP�(�.������$;�^j��5B����l�X��3�#�ƖR_��/PQZ��{�fq_�|��RE�'7.��5���ڎ`QS!�:��eČ�J�M�vM�g�y"�����Ed��d�U�M�]` K�Hk�1zM��CL`��G�A$��P�V%Q��?�� F3{W�����C�������og(��@=�����o�trB6(Kt.ʰ���q���Fq�Az�|�I%�����A	�7+d�X==�׵�Kf]��V;�j4��ã��o)aFn&�T-B3z~��)�����L�D�7�B��uH������e�Y�f�S�Ha��ǋ;��`���t(�"�e�aX�{��.�O�˥W�N�$�NQ@T����'S�>����ċ�n��k1Q1�=��^��˫�$�{,��aAHE��M=�q0�~�8UNL�@@B�KD�U�j5Hn�+Z��|�Y�i`��)lm�Z��76���k�/�I�릘���-�,	����]�{�P��Q;#��Ⱦ�;��}D�uxrb-3̓QI�u�
�n��/���m�����U+	����-�C�r�ʪ�8w$��ʖ��CͶB��֛~�̙/��˙�ua�U,M6��!���=N֔��������E*�{(���j:�x=���C�`6�&X��}��Cpk���4,������2�̧����d�Z��j���>;�F<�z��:��3NcC��� c�1��n9�Re��-B5&oj���W�!��٫*��Y����rP�������(J�/��^���T�Ζ.l��UPG	�WH�]�`�P
�kMX���W�����A��i�dh$ýG;FT�Pr���_e�һw�c̱���J�,5��d5 ��)�m	5�/��f����d�1y�7i��R�}��t��<jK�:���v�＠����������g��Hݰ�P��m��#UO�RO��(��_~�E�`I&x;#3���>X��b��7��~E�#��iXoj�2�~BC�D�"N)���EPG3.'+1���ż@�_�񽸆��U�J=�f˛�r�?|�(τ����G��â��F%U�e,\z�� 5f��v�4�1�%���jI#�P�s.B�P|J,zR��p3"��j
��O�<u�7O���xh[�t1�l�j"Em���W珸�����(p(it�W��K��+ŏ� 7m�
����%ONf�5�5���Ƃ�Z��ؼ����*�h��֎E�W�O�1�5���˯��"����� ��Jj�B�N�n@3k�g[�ë4b�H�C�j��r�����T�lT��\j�KP�&0q��_u�Ϯ���.�M��_�����עB�B=]�CU���l-�ci��I�����PoC��x"�z�5��T�Z�i�C�{n&�A�<"n�5�xH}��4���e7��e��zz��C�a�ELFq����uY�ۉ�Y�?�	�	]Mv��b'�Bƙ�Mj�4�;����?���m�n7��A�1�⡱�k����?2.q���zޫ�?��5)b�����s�O��ū����k�4�j�DO�h;�� �m&j7o⼱�p(ݸ`��b�-��H�YKo@���iZgH���U֣����e�L���-�m�V���K�1�w�v�41��ű#�a��o��!�s�9R�X���⼳��f�<3�Rμ�����u+���b�u_Gg��wV��yI�+`���u-֮=x�wb$��A�ĳ��f����
[�H�Dg�lڪ��՝�:0N��+X�P/&Ծ���uއ�!��������=�k�	S��|b��H�d���F�� m5�|Q��t�MC�,��T��������y����PA��B��׉�'ʖ���$$&��K5�JR~!ћgT�঺k:(�P�U��kׯ���1�*��qCZԸ�l�{�ꘁ�ߛ�����i�	���`\ԓi�Z�DTJQ�9���we�ٰ9��XIi�n�������7&�b�x�n�量Wċ�%RZJ�ϞT�O6#<�!U�S��5Jq�]^�6N��Q7T��<5����H�\I_,>i�P�.��R�R�V�xEZz
���v��X��?X��� b]<r`8�D��U�RA�u&�R�H��4�����״�i��'x�b��rh��]�z���7�a�w�\2�t"�fr���ږ��"y���Q;[9�t�R���'0TD|��x��t;S��l�0Po�@��Kf�pR�����W۲]NY5��A}��@l�^m)�J�X�]�n1C����v�Ӗ�I"^�J�Z��0��:)ߛi6%�qd#��y�P��\�0�8�U3�����س��0/�ْ�S�Q�FLi�Zc�v����W�4N��'�Ji�UZX_�5hYQ�0l�r��R�B�h�Ӕǹ!�Ny��oL��+�(��<!7�C��/�	G(����o�T/��3
�k�j�f���ސQ����3���?����sd�D2*�Rt"Z����`P�.�E(b5a����.�DSA:ʾ:kc+]m߽+�?|c*F�4m�>�N3�L:�fHI园clW���Vg�LIht*L�߫���sZ�]w��BJy ��'�f=�7<H��3Ƶ4pQ��`�T�����Ū��!0W���ئJRl�����já�!�����K��6�w��/m�͋��m�L��n��J�� @TJ��Ҷi���e4�W��*@�,x�Ha&W�Υ{��u���;h5�%N�24�B������OdD=2���������V�x6Q��Neo�l'�����0����4�[(��,F�!��;	�᭛�|v/O0Kc#CI����Ѩe܌ղ��������Ca�h3e��24VS��N�[�U�a�����?Z��}���˦-���=�9�z�Q:�����
[鑆!%��@#��)���L�ө�H=�X7,�Dx���b�n��+�e��~�_5�%dt� �=��ì0�(�'�w��"iz��\�b��y����=ca:E��p(��I����Q����}��_���?�mn�G�lи���Y1y�H3˅�3�o=R�rwƱ�Y̷���j��[k�j�M�(~8h;_����)Q�n��ꕃ��.����7��oK��q�i+Qן'�Plc�h+GA�U+C�ڿ�^LjP?�O�]�ͫPzEm5`��.�$���/]�2���Φ)<ق͘��1��H\X`L'�c=��3�C�zrK;t�B{b6=Ofz��C��%K�p3p�`A������emH)�C�D�( 	�����"�y�����I��[iu2�;�E��|Eb4�u�M?fZ�H)I^���wQ?���F�;1��2��<T�d���G�`&������*�r�ar*��������L�_=�4���KU2W��H��Ƃ�K�c3,Q�$0��Z�%��Y�)H<Ѧ�.��j1E�ϫy�����Y���.�'�۪� D��S*�j�'�H�`�OD �:\7�)�(2�W%��-�a�o��S���;g2M�{����eN����!�P�H�D=��GԳ�V�0���4�70�U���`#~�Ŭ���48n��w�%�&�&�$f����j��l��Q3�}%�bGʨnbop�DK�p��A	���;����xM4��|�����J�]ʇ��G�Y� �01�5�[�ɐ�xR��h:�u��X�K:8R�,�/[5����g���]��������F�����z|\����C��b�q�RHzу�����d�Ӑ���d�zJ�U�����|0��M6���-���MQ*�V����ĈN���j��Ѝ��HkQQ�}�q<���10w�/���S"|n% ��j�u��� T��O9 *��͕�T�I��(�Ŋ ���G7XjH�I��X6܊
aa��!�3K�^(��^��XiL��i��>���ʵ0L�t��w�T�a�R���	�h���n";)�^�{TS7�m�ʹ��,e��O���mi��Z#�����aU�~����b�OM��O�{5&z����1LL����LQ^y��T=H�����H�4f[����%��f �Ι7���\B�S,����hl�SP���q�Έ�� ��Ma��=�Ź��?�&[l00X�~�c!�Em1�+X��'o%p�U��-VP0����9��@D��R�o�-]�ܯ�������Ÿx���o_=���+�$�k�*,��ãy��x�b�Ce(c]/��+B��M�J����J�l���:�)ITU��b��d���YՐ���y�h�E����8m"ƣ�CE���u]��8���K��[g�L֌�&\�I#��j�1~�6��t'��m�a��p>ԛ=�sT���#\�x�r�*��������ٰh=��/_�����"M��B6�ꑑBOG�WXV�]�u�|U1��A�(�u�
��z�/4q�}<���*3�GG�|K)�B��Z;�V3�az���dh�mf�2�?0���#�i���@�i�Z�&�Cy��zɖy���^�����#I�"r8J����c�Ci :q���Mc2��������n`��eRY��}�e;&zT��-����v���o틭�e�a˂ـk�w6I/��W�u�QO�p������ӏ��p_�[K/W�̮W�~�=�x���E��I����B�&b��X���J�sex�fՏ�b���D�';�4��}8����`�~�7�Ҁ4٢��,�2�JTiZ>���P1T)�02t�p�e5��(��K�Ř7fH�}Q#�r[4s�6�øfN�qk\��b��XPN��tVo����سH��B1�! �|,�ǫ�#��������gŅ:	�U�'�����������>ȸ����A�k�b�X/�~����͏z��umy-���݌V�㠐���Z�o�*N���x�}�o�Zܠ�/��"�-S��%�w��V��Lո�z��(40M�$�`��;~z)o�����gZx�t���ܪ�ʗf��U�4L���
3>h#|���5�nlc�D���XX���'��|2��<����#�I��<3����JC��yf�6%�ofH��z�cKb����p��h54$�y�sY�[�k�n�6�c��4�t�����?��O���?H�
�X	����U��?��,�=_J��84��9�)��'ث�tٍ�Y�M�Z=�H�RjFxoH�_��ؐ�o�-��e�s����$R��7�W��Z�x����Д|�&Ja��xJ��Q<m�B��M���#0��M���i��W�*FN�4�Uc:�uVN/Hv�i��s$)�������ہ�CL��,�"��jQ���{�����}D)H��*��?�]��~�8��Y�&M����&~Fet|ch���{ߑ3��������vs�OKy?��;��]8�6Z�7���"QC�kReP�D,�&2��"��][Z����3��]oC{���u`H���~�v�{0�՟�_��7������K)ZY�u7��O�5��;��<5,B�r���<˖ԙj5ڍ�
�4Ƥz8~��l�z��ܚ��J,Qf�Đf�up��w��LcK�F�������:3_����M��\��c,���ϖ�G�$�&i!�A ��x�e�="�<T��E�����CT���ry8���I�v4���ߜW�Yr�LpW�U��U*����YaƚvQBGc�����-�I{����.�G�жf	Γxc,)h�X�J�MM�Rr���I˜��L��b�Đ��ek�\��a؂{ �����'�#��
��g���}(�?~�q���_d��o׫g�5IP�NF�:C�[��v�Ƅvb��~�U�ᒯ">����|�$��YD�:����s"X�Z���Š �a�4�?)T3֭��!hs�=����h]"z��zt��Y&�%2�3Yk�at[�����m��LhoL;�Z��l�w����xs;�>v�ZW	�섣�Q�H؈0E�
�bj��&�x2	ɸ�Vb�^��S�!��ʷ����+�$r?�S/A[n��b�A��&
{P�$�b�� ����7��8��"!��@<Si����x�2�3H+6�EJ7a@�U9Fwt���vՒz�=��'��J1%���k�<�CK<�jٿK*�d�J2�碛�4�&�{tC��0uS2�0^��h"CiH*\qxÀ	���)�r�5L=̲xf^�2�|Ґ�#n�#�<�e,�a�<cO*Y���ma.�J<�B���)�g�PH(��tM�K��֦��"\&�ޤ'&a�C�����Yg�~�۹��aӹ&^�u�L�T=lD{�)��(颂4샦̍�Seu��}?P�
�1}=�,{o�e��9'ՄEߤH�Jc����8�8�Eh��}��ù	�h�j�7�	'��7�����"�B5 ߪ��h����EB�}�D1�d.WK<�K��{V���s�v���h�<��"d��� n�V�(�I�ϥ���3�LR3jƕޝ'�������]~Ag;e�Ԓʁ�贿~��_m1|o������B5��}�o<G�X���UU�����_��p�G�Q��τR��x��|�w�r�'{O�<�(�T�d���_��Z�IgR#r�y�&-�� ���u�M���0H��oQ��D;������8,R|s
�N���Ԡ�
�����FՋ:���M ��a��Ć���K!�f^���Y�2��Y��t�b�`l�����b����R��ݑ$G��� 򪬃����?0�����/;�&����k]TD�<2��o�De&��������;R�.d�\����z��������])�'��E���k�]{I��[Ș�=A���a��o��lr�ܔ��J#f�U���9\�����h~}�O����.#��J���W��
��aѮ��^����
�.�އ�����Yi�S�yJ�H�D�5;�3��	����v*�fbs���,=�FY�����h`Y�'�L �v���X�I�R ���43��*���^f�K�5���SF�4י8{w ���l~����vL��
��k�h	��c5��rMR�Zn���7�9��pL_TfK٭���Р�����n�Ĳ����n]*],�0dI�ȼj#������Z����-�����	+��--�K��4�\|�i`�i O[������eC�h�A�Cp�9�e��@ry�i.WΤ_,��'�&#�I�Jgr��Yκ�C4*�-�\|#�ȝ�O��l-?W�{�B����?X-=F�2ܕ�C�� ��?��z�ʻw?m�����)���0�!�̃�"�<���<�pZ'�h��^�����k����z �@?����a��t�Wдޣ� )�m�CLzx�����v�����N��ѵ���+~�C��u�@Js�SIO�E��0���C���L�ӯՇ�>����?�H3#m��A���lf���	D�y��A7�,�N�;3��%L�޹؛�a7�F��Q�,��i��l����=6�4��t�w8���nU�����֯��
�7�*��-1�h�!�Z�]D�vF���=���c�Oκ.wV_�����s>�'u/������eGsjd7�D?}�F �G)�}_�e����<���}aw����o�����?�}���mz����t*�MU1�>�枲Y���7o#@������Fm(Ϩ:��1}�z��t&�r��N:7S��v�4�p��L���sr�un�X��NP۟�p}�_ca���D���s� �O尖��c̓#�����$��X��9<���u�-�"0`M�_.�_���;��H##�5��A�zӴܿ���df����wp��kՐH'�Ӽ��t���8^sO��nt8�eL��͛&p��9�6����0��R���%��VQ��,ý�X�V_`����Á�o��a��w�޸�6�}���?����wi�.#�۱4�T���:pߒrR���.$~�©��¼�;Gj��1����8�MK.����ƦkY��+K�l�i�%��Ve�f<���BXJ�_�,q�M$�mf����}�O�-�z�X�\�b�h�,`?.�nĢ�먛]�oA�������7e��tX��zՄ��|����LK�7�&�߂h��Mf����;�zh�=�Ad���
%J�q�>�fR�M�ދ�1694�:]����+��'�Ӑ9T
{+�,7����Q� v�k�de���=-^/���.��jRIOn{;>�"|�/����ً?|�#�,+$�+Ma�KT�� ������#X���m�`x�Df%.݊U�����1ف�.���6�������6�ɱ�8h�����3����J��=.��Yi91���\�l��������k��c9��^�D��+�c4���B'��=�q�+[��͝��?�;�ӟ���3R;t��������S��D���yU�t��+���O��JA��6T��vA/8�ۦ�ʌ �bEAT��H3gP��v'��\ѣ$��kn|�NK��5�M
J�-H�l,*e��UW�a'6؎C�l�n���Ȱ��	(I��U3�([��	���>��p��G�1ɑ��8��X�bbD�m˦�o����ّ�|�t�������*�l����?�/;�J#��GI�	J�#�\�;�J�^<l� 69����n�#�0�M+��j._.��l0J�LmY��^�J����<�A���4Z5��8֣6 �^���qb��~�\gsE�t�7�@H���Η��(q����|\�qbEC(��c*�A�����{��U���>'�b�9�ơ�uM��xj�uXĢ����π��
 �A�O�[X�ကi�~/88��2�n��7ǉQ�4�G�(��y0T���.����R%��,R��K���g���?X;��]+���s��av�d�yR������e?/����Ha�$�@�׃P?�ܛ�N�Y�c
"6�r����<yl?p�_tۍ�@�-X|:�l��D�ؘv,^!��m4��x"�)26֘;ŵ�yD��4�fQxfe��&�n{G2o��F!���ow���$<��&1.����R�[���K��_�'V�Y�5��^
��,�b̌L���V���A_g��2��H��ImsR�=8�:��q![���-�?C�S�ݭ�]F���|?��dmv�ﷆG�,�\8J�AZ� �Z�E�Lo,B-�1�����Q�2k�8��cs˻��E���������+�O����e��P�������W��O�JR���ӻ�}�>��c�S;׼��Xm��ٳK��W�伕~�n��5̮���H��-�`^2��p�[�g�a�'��i 3��8�\v2W�~��Hϲ�:��$�����o����˟�L�'����x��yIB0i?%O�t\)%���p�����Yj�H��wYe�u�Ԯ.�>S��ߟN�]�Aw]Z���ԍ�&�*45�֤}�>Q�e�b���
S�j-���^�vS�(/ڌSIHV�;���V�J50nM<��Ԁ���)~�Y�����b���"�y���M�=
�)��CF^%,�ospa��P���YY�,��9��u�Ԭ9<�4NP=)�CH���dH��5��cA�8�������B���ɓ���u�>h��咢�s(��p̂����Q�����C��dh4O;6��QϮ$lJ>�d_�9�W���m�a��O�,�Q/��,���C�����؅*� �榉�ƗKޗ�	��Xc|����ᢱ������|�K�x'�1l�y��I-�c�Y�D���v���M�GZg���X򍱑��TF�VJ���1�fV�,+1�og���y�9h�NT~4���F]���öR^��|9{��I�l�La��ŀ����`��Qj@M�ۀMs���gd�m�צ7��^��- 6t�����.��1tWr(��ţS�,tQIn�4�mи���eyǒ,�FY�R�*�g�rO�nHq����4�<����C��Y�E��%�� ӣ��jd��o�d��H������vc��и�s�!x�7���3a3>|�(K,�ƵZ�DUrf��������qH��Y�ڨ`��5� ��a���� �@����UT����ǿ#8˶	22�:�H�r����BM��l�с�\3���h�g�#`����Vt�����&n�-	�f��S��-3]E"^`}�����������P<1��i�
jU�Ċ�]j3�<v'lv���z����V��w�w�����X���B'I�;���Mf$��, ����XG����{7$F�b�@� �v
����yz.;m��lLU_�!7��>h���[k���K��O\8�C%us~�U�/;����!��42�X`[G�[��\� ���ʚ� �va&����uޑ���#�h�n_��h�d���]9��j�9�e�8�l���A����z���y��3�M�O!�|H:�ihd����an�x���
�\CS�d�J#���Aԥ�Bgs Tm�z�wwz�]�_�𻠰_g�T�/�w��Z}�wQN_4;���p5�����\gɡ9yt��#<:��$�t`�[�̾D�������T�3��볭�����S"��zX\7�/#q}�n���xnc��G�]9ዯ1GfJB`���%u|�~�=a�j��{�VS�:�{�ZhZQ�����y����z��޿���WC�T�v�o?������Q ���Q��ZjF�uҡ�F�7eC���n<�/z���u���/�9�O9�{�E� ��<NQ����1$������q�7/��Qb�ӑ�� ��^�͓�Hrwu(^ˋ������Y� x���:��w4�62��p�&]7n�k�� <:�u*��v��L��|?��W)T2#�f�vE��B,�����H�������sl|�ldg
R��H��E��$v&��u��wx#}-[56� �;�����Q�4�84��
)9�����޲[Cn�N�\�'�JX��&�����c�u�.)V�!PVeշĽ�!�D�%��������Z�#X`�Ә��j��ُ�Hec9/��3#�5]�����=����q�W�mG-��:�z��f<�Y��O��h�:�T�]D	����`\������s|H�kf�*���iS���Ã�b���\�� G���k�k���'���v��q Uv��
�u�m���p��id������X4��$��bI��dwo�^��}Hn`(l4v���э�m^�x���4^��F)z�k��O�c �'��~��X)��<w���1��[I�4�g��MPe���*\�D`�F���ޤv�7}�mY�+�%s���s9Ks	퉤��ՙ�7d/UZN���ɴ���.���~��.�Yu��,g+��-c�������(��|怽��{�6I�x��'K	{Y�͑��w��$�x�&qI�Dru�sҽGA����Q^O4|�qͣ>��y�f#k80c��A�ް�����;MX�HW�A	��{��	��ʽ8*K�fƃ�2p]p���ߓpC|Y��C� ��~�ܿ!)O�dB��i���۽��1ꮦ�l5ǸՁ�k^�8�����u�
n�`�c~:9K#h����>�
x(���$�����ת���71]�뗌�8���Ĭj����:Q[�j�Դ�1*}�{qu -��]֠/Y��r�((ݢ;�r��mGpR���ݛN���7^�Y�O��Ҭ�xΓU
���M��d��1��:�榅fy�W�F����!0yJ�
�i\����3�ΜG�=ǴeL̘�#}�ad)s6\<���G��+�d3��%�����A�����qy�@jQ#�s���\��Ȅ���QM\c]<k*& 
�ă����c�k��&e�*�W�L��u>�����q��t�%6e`��F��.=����)�!y��)�2P���+�4Kus=K���� y�e�r~i�P�y�C޶�_댡^J��� ��-Mmnb#�p��8�!��Z���쮲hFׁ���� �G�H;~��Ǹ'��8�6��yu4��Q~�����"]�b�V��dU����r��@��^n"�Gm[�@���������o�jV�D{��]eJ�[�1�{h$c��c�K��ݹu]����������=�X�-5�\jc��GQ��%qFf���]��s�Pο�J���Mcr���V���	*�,2�ZC%# �T[�9�9Q*� �?D�B���扇��;�&@Ykd���X�5p]�M�1D�جS�[�`��(�,\f�Ɨ�|?��H*-�bT����%1���K����|��5ARp�y7�r��A����<i���d�uh�����w-ŗ���(�i˵���p�e>#� M��>[QW�����y{<�(a,k��>|L���� ��-�!�%�c�8z��7ԦE���}Yc�ꑎB�R�%r���x�j�Yc{Q���T���Y�-�Ӝ)��,��p���@�*�Q޵�=6Ia�R����D
����Ʉ2ҁv�P�q]�L(ͣ�)$��k�6ÿ��k���(���}	ap�ĵ�z�Z���)��4ơZ��g��,�V<.<���1+��g�"�-�Yֵ22<���.d'���zt6���7%�:'����c�u�mv�9��F��)^��2k^��k�"�]��U�]I�~��4�rJ/�DZ�&�~¼��N0э(T���w�(_\�A�����CH`j��p�k�3G�?�s\Lb�7=��8�pL�����]�yɃ���r�:�����:y�qZf�z�ӴW�!�Z:����ǇtU��ꖙ��������������+�<�Y�����^)s<���gP1e����Sor������j�Y���þ�yc��M�B4H��%̢����17cwf��Fs�V�2�;e8��"�r
B�|
�%+��X� �iv������XP���APP�9"�{��^���$fI\5���T9�p������^��%��pf�x��UR��$�׫�7�2QȊ��N�dӯ*�*˦b�����jg��A>����Ϊ����1H�SA�\{C�?>�c�^�o�A{7���l���x��q�@��ْ.���JS�7d����J��1���]&4u���,��C<?�҉�y�"=+����Ę斲KI����FW�������Vje���7;��2��i��Il*qH�-ʱ$��s�-5_�躯��/nN|�^ԧl����L�z��?�9Wd c�f.�����m�r775�Z���4p�[�Q~]���Q2���
,�&ۦ�LR�0�&Ӄ�8lط���� ���,�v�����A��K���Y�ڵ�����Y��J���Nv}f��J�x�~/���U�����f�w H�h��oqRO��Sr��v�^�8�j��s '�@�5I;{|�/0X x��m)Rh�!�o���V��p�5]��ƹ9�HǒJY\>>(����@��b���g����X�]�N�'����zph�XGa���9��Z	��G���)iejܪ�h���q<�lyX<�r��ˎ�w�������vXկ�:afw�R �}�F��ZLJl�?f����)��~z�����Ac��+��1
l�[/�-�:��ܲd�S_���_��C���MY/&CV��<e�!i��F�M�^v{K�9lřV�&�@Ja!ꡇ��䑣��?����0��6�G��-;��{���A�� �%]�{���Y�kLIy��WƟ�	��9X�=�ˬn9�Y��ṏ��p�!�Ixnϝ�@��S����T�gC#ș�(�Y�~u}�QJ�Gl��e���ln���I���q�`�\�cN4��P��U����`��ZCe�k2M�]�G�>i�|h��i����T�Y�3��ʸ!	��YG X�D��,Wj&@�����3#�
�b@rcmNH(�z��0R��N�jVM�6U�G/E|�|�x���J���1�ov���i�v0#�kNӍމ�~`�����=F ���訆r��}�Tj�>#���CǾ�~ٽN��Q�]F��?�\�e $w]���d�D[v��{��T,֯_w�As��	[���{:�Ed{>`1�zy�llf�m��ʛ�JZ�J����M �N��:fyu��Bg��7�Z഻S��#�H�Df���c���3��c�}
΢�q>���':��S�Q�����ѣ�C�;�R{�F#`���j�q�Aσ	�y��`��.+�����<�8����<=>3�GС�7X8F~f3�f�3����Aoc�<;�Z��Y��W��#g~������?�5W���r�pů߾8��#a <�_�(	h��H�JS+�fY>�=u���'����8̿�:�7A��,�B�ǫ�I����UFQNc2���]���7�F�dҎH?��ⲗ����{�����0�%���	� 6J��Uc�����V[��x�rI�i�|��ȭ�S�f���FV�j�c�z�\�����i2�'КA�.�5�tjxC��_�%~
5��=!�Aՙot&������t��7c�y�{yΎ/�`V֓��GNK�Ů��-G�4��0nX]���Ħ�x=��O�IKd���{�y��UT�)L�nA9�f��J���%ɸ��qV⛙�,��.5E�|�1��.60K�.�X���s����-��j�9��dHe�dv�tO,M��	��D�������%���������uh�{P�����G�w̆�x���\�K�ן����w�ބ֚�60�`�(�Aխt��k��W��=�3��$��i�՟�����,k0�I�V�͝̊�X�}�2�Q,�UA����\�Fj>����k�� >��7�b��I�Y[��4��׊��}<D��T�%� �pu���D?�T>}�\>~�P�����?��X�v��g0M�Ti�Q����;��׈A��Y����Ȳ�,�ԞʾZ��F���ɘv�i3��lD����0�f��4&JϏK\˻8�����R6^�dk���qk_'�yh�!��B)�w�����O����1p�HEc|Ee��D���y�ωmƂ$
R�� 8��.���l��[T�$-�����o�\Č�:`�XT�.nGy�[�zJ���۫r#��2X��ܟ_U1c�31z��ˎ������]�&�zDݰ��b�m�O.M�Fa��"����i��J�O�4<��rh"�"�	��0�wJ�y��|��	'||a�e�e�_1����{�d�>5t�z~�[\���XcM�����ndi�Pw�fh�M��v���F6� �%��׉�Q��A�C(C1�V_m��qp��p��,A-6��]����cTfݧF��5�i��K�=_>2D���'����UڧO�@�Gdc�w/5��a@�o�0=��R�����f�>8����k��0��ب���Rn,%�l�����{	�Z;�h�]ǔuM�J���>=@��Z��UJ�U���%Fp+G�7�$���!�Sgb9����f��;V��yޫMW�R:��(p2�LM)bXq��;zؐ1�B�9:�=UR���@zJ�!,����sy��t�Cc	�F�Jn���#�/���u��D�_s]Mբ��H������s��n����. ���H����e�^����Zɡ���*�u�!q�i��aᆘ;��޿��"V�x}�៴8����p��)��á}�h���eӇ�tz�~�`{���nZ8�pꃃ9/c�?��m��3\k����y������V��"o��Y���FUQ7>ab�S��glp7����d��)=]�56�i
Co߆%2��j�2�~� �g1E3h�w����LJ���*�0ǭrz>n��`�%����7���O�j�rKp��!��H��x��g�F�(X$E�c5o��r�d ��4��lٴ4n{���dbs<m�|U�=X����#4�)��c͡j�>���=4�z%ؿ�*G�R��������UD�/5(�%?��*�^��N�}cc���R�x��徴�t�k��l=�D�F%َ�'���A�}�.�U�N��bn����X�A]�{ʂ3ep`�� �͚x��?���n���Wh���3�q���T�~�ٻC�窇�zCX-|���pTUM��g]��d㭨�1W��p�i4W��t�7���<6����X���F��.dĞe�q��Y6A�QY4��(�X��ۉ���by�e�kC붧 q�Y~�H��u�vҦõ#�J�/M��q�)%���Ą:˫vVݴ�v�Zl��墮}��1q�h����$�uR�R��%��9�<��ڊ���E&}b�4E��2�V�:����d���0#��p�Feૂe����������ݞ�k�ɺY#��y:����$�F�U�?�ت
ɒ�=_v�>��q�(�� J��1Fk)���y3g��>��O��e�{��_x���^~?DА�3��k�A�(zI ,!�F���7�K|ă���m��L�3m��-��`�����g���dԙ�l��/�%p뚳|*�O�]f�IL;7y���&�鐴`U�`0�Ùl���������oV .:X�fǛ:��ۢ��F���,��B�����T��#� jH�.��$��ق`�h��)k�͜�F֪U>���$�ɦ����+ ����Ui�&��Ȧ�ϊ��Ƴ����[�w��s���ɲ�J��8��fɎSl�mVQ���&�ϴH�"�ŝ`_3g�{j�K���gЙ�0�s�S���R� G�nޕ�%�t��{��0G0zt)�7w�|�hg!FYt��Ӭ�LL�m�5kfY��L�s�>��[���(���R�3H�g�E�D��F�P��ɭ%�,�'1��s�J��w�
���O�YS����ÕRiJV�Mf-E��%���1��pp��������q��ܬ�~��dN�?v�@�Ct���������Z�\�}��((�2�ը�I��H�l|�b�j������Q�k���_S��� 1���׳�cW+�m;�b���aǪKm6��U7p��0iS}� 5�,׻&�u��74X����bS�f��M�(o�0��t�I���â�:�$��,�+o��_�ZL"\OAs��l�a�������Hc�ȅkML+LׇX�+������8�<�uQ���Q�"������֕���#�͐r
C��'�}��a�s�O)�>��D�A�Z4&��q9ˏb�LX��w��Y��C2|o𜸖��q��#;�,\ʽ�T�^�^�% 8���m<yj�>�s³����ޡ���.��[՘�Ds�r\���,7(ӡZZ-Fi/��.�&����y9�fW��hA����ʺm�<��~�Nw�P�����լF�4Y�����:[�1�`�Yo��P�H�s�F#h�Oi���R�{Q�����y��@�
�V*�3diW?�
q���r��*��_�,�ۿ~�Nj4MJ��d_!�e��#�(:��T;�Z�s�f�LwR�m3`_�(��u`�p���m�`���%������G�Ny,owYW_�k%�CV�I����)G"�ɰѸ]�#�BN��^Cj� ߁g��xe�M�Wt��e�'>�\�jFd�M͚��Kl~�=<A��1��M
�~#^.��[Wy�e�s�Yo���U�m4��u�5�E<��CT/�	lbb�$��K�GŠTF���/�ds��ڗ��"h�a51�$�IB&�=X�zJ��+�A�bjk�%y��N�(Ј�%��?�yS��@��{9_�E��f��q��J��U2U��� ;�A���x0��`�\�X�h�ь�d�Uto'U��]y���k��J����FT-�w���ws����:�S6)�bu��p[��g.r��҂ʅ�@��(<d����ώ]`M͟i�Y9��������t�#��o��d���ɨ��~�n_�h;f�!)4/2�m�6�Ng�@>%��A`�5<o�_�g�7j��y�p���s���F��{�a�b���\��:�p��w�c�{��M�bǼ��/�yIE�4Uyfd �\�U?���i;�*h�Mˣ���)�� ��I*d�8x�q��3������u�D�Xk������-��(:��*	ƀDg4nFEc�\ٺ�9��� F����C?РSm��[��1�-����t�5���3�z�y�p�E�-^�*�/�h�|��'��h8�*�	" y�EKZ*���]E3|S3�"ik�{ �9*>X1�fJ�t��!�1ɕs�fVt=�EŜh+,�&�^b�sd^�b6�SB�{��M��ؗ��HYU�fl�M-���:�C�������F�
��"�� I|Ɔ�B�ldб�1\���1G(���<�R�8��2�F+I����8e#4d}Lb��ٗ�ۗn>UA�Ppq&��%n�u��\́�f�GV,���E5���l�X%�>����(���>df�d�8���T�@��1�s-Vl����:�� �4���ý�%�7q�ѽ�x�(%�����y4��4/"VS�.�s��S|��>�|wX1�cP��}���<�@�~�� 43�ib�:�x/��^ơ";�S���@�d&���j���R�ɠ��	���o�<ש�y_Ƽ\�GY�r����Aّ)��4�qݪ��L�.w��E�:8��{g>D���N�pKH���_dA�y��F��9s
�C�Ǹ���דБ�A�b�tHH���]��3u�����������3��$�6}��;i�PlYgx �/�﵎{i�Ӎ�q� �Rl�G��~(�7�\���؝ɼ��{23W�xZ���r��(�Q���1'uQfp���=�,2��-~7�%|���(��\*�=+>H�
�����&�L�cf��AA����p���nFJt��k�$�f�mݸ���~~��y�n*�a°�g0xE��RM�W��t��&3���ڇG�9�k�����yx����0�7񞱠LcX�xX�ɗt�ٟ���/����m`�q�U���02����m�O[����V���v��b���H' �n6��0Lï�� �᳚^��<�}��(19DNs�p�e*=�v�������i��7ǘ$�.1a�[�k�������f>�}V߅>�J����Z #�w��_ޝS��g&(��"�Z8���<�Hi�Φ��A��`F
!BAt8�$z
3����RLWUZ�6 MY�B��3���]м֥R4;�)�vY10�*��u���*�^Ѥд�l�+�ѻ+���m���y���4��2����iL�K��r���v�i�k�>�)q�n�:�2X8�4.jL��&0W��lASX��?_&0EME��k�v�n4����d/�zeײm�}���{��������I�.��Z�B���֛�"d6VnB��Q\;u��؝��=t�-��쭸w��#�1_v������zTu�yM�Tbd	L"�Y�o�5?�qoc�Ƴ����F&)k!cL�^/�X��zt�y�.�!�Ri͌1�D�?�h�8���;�I�pG��E�{�]O�����F�3_כ��CC���Lp�֚��.)G�l���$�o3����%����	��nG'���3S79$����ł�ϭ �~��cnrf�n�x�D������E�}W���#�t�)�k��"��@Q�lY����>�����,�N����A�Ǭ�Y�Ѱ�!�I�\�7VZW5�Az������ׁ��]U�k\�)xw	g).�F.�|A莋_
�6�J��jR;��t�)wd�u t��*��ܠM|�|_\h�8��R��|j���`v�'�dhJX+=+�!E�z||�)��U��i*�P2O$��ƀ���x�� �ΐ��n���4׸K'f�O�V��NQ< *lpkoq��t"�	]޿����������̸1�����N����e��r���i�5j&޻v6F�^�P���D �R�&*I�[$��h�ވ�I�視<�S��hL����3H�`�t�e����UH�p����ƚ��� ��)�JӾ=((�B��vɹ��|������x�ǫ�����9V��*/f< ���_��c��ڊ�y
��M'�2D4J/W�4jP�o�����ڰIzȊ��*�z�z	�ε�2�Ai�k�!m�A}��Z+�?>�zxH��Y(�k���M�a!b���DdYN�0cf���������PN�k�4VD��yW�e�J�jD����>�V�	��.P������Oq����MA`��=�	�O���]��
��A��aP�V��Yɧ n6��[�$�Ts櫭]�"%}��6�ie��G|*�l*�(!cOG��:�囡[�ch�ե4��$�߼(�g�E,��8W���uG.���O��g6�r�y��v�H����x�a�`�>�z{�+�k��3_2��ŋo+�MA��b9�9���H�;��C���9��^�6�S_gqx{-�%�.����|�M�t�P2��J*����Fv�T���3VT�L���I��T;��iP�>�f��=F�Y~�]�QԤ�x����/��WKYt��mnZnТ�� ��12���%���G�����J)E�Y�x�����Ш�5��՘��x
�=��/�8��|��&�h������kI�B���l��u��Ց�.sML*8;��,�:���w[Ȏe��C���3�!� �pU6���7���m2��e�w�KֻR_��i��I53��ն��8p���<>Q�	�|4`z����^����~���&�.����A������zj�z����	�k�B��<	�<e)�����.*N�V�`�΁x���p��9z��ˆ�o�t
����!2�]��P���4��l��6"��(+G6���:��*�#��6�}w�=j����+8�6��7�N�a�2ԕ,����@=�ڝm�����q\�{=Hco�._�M��U5x���m
�Z��}��_ML�,j��A��0{(��`	ʏèk��Sn"g���pl�%�h 3�^�@U�n�ޣw�ۯ�qݲ���!��z�O�|���O��9���[�JhMz~����N���X�'㐂hĊ#b�P�a�iAc��sJ����XaVٲ;�'(��'�Gqm������W�c�
�<*	�*�4�r-��WT:���[���ل]�7pӵk��:��5Pa�:Wʟo�n�<jCJ���Y��w���jS��'6g8��X��۝ܰY�l&/@�M�j�Դ1 �1N�Ǉ�(+��q��3� 1�����:k�\צ�#��m���iH�b�L.�TiZ�sC�F^�F�RWe(�7u=K6炏��+n���b�r�.�B].sd��c3E��y�}o'p46h�G3kZ�㩜��M�R���h���>(o���#�7�]��]�^���ِ����Z��m}:1[0Ab�����sRrz��[�c�e-���X]Ib~\7��٭��#�l�3��+�L����}�qM�P�7S��l0�PXc�����C�$�c�^F�:���$W3����?�!̔m�KŽ��!,�^��� �O?+㮬�'���T�7�uK�E�Nd�&��F�`��`��������Y&E��a���TK���>�tÎ=�
ٓh�`I�Hǿ���G�X��e�Nj1	L�r�F#b<���YK2a���R�ŗ��j����.ЖRR������s�`J���FI��8���5U@|�*��@z����K�.X���0a>т%:��n���v�SQt��z�)�'��eW'��&��8�@j:�Md��h�7�W�!�D�*&��[�<='A�J"��<)D0�ri����!�LM�?O�f9��ݟV->�"��V p�(l���nРM:�2�8��)�(�#'�E��0�XB�H`JP`�����Ǚ�y;Ȟ���{��4ω㽄�t8h�� �"O~sX]2[�ڭ,���ɍlR<�&�&~�3�Šr�k{&L�C�X��JCR�G��Q�5*�q�g�Y%M���(v�!�"+�5�\.iHeF�Oݴlh��ow�^��v�)�	���(�쪷ʘ�Y��E��y�
a��J��$l�@:�3�Œ�YD+ޘPC�l�y�\��,�ܲ�j����L�*X`����������Q0�5�秤.�`�A8 "ǻ���d��J&�Gsn��'wZ�wu��x4Vſ�D-w�ɫ����X�d��ڡ��?�㓴�_��.8�<Ŵ�z�l�9;���.%|��	�X�p�H��\&�:�g��vx��<Kg�#nd��c30�R�.v�t�L�H�K�R\�1{�F�`������"���0āt�ǒ���{GFa���Ecs?�����N�����n�i�����5�'&�ݏ������5�{䝟�Y����l̊)�d	mL�g�[��}ɮ��I��
	��ri��lks`&�?c�=�������{��"��R��}�#�}��U7�A࢘�9F ���4&����q��Ш�K�FG��$����'�6xmX�Y�`��� \�U��Ɯpg�kH{1� �@O��df���`��.#���G�����l���)�M8�A���A+�)I�D�&nʌ��pcSd��;�1c�
�̷�<�N��U[����g�Y��σ�.���ϻ_�Q#�*F��q�!P�M��n؋���|��-6�iM$y�wY@���r<mswu�ƿ���� ��t:s�rMgz��ѝ{p��Kw� k,�/��]�Ez�o�]�4Xr���
\&W�m�`E��c.��N�qΠ�fU�3�q���4맙�Tq�I&�u1,*���RV��Vxy3�`�rw`�E#s��-�hj��xM%��V> ����O0I�������x-��(2"�3un?������X�bg��Z���ԃ��a��Pח 冉��Z#K�rG6�<ΜS$�Mgw&�����l��!��]�Gݟ��=�j��K�G�/*	���k�}R�l���9+6W����ӻz��O<�0N>����6��)`����Rs��.ON4�/A��ǽF��b�WC�x�N�7a�mc!{VN������Y���.3��&�9�?R-��PV��£���=|�JNZ.jd�X���bsyQc�B�fIf���/6�l��ϳ�xT}�Hޞ�rk�hT�Ø�G�G~���M4�EZ}>N
ڕ�HI%3?l|x$R�9H�[����c��4$�(sNj� +w�6d�P؜B�%����]g��E��KG\��!�3ZK�jQ>�ݭn�^�D���P��@0�"���a�"lS�8� �_oȠ^��ڲ���V����y��FD��p�=�v�0�boD����^NA|����Ƽ^nY����tL���XV=��Mì�vm�x����+�W?\���`V�C�d��;��=�	���)���7z��N��Sz�kr�G�%~����i��m�� �uű?��bd�A�oB��p���0����~vӵNq߾y�U<|�E����+d��'�N�J8Goļz㧆��su��:��/���!�oЂ@���d��L�g0g�{(��] 5���Q윭�x�ϧ�*����`�&�(���$ʒy��@���7�F�|�ǿhG 4���<A�i�Yb�?$�����-2U�S��4:e�?��sy���(�@��ж�,��i�͋H�/�m����Yɷ�R4t����e"�%4�x,��1�r"G+h�Z��.L�#u�d�R.`�<鸵�I��(��<v��Q	�)r4D�k��%Cb���Uv�y��4�~�$	�~�-�K@�ۙ���;����ئ4���-���X��B�(9ֻV/�F�Q���<�#����,��FF���)�&4���l��a���We�U�h������h�$��c��_r�ʲV?Lv�۸�X��#G�	�����RH���Yh쿆��(~+y�X�*�(r,=$HG�S_I�/و:�s(�_��v���(��?�Q�	��7p��F؛����_��_˿������?h:�����.>n��--��3(fpDG^��0(T�A\�l�[';C�YsI)������V��@V��5�Y�_��'�J��d���JT��	*x�#��`��&���������X$�m�L�9�o��]��a��Es�(�tZ��*!���es�m�:�Q��#���@�-N�����K���_4�Q��9��X�ӀL2���׽eh� ��2�Sw���R��wc��\]��+̰9KΘٹi�{1�H��,�Z�	Z�mɥC�z8��.�]hg���AgM��I����r����n���B��A��ٞ(������߷��"��K��[\�V�ʺ�ɩ�jc���p�际�D峖�f 6α�r������)��;���f! �����kq8�?��G)ccb� 95GY��5a����)�:	��s|��Ici.��:_��wJ�q�cP��o8
��e���)�xO�o�����R" 9{w80~2aL$@p���r�"�W� f*���U�l�|��޿]~z��&��@�rp~�NG]6J	�`�c�����������?/�kY���ګWo4��T|���.��{M�u+j��n6]7�R���3%��jU^h�{N�v���n��aSi_;VĳL����#m�����`��O�y��}��I�4�5H[|��MVT򃯆P��'����x#TP�����-(�2r�3g��CEo"t��B�c|úLA�Y�[5�uYY���xy��m��
%��m����|w�/��$���E��:@��b�yv6�MVa��1H�Mǎ�U'~/�+�fj#*���)D���4U�jcc��\
��˷�����@�>�u��7[�1t�ew�#MhH3�V�v]�Z��-8n�[��Z	k�F� �	9c<6�m=����2���Q�}���D'}(W0zz�)2�=�:��w^2X�<�Na�i�����D)���bqo^me���NhԬ]P��D�h��M��XS[5 ���Z�{�j;�ߗ��_c�}�C�����/�}-9�G�<<r�*:�`���F#�����ğ�IPI`�:��{6�^?N$�*:Xa���-�_~�u�}��޽����z`C7�n=F�8�z�}��A�܍ʘ����V��%��X�Ț��o�������3�- C��ʰ����⹖�MǪk���q�����2o��\+ºTity��!?J"�7S��3ZsH��f�X6Z�6L��,[�)���I�����8�K�ɲ�$&1�� 6)�v½�V��ӌ���YoY�z#e��rߝ�yT	�aR��:�í����kt ��m�73���$z>����i+޼~^���	��ϐ<�4K�����Ix �M��|t��0a����S�H1qS�$�E�Q�k�������.n��%����ڂhh�g(���yY�sЀ���}�ҟ��o������m9�K��x>���t���M�n�����)��o�x�~�2���O���K߅FԒ&�x���n�g���)�����i�\q�@���@̏������o5̖1�~����C���6������(����so����*��p7����_~�����+9���h���K�I�Y�?Qm�޻�8Q�SE������� ��K�w7P�u�@z����9/�����K�1�h��@f��*=����䙃#��8
�u0�e���W6��]׮�xݗ�s��^��@�4W@oB.��˷���{�ödVW~f��G
"N��jTA��@:O��s�UI�w����Ϙ�R��E9f5Y���^k�74�na�� ��Q.6M婉�c\o�v 	/�Aq��8#%=�-��W��^c�����[wZ�9�"���'f�[0����%��>��l$d����o�7���?M����@zN*���<�OIu�5<0]4����Ag@-2�-9mAb}�C�95�-k��sl�w�^��#!�V�@��?���!����S�}���Oa�Z�~p3<�>p��],��n�׺vKl��rbd�v(-���K|�N�3����[@yS~���(���z��t���v�##}�@ڔ7���m�����QB����wRf�6�����˿�e��������ӑ�>�sd�ӈ��E����c4N~���@e�n���ˉ͋5�i����ś���U�QU��իf��z�chLt�c+!��脪�
��/�v[�NCT%?m�_������#�iD��X �Ϙ~K_<���m��/��P�{:p���<�Ên3p�E=�C EF�eF�@ʾcW��D`	*�N�6*z~X������V���۶6����a�x� �@JX��?�N&u�Yaܶ����Sf�L`���ç�ш�d�a�:��"��~�i[�2n�����f��k�hI�����fP�����(4S.���/����I��^k￫8,���H۽)'�&J�Kz����
�]��6z�=G����l47&�RvdV�]�.O!)tgm���X��JL��s~y.��~���"�SL_T��w�۫�C.�Z����ھ�7����5�[�C�Agz���|�z�r3H����Q<�,ż�F�&�O��!�y�1�<ؤ����Jk���<�S"��̠���m�j�U�bNz-�Zl�]iM.,��wB�8d�(	�>����o�y�=�c�������i�D0LQ�c����:^�����m��0m��8K� Z͛�~��9>½X�IЉ�z�d��a�ulb��N�3�)�	^W:i������W)�N����iZ��֑+��\hd���(�(F�fqǊ5�?gf��γ�IC��NF�0C����X1-���|�"8d?$�=�������}`c�Kiuhp�1f�0{;�NW����=.j�R�.]�Ĉ���&����k�t�5��K�+E��h���N,��Mpu⋳���a���6��?呺�'��h��߲��aG����N��ݰS���Y�96�^�VG|H=U��W	gopT�3�\�J'����*Wp]��,M��Ը�3��3���Wuc	|��9�	W����󘔞1�5��A��g�������`?��l�R�j���k�ej՗գF�� �f��[w����݃�$��P����2g�u����ܵ�)�}ג��nWg5M��Ϡ�l�����B�`�ؤ�)U��f��LFDP\N�����p�o5n���ǪVy�������=m�]�I3�<����ء�R�M��t����W?~���r��P�u�K���p:_�a��f��]���[�"��M13M��9d��T�gL�0�gC��T����?g�flz5"�7
�	ԩ������U�,���>_���n<U�xG�"�z���jJ�FT[�hc�j��R�����Fd�K5����ņd
9�6TI�7-ſQ)�;"����?�'<7��9�{��B���Wq�$�	A�)R���J)��m�K�Q�������j�$��kUI�]͔Guɉ��_lQ� �#�>��L�"TA��bnN�
*iT�.����!�|I��&5����@���� �'�~_���Y�j��ēNH�̣d� F0>`�A=z�i��Jk42�8����ˋ#F�>xTӐc���YV9\�+����o��Y\=CIn�x �C����������h^<2���_�G1�<k%�Ǟ�L��!>�u����|��AR�>+�p��5��ף"���4�e��L��e�ւ[uc���|Lk �x�ׯ_���\�B�ɖ�TΩ��u7���\�M��8���M���������H���ש%+@�Y}x8��l|�p���z�d�����dFO��]\���)5b��Rtq�B��U��b�'�i�
�C����	�h@v��{o�gN0(rs6�=�9{�&3��1Z17�v'��.͈�0������^�s%�{�{V'��>�4s���i����$��r����V��^�]�K`�R[�U
s����<+p��qy��F�|�5�����Z�0E��A���x~��i��l90�:�I� 3��&<|��]3���C/$4����<_scǂ��}���3m:��f�_�>w0�AOI�3o
	%p�i�]��bYY����a�L󒙳-аI���=E����C��ô��e�q�����)��_^�1���M{N7����ks��M#Jl��2����qP�M���\!�<.�|<f�ya���CH��jf����}hB����a�A�����L=�G�꾶���TZ�B�1��"��A��n|F�9S�O@��a�ϵIr�黔sN�C������[a��6�p��Dubl�'�2��ӶN��D"����}!�-%ǌDU5Oym��A��J���X���*٩�3�i4�3�CS}ƚ�����^����t�u��f����ˬ��9��n\
1{\4��/4�F��M�����pS��5�0�Ʃ�3����j(U:gEĢLҋnU�A��1���{�pƆBV�VC`��"�����B'�++��Ў�C��?~������pfj��n�,7�M�<hXN�ѝ=D���51���׃Q%6��m�?>�Դiw���n(��u��g�����z8� ��FD�����^�;��,F;�T�� LàU�5�(��-��r8B��^�9\�il��|�v�@i��5��7^��P���2������9�~v������m�|��8��2X=�ʞ��P��euPxtr4à�[�޸t�Z�Z�qEײ6�o�.�q`b�c4W�T���½9��U��w�fmR?<�X���#_�F[�wm��i�ML����ГCj��dw�-9�P��19����YZZk΋���<��H��Y�;������6�E���m��b��Ҿ�d��ǚ�i�;6��6t��	\����$�e��3�N�4Q^�β���୪w�q%�Pq�.E�3�̼Ff��j��]��K4^�m�Çn[��.H����Q���Y��^wY�:���(������<�!���j�ǅ�/������k�^8�?sb0A� 'Й-�{��)�.�y�E�)u�n������8=���~vL�P@"�,����%,���I�A6x��iH����v�0���E�,~F ݂l���1 Yed�G��)Ue���<�{�`�v4!o���n��!��i�Z��s��:ˣ9x:��Y��X����6 ��J�ƃ�uRd�}'��ܙqxZ���8�T����w$����L���Ȝ!�	�z)bdظ��3TJ�K}�U�	P���mò�Nd���ύ��l��zl�-@������a-G#�H��� ֔�Mc��ʘI/3c>��63�Y�	�n麄
�edc����-���;)��'���>#����=BZ���k�J�c��,���H/��:�#s�r�vl#�@�N:͈�4β�C��5q:R*_42`��vZ�{�B�f,H��8���N�A��ҵGJ�^��0�8IA AY^Y�������E�����lP>�����^,�&��ʝ��wHi��Y����s�!��t��%���O����`��#K�x��l?)"�����ebm8��V��[nv���9>�R�vI������Ꮟ @k�U�n>�Je3B�%c��X)`���e
�f �M���Õ�(lukX�ȶ;n��H[��4����� ��`���3R[c~����Te͚��fR4˔4/�������?`�H���V���>F��ږ����l�q����
�:Q����dBCW�>36V�W�;oA���n%��>끙v�N�2���GŬYM���s��3Ҩ<�hӢ��)� �v�HW� ������O��8i6�ܽ/��f(mj(]�w�}�b��^{��0������n)��PQү����[��<'���z�w���Hu㑐;%��P��$bG���'bVi�- �[���#���_U�]�"���>�{0��%iHwHm�Nr�:Q�23��k?����`���~<9�hɪ����(�	�tS#{?�%���1�0C?�����6)b]�#x$�mg�7N���La���"#
�E�E����[d!qM�����a)`3s�����z�X�`3hfX+��j��13��5�La���zq6j+���1���H��u��t��\O�-'_[#a��oǷq/�:���n�9ع6�%��>{��V��M=Ⓗ�|Ƅ��3V���o�k��~�ؐ����`h��~݉��XҴ�"����B���¦B��u�������x�Z�y�����tHKS#��f,��o�u[;�m�[t�5%�!���߾��I���A�]�i)�X�M����>������6~�U�j��ƙѺ3Fm�t*��� ��q�:�@#���4a8i�9O���.=�i�[�����*CsqCf��%�h4<�a4.x�J7]���&�ϟ5��V�:öV�R;jګ����s�gv�a��z�`	��A*���T3%�^t�'a`si�%���&d�[t�ϗ,�<������&ɤ�=Ǧ����5yKk�ɦ)��Ĭ��dS��,6�R�'�dP"���}`�8����������o�;"���� ��=�"{��ŃfEy}9�y�Z��2����X+iF��#��6{��Y1.��[���l�r�2k䦹�O�+tW���焙օx���i?�r��f"D��I����51�i�����9�oL�.��뗀U��� ���/ |�Q%�T�,�h�tg#�ޜd&&e�|�Ʈc�*�=����ܘkS$Ęӫ��O��v��Q��'Lt�%����IHk��A��}����D��;�S���Hk�]sû�eg��L20���5Uv�p��H��{��$�-6P@I�]x[;+|�2I���'^�\w��
����dt(r(ˤ+���X��7дF�B�ɀq-��9�v��� �52(�<�T��컃��#�6�Y�?�c���=u���"�`��zM5���0�v@ P|�v�ػ3�_��Ee�2d�N?�����U�g�8P�\�H�7�jm|��e����S�����wؔ��]m+igN�Aj�>�Qgv�*������_������P����aݸ=����,��ۿ.�v�&G���f5�YW�V�M;��e��9E/�����-pu4z����%�(�i��~����XO�Lf��:��6��wb��1K�v������C鏃\�����޽����L�*����b|�O�?������NSXz�b=A�R�dʵ�Q��Rlc�������9��9�\��&��Hh���۴jY+=�Ը
���qB'M=�=�k���x:�L|��c���Fxg��:wAtG�7������ԯ��)���^�:z(!��Q�͘c�S]��@{w���3��f~P'���\ߑׯ����hl7�S=I?Dz���.nT�1���31H���!O�jW7Gi�%,����#�{�˼��� ZZ��W�P�_q�8Xf|�y��3�?Gv�q�ɤ�12�1R+%�Ѵ�kHM2#}�F`��WP��x#b;84J����Ÿ�0�Q�������DF�������}�Ph�qPE��]��8��C�l�,��[�I�����/�Z^�Z��FV�U޷�J���Y�� �ݷp����Ru���4���v���-��{7Cl����C�+�t�)�xNg�lz�*'=�`�g�?}I���0㰬��K6KuK��1�l�n�W�,�0Y-r�{�~�f�>o�Ћk������B�L��2��7=�HϚE�Lt�d�9|`��P��+b�]2mj�f�C�cN��#	�N}���\*~)�1�<z�V�<�F0M�V�sF�a/w��{e��˺�F��t��SҠ�E��%����5B���&��$��+K�QR��*�����=`8�H���&�%�"�������u���n7'0��B��vh�������WX�9���ȑ'_s̱o6���/P��v+6X�;,Z� �g��孊��y�=7�����Qp�i�귺['���9�I��m�ֳ���;���!' ��A0���F��_!� Z�[K��S�~���/a�ۅ�}���~���,����ʓ�Ԫ�-*>�As�a ��������ޜku7`�����gr�����Z����qݘs�a@}�n5MM6f9�cm�σ���l�����*�#����ܰ�D	������P����S�LUς)�L���^�5���ʊ7��[e��He�m�ihHҧ��>��}}N��k�15w�~�d�7��p\���Qjj�%��{��P�t��Q�P=�ȱ9V'���M����4�C�9͛&V���"�I<���z������u�����k��8��#�ҊL��v��C��l�G��x�sZ�B����@���x�%�OG��W:��u9�z��BU삇���u���@fX_�9�酓�\����.�6�<U2n�y�"C�شȀPb�$'<���]ޘ"� 8��ec���������ߙ��Nq�id]��\5���͡��ղl��q���^b3��$��Y��Rw��EC�S��7(�b=�z��uMI51���;�ͧ�W�0b�V��g�,�z����0���,A����C���<�dV��\(�>|�������u%�vpŖ(�L��ӈn�&�F?L�����~/�l�~%�i��Аk�x�#)a�r�rȃkq��b�{�'��k3������C��j'L�6o1Ew�M4w2L�	��� ���hnĕ	�R�!R��B��f�a����D��^��qT!�(n���(�/\�5��1)@���.�5	��1�/�:]BYg�Ȩn��@��l�!R���ՐG��L��ݥ�H�d����z��=�. X-�*Ӝ1���x/�t��d��͈SZ����Y���|δ�3p��8��#.�\J�*eUK%���-��qd�()�a}��̚�L:�E?�H���I^��a�7�'}O)��d���iR�Tf�z��͈�BN�c�;�F���?���
���1	���2�%sμE���>G��,%���f�L�ˋj`{^�)��{<���xDW��-2�e�xxq�e������Ǻ��i��Lь�C<̍�cY��և��M�k�����b�8��w�ky�X+��hd�F�s:�}=�J��ԅ�?;��P�1k�-���~���{����V%��_���#pd��7y�j^Z�6����D��qih^�J-YyCދ��g� \/l�NI�µX`{ JyzE<�x*�TJ;ՙG��kC��+���ԜS!ƒڊ@�Ϙ��1<������C���1�7d�hV�*�ką�MԸ�k��%/��ן��j���>#-y!҉f���x�"��k��� �NBq�J�
�QF̤���ZeR�d��"iX��j�̡X�?�B� m#W�^��&p]�X�wV�6Nl�8��C_g)-��-K���Afㆰ/{~�A�����0� 7/�)c�-�ʮ,62)4�jg}��}v�1��WHro����,�׸w������<׸+�����鐝�#����i�;݊�ʱ$��/�Gl�qS*�Ld���r�N�6�b�?��n���B�3�%�˯����r���}���D4��@�'M�r����VU�F�D0:�˚��I#�#(Tä��Kn����f|tM�;�[��[��x���+]����?�����~� �7G!7Ɏ�iБ�P[*������WI��'A��sϫ�v60��=,�u���>�S�+a�j
*����a�vŬK��:�I�e����,�[�CW�O"��8y��Y��@�g��^�4����5���Д�
��!���Z�'&�ݬ�:�8^����ܿ�]����A������{*"�*��$����ˉ%�G����+��!��lz��녃x&�A���/��z	x!M�j.��6���JN�18r7�� �.��$����ٸ\cu�Y�Űr&}t_ů������(��:M���Hhd{�# �t���-� ����-�5�#^���9��2���7N~hpHoH����==kP��>���pP!2!����8��Q̮�4��;�C���X�z�3��`�����[�fѡ��cV�Tp�a��\�1�T,��Q"�Q������M�n��������m��;�d[ra�N�������3.�������͟x�at� ��V�R�VR���*~z<�q2g@�!���~^ ��z{YF�:�mz���Kpzeds�w4���>�1,��>,v�Zv|�]0�7Ŀ�j�&�����'7�ڦZd�zB����0锜w��2[�]�n4�4>�g�;��N�Pu҅7}�wRυMao�ƀX������c/ը^U=���_������&)�D�C9:���ֽg����Ɔ؁g��#4�-�uB{5v��+���!G�DY"��1�F�i��P���r�۾�Ħ4�]6Y�;������N�Ğ��*$����3J�5��Sx��~��(��c�^gN����l���[�ء5����������υ��^�;����⠒J���5
�UB�d������{uӬ��nm��/��hM��d�l�ֵ[�C�a�AqV��I΄�����yǔx��U����;�zF��ό9H�j�����z�>���������F3g35�Tr`���C��^_ϊ`���&��I�kCI���Y����-��ki*�ɞ��]��>g�M��6�c�`��V:�.yHuR[F�ܶ)3�x��{�>`�W�_?�$�+p�]����#NkPJ�V{L̶f��~���l��z_��
6 �A���\Ԏ����J��g��h��t�_��.7�8>N�r\##�A��4S�H"�Z�E�ĿXwfn
W�#5��(�K���Q�t�����ڛ��63S����l�,p��BVw�5Y�y�?ϻAn��A�\d�X;��-���*j �#�8���h}{||�S�QY[�_V�g�2|u�W����3ز#\��0
j8�i��{3i�6i"8o���8�Х��\��F5:�Į�����2�tz����1k��͢�V��xt�\Z�4�HOT�q�Fj��{@EK�W��i�V��=m_�8�no�|l.h�9�V�������pA#>���(c�L\Ψ��&�U�}��C+�N{_UU�=�����8F��Z`xI1�0�p+A,��;�I�2]�P�6��7	�9pV/XO�e��d/& ����բ�]�қ�!���zP�����0jG���mL*Ⱥ���dm�/ ��fV����8��F�l�t�k��G�XxZ|�^�����J�nr�)8}��k���Y�X5���-�{H��t����3� ���N��|�I6G���;8���b-A�Z��$52��x)Q-I\e~cc�daFmG��Q��R�*1����F���}t�=�oV&u+����LR@T�ڬƣU~ �Kڲ�0WA��]�e<N�D)��
u�:���I���|"n�Z�4�����=E��2�b6�\^  �[%�}%�;X�I��e�+�sx#��9d�o�8�PUq$L="��_>�l;H9���D��ob\�LOE~��%Tt�t�b;�а��	�'�����$������~Şϻ���O���`b<��VZC����hj$*�r�X=P�c���/����K�r��ʿ}�a�8�0�n�<�@��;�9콹9�m\��l�&8c��HVM�e:W�h�5Č�P۝�M���{�����"�wi�C@-:q�%kt���Nt#�N,wB���|��:�D>�������'�=�$K�$1$"2�XW5�r��;|  ��?�Nng���Y�d�����{d�άr6���2���nn���Z:��ٔo�d$��-�R�kz~5/CD����c�B�����T���Y�s��Wwp�@��8�	�A
�hRr)1V�V�����&�>��|,t��4%�^R����
��VM��� ��[F9��=�A�3�#�ͭE�}6Ʋ�8J���V{bun*FOp�q��TG^WȊ�mQ�a,Ȯ�1�d�\a���ZT�2[!��Ї�����9߾5�M*���1���cR8`�|�*|����*���b��3��s7�c����J~=϶�a��uU6_�!5��V9Gqu#�R��u5ӥ�+D@f���)	�)CW���2�"��IK��b���߷��]$��hҦlq�I�(5|i�Ä�+���J����QL�!a���/�CUd�
3�z�0�����0�
��B~��M����CH'w{Q�z����������7�.�%~����?�̽��+X/Q��ǵ�,39��Ob�<C��Xl�����陑
�g��)ͅ?��.%���fQF^w2�z���._N�o�����!����Ϸ��26��E��2�.��^ #�>�7��{��h׿��m�>�%<;��$B�4�l�puAn;��Q2������3ǂ�G��
,*:��XD8���C�j^հ���2d<�%���u ���U�����5�@��#Ow/���U)�� �q�>�v�N1,���Dխ]26 ��j�V�>� ��vmq��$J���}�;���<ff`�'���`{�,�i�5�
uV����U�v�<aD��ߞE�@�on��)b��F|��ny���y�}���k����/�R�Iה�TI.���s��S��w1�n3!��\4�F�c</��0W���GR����5�!���+�5%�����3��A���A�mf^��3�u�C���'1S&A��,k��:P2���F���7q�e@yV8��.u�K��]f�E���S1�)���OmF���5�67+�,l��c�`���2K��)R�gm6)����t�R���1��zqH}�{�%`l�Ab��DK��>ŔgQ&R\E�T����u�"�4K;*�?{u�X+�f"���˵p�2�Ah�����R4�4����(>n���!�� myb_��(%��W�v��uv�Đ��j״+°����$�C�X�U�M���ʹ��ar�*M
v����E����oʗ_}U����f"!�����Kcf������t�2�X��3�g�A��].6ǪER�|�{�[i>~.T��t�e�ud���ͷ�w1�Ry��TBõ?+�DpO�w�j��=�Z���Xr�!	��,�oe�T��7�1נ頱�e�i�~AS�kf���4Y[��셰z����ɘ��ʲWң��4�6�3�<�wr��}��_I՟VѸ'v;�:�CI�ڽ�b١�Y�>3R�\`�
$�]'O�Pm�\/1�6���\"(��P�T`����h>0X�t}�cr�D|I[yf�S.�i`?�n�!�N�۬�ﲴ*���O�1��Q����k�R���g����]��t�W�LN�� 6U��HTDv�k#��_�����
E�U�+��%����1�Hky�j���3��mR�w�Tα���}쎕
���42G�#����i{��1�c�XV�w]�Fd�z�����)hR�ؘ\�ѹ�Pp�6��@dC��?�<H�_~��p�.�'�`�lh���.���6f�����rCo������ ��,�r�]���'��^�q-���(���:{/1>8�j'��KEN�<��^�/.��Fp�ȫ��E �I@�p����&�"��b�
�4S���e����i�{��WG��iF���?��RD�/�b����3@�ˮ����zftrk;����EU\���ILZ�(�)n�5.ɟ(�?��`���t	��Q��j6�@#��Pu)��W��bJ�*�ոp�x{�nB5�c��[���6�3J��8�����esg�AtI~f�g��R�g�����$�E��}ۋ��2<)������Nn��_Ӕ�e�:5^Gi�h��C>"�ɱC0���!(|��Z�
�*�J���]Փ>`� l�zaQiة�!c�s�#����eá��)�㺤GLN��U ��r٥��h�Y��c�
T��_ �~�eS��'�ܝN�����Y��s�c-V��}]'}�1�e�K2��Px���ShA��鮀@�&&���cb��H����F+o��@�Z�>���^���^��w����(�4O?�r �Y=|�Pt���Iy���`:�@,��� 0Zx?A���HS� B�<�X�do��T��@Rr��t��l�@��1��P��Ϻ��)����>��a����>���2�����賙U�\�}���^��m���?�M��	�ҮN�[��n%V��J�馕�7�J3.����ԤL����Q�����F	6���	��W9^����a�9N$����T~ `A"|>)1E��@��X��$�!;��4?$	��]d9�%}�}=��^�@VR���1I���1�Z�Q����<��#���|C!8�����p ��)���y��dJ����D�a�'��SG>�"�$ ��Z�P�r�Za��'IJ\�_}�uy���?6���(Rr��nxP�T���Dd�] )�HG}G��:!��k���4��W� 3�E&q�C�Al��i�vb�̂0��$���#uW�'U
�����^�d�Oܲ�N���8T�b|��wܿ��ǐW��K:���գ��)�+3�]�W�N� J��B� Ho��5�#��X�H�T��pS��ٳ�K'�`e"������]%ܻZsu[㝼��KWW7���j����G�Χ������SoI̒|�zc���'Ƙ�z��}<R5>�m�3�?7��wv�Jxٳ$%͈"�3F3d���0S..���6(����H�FJLż��i�]�vĄ�}��j��OC�G�6���W�6��U��=`��c�-���$-�^�S(�������I��z��Sb����7&EۊظVu4��J$,�(�d��	���Z��5�Ȯ������6���R�~��uh޼y]����}�P�g⣲�� �!e.�]qI_��8�ҟ���%戓�JUW�釡��la1���"��\��)鯂Z�{B^.($���ߙ�EtV�n^i�ٸ�iX��i�s�1{�ݻ�K�=��f[��a��݉��2��4WQ�vc�|:'t�����F��Yȗ�$�A�g��lpkۙۃ
�O:ݖ��/>dYZ���c%�fs�Iy̞�O0E�р����db5J�����Uoƒ}�j�S]3Nv����$��I��{\��mZP+o�{�IU�gNC`E�y~/y���HP�e����`�1nܜ���t���w����~���3���b������ǜ
��)'��t:j�}]�ᦅU�,�k�~���n���  Y�$��UM� W�pgp��e��"1L6��@?3�DJ�Bl���la`��8QW�k�-�r\��.�.rd�]:�Ϛ~��1gy���_|Y���?�?��O�Tr3(U��%0��\q��&Z�p�օ����C�h����a�I�dp"�۵��U�����V��5�n)�գ��3�k������Tum��8~}�7�T*<��g�fF����dS�f߮��F;�p�Qѫd��t��l�D���Pzᒻݒ� y���fե{p�
�n�X���J�2ةՍ٪�asMR�Xq].&洷�	��6�R�X��t:�����4��t��}ڀ�C��,Hc#͟�H皑*史8?춱�}r���',6B$��,'�lD�v7uЇ�mt��|
���Sf�P��v���e������b��/>�r��w��%�����sp�t�r�n��_6���!p���5	/r��0�V���[���}8>^ܤ��L����M/���#1>w��Ƶ6�9'�<gl(����(�\���M������f��t>p�����++��É���v���G���e�/�b �o���M�ԴZE��JNnН�Ì��d^J��g���;7F����d!���J��`�� s��K�y��Խ�58hڪ�Dq�555
�tg�p�%�L!��(�1T�� �� ���9��%v潦�d5��>�2 ق��x���y��=	�
]�zt��I�S&�~5�P_���{�6T���k�7&����CO���3�,Ϯ�^��PQ�8ϱ��(�d��CN#d�h.��)���(a�s�����ݭ��a��ګt�}R�g!�$���:w��RiF�q��NJA�ٶ���:��+&%��͖:�kl�7b�����T�o��5;YS�ҍ7dor�,�� x� �]<�����z�d7W�L4�ʪ��vP����C��t��
ݶ\5���R�����w
�AX� ;+��>����X�*�Q�d1[L�"������`yˡ�(�>Kc �E`�>���Gy����F(�o��_~�e���Ct��d2�r����Z89Ǚ��Z��'��˂��o���&�M)]�Ъm�:щ֚qF��B��YdUx>������Kz���=��(�l��)�#V�ڭ�b�I���"��`��LG�Ԁ� Z�Eާ�tUF�1]s%�,�{�U����c�b�@7�?���}7\f��R���*/�#�]
�X̥���ZE�<�X(�b�\�Sƥ%0}�����;U���!�;fN'�v&��|�����ϧ_c�'_��T��ʵ} vI��Xfv������.��D���/p!�� ���x7��5���oI�o�wڬ⡜P���B �%I�[m(!��4Y`�����Ƨ:N���A�6HD���:�Yf��i,�Hb�S7�q݃l��61�;�Dn�#�J�ɫ0O�r(��l@
���	c�^L�,����:��ˑYd�n���w�Cd��}������hP���"�qTBȈN}~�s�9���X��P��n8ĵ��k�����p7w���%;�Y��ӎ*��Щ�� ��/��u���(�LA�F6�ݐ�7JI��#��������U2GSe<^σ+�Ę
(�-�[��y����v���Yڡ6L����x� ��`腁Q��M)9^�Q6��~UE�#�E��R3��Ś�#�� T�b|����>�]f�����R�xiYK&O�x6*�w/�6j^6�ڿ�w�i -Z\n$�x��?���c7�"�i����p�&�H_���fѤ��ؕ�-g).�[a����˙<�H}�ścS�
���Ac^2jL�zB���*lL
�:�p��3P3o���>p���o�^{�Sӕ�q4�J�X`5X�
��(�p��L�&;
6Qg~V#/ؔ���.�R�&��i_���iX���]|�8|� !��Bbd�. '�j_n���7[����X���������F�e�����V����+|�;V�Zx�w�������~r��Y��rM����t���I�]í�˛����߽�o)(g���pEљȼ�U�=p���Jc�e1)@�Ɂ.�kd龜q}�y�/l�̟�ا��Y�I@�,��q�s:(8[�dW[jv.�=���sb���?�X;sD�6���0��Z�o/��I��B�Xjѡ�l�V̲�j6�/���a������:-U��x���~WZ!�� ��K��fZ���������_|i�`�^"2QFw_�q����.��i/����t'��`-��`�c���g��Ѓ��E]=�j��z��KN M�����cu�c��S�T�l�>U�}"����#���x��!H��,K2^
Q*�8�#�M���1cJK�15�������#���y�0���bk�<���dU62I��uh#�%�:���>�����TW��88�8��|��|�����o�)���-+e��.��b�t'=Җf���ϣ�Og�47<R,F�LuS������ˬ�,'`���';K�Q��B''��Fq�l�-� W��������]�(��^!���X��KU�ծ8+�#�&M�9!p&�{vZ9wn���!nP%�ǞX�=�c�h`w(5a�#lU&�$-��0W���8y�J�t�$W�Άw�)�z��:��ý\'���W�UP�ɫU�}c��9�yD���覥��P������i@힆�� �Ͽh5���."�%��O�2zi���.���w�4x֤Ƒ��6��60d�l <$Ԧ5q!kS. �g`>��m"�M��lw��5?��շz��9u�N[���6{,��:Q4��+=e8�h�J;����E�q'�D��1��q�>(H��ӡ����2;M"��Y�8zӒ��DVv�7ؚ���X�ꏸZ@P�Jtj������W�/�,_��H���#��lo��X(�}8e��'9Z��M�e�����Xh]�V\b��5���5�+=��@y}E��gG\3>���N�Tv�#�-�����N)�7.�"��de�w,K�JO�o�����/���['�����V��A���-4⢍�f�52��0	�\�������L}�OZP�n���V46� �1�eQ�}Ⱦ��ȠI؅:Ʀ���u<o����d�p�oVezd#
�Q�k��>a-6*���+�{�Z��e@-������I6{�D� � ً������]k�fr�SŌ�3>�� �5&���o\��=�Qr�{��Y�.�L�o9_%ݖ=l�:n>��P"G�D�nܨ��	������H�8f��kh�~�)V!x;��+�vj(�B.>�3*��!Q�J��}�4�F.d�M����o�ʼ��t�Bz�����������ge�T/�H�����eL&}��oが�����&r��h���J>b�R�Q�I��#X�%��	ZWBL5k1¥~� �g|ཪ�ws�&ɵ��xU^��yL9�M��3a��ͷ�ˀ5��6��<8h�bnqN�lȞa��e�o߽�.�?���H�;4	�:i�Ƹ\����]�A`]=�.������(�h�.�`�Ǟ�>0�R���k5ՌqY2�ζپ��E?1N����-Gpc�e��Y
�s�>�zxo�ў,�m���8�{v�����9���:^�$�^�Y�
�m��$��K����0%�7J>8�G�f���_�72��aB�0>Q����)��Z��ΰ	ئ��*�q�Ş%pB�*6EH�o�qh��@?*0/�'~H����>���b�	1���r�H���r27~_�/b�D�����C�q��K�l@} �`��k'�6�OĵL/�~����Y��f1Q�C���B�j��{̝��Ed��~�m�/�KR��p�׃�w��x܆�2�un�J�?H�"�In��r%%�:g3d	�NQ�u�.����GM0am2#�TȜ�D:��^U �'���9,�HƉ�ב��),d���Ͻ������~��
�T��������;	9����C�Uc�&��;������b�V�������3o���DՓ	�jRЀ-�0���{h
l��W�Y������/��]K�����ۺ��J���^=4��Ÿ�I�ԈFs�]�j���3K���灔�88�q�r�2E�L�v�a�ՓT�̳��!}��6�dŬD�&k��䚷�Ժ*F0Q�/�p6MS-�"��{<��av�n�!&DzbNv+�f�y��:��/;����Jw��Eb�KJ���d�8�0��|�m������w���i��^k�+!p�:lg�Ц�T:-FJ5L�'�rlF�8^���'y��)��s�gqo ����#��S�3)Ll�yD��c`�h�{� � �&�\g}vO����ʔi݅UG`�UZ��뗋��� VQo��cε��1P�n��g�s' 	�'�L z�f�9x�&l�,�}��e����{�D=�_��iw��"�7lJ�H�=f�6��'�$��W�#�"�A�C{�*�Ҍ+�+��4ߙ�ui=��W�?kO�f��@ox�� &`5Nu]�-zUN����6걓��;�Z��^i'���e^�f��P�eD�'�Ԙ���[	���l�G��#�eǌ�s��dɸ� Ύ"6p�l���Ml�lH�FT/��|�X\�sl\|������Ѱ	_�+5%f)�ω��w�(B7Qe&�*��9��43�����J�Hjj�n7ʚ���q�Vå3��97%(���jZ�Օ(��H'�5��(,�kS"!Ԛ���,Ia;1�ƴ��i8RT�XU�����1'��W_Ei��3	)gٮN8�����n��`��(�þ��j��f�F����饨Jxɜ1��]�1��6���D����d)���������>�� 'R\'��P�Qk�?���=�� l��O?m��?"�����/��x��V�7џ����s���}W�pks�������5̜<3HUq�>3��Kb�e''�Eb ܃{x�B���W�yj(f��x5�Di���ke���������>�	�Á���0Ǌwנ�O�~��TN|~��jgtL]��eT��@����@ʧ�ԏr��ޤ}}ĩ{:�EFc&|�����b玞I���<�v��1�����1��n��+�n�<z-4O/����x�'��K��\ѿi��zՌn+�� �N~�Zdhp���e(�E#:o����i���򔿍������J�� �$�[nrQg�1���T.f�Cv�9#-�(�P�&�����>pb�2��G���������W_�"�-RDQ�#y�75VZ�u7�vR�w���n�aټ+� X>S��T;vd=���>Cq���	�f�rs*nYYF�/����Q�w�u��s��ױ��P�X'���w�`�������DE@���\8�`M��,�df��<����f�x�b\�u������ ��/Q�@�p�����z ϢҘ罻��{mHJB|Ʊ"�Z���Y"	�$�N);�hLo�-�)v�X�j��^����5�aX)\�8]xyP\6��D����7�&(��'�3��9y�TJN�SZ��+gZ"���El;dO�R��V�.:�A[��;C�DXȸcp.]���s�h 5d�s�X�.Iڴ��wv��M��l��qJh� cb1XX�������IE@8��.3X�ۄ�5T�e�p���}ƙ�}Z<ur{�^��U�x�?�}�0�s��X�HX�gN�`@��C���u4���6��/o)k=�	 ?޾{��CfC��+ )Ȟ�+�+o6C(�n,�[e�l�)�-�b��Y�4bcv�F-�_�Y��5G�����	3c��f�� ��?��K�e;P���6�d��pܴ���>`5O�=�cvW�actUF������$�2���k��/�IЍ�R�=k��	U��b�>�Q�OVIS�ꈷ����z0e囈d��<{�����1u#�����Y�������{͇���<������D�����_W5.#�����k�i0��cvi����Gc�C�5���:�x�UŅ`G�����9/:;�Ke ��MЏ\��TK�dL���8nx�����5ʗ���ZO����~t�ƀT�����_��x�5kX9N2�a����<��)�րot��'RJ��£�������@\�P��dH�^A�Axɉ<h�A�c*��i�@�Zt6I�;�E���\�cˮt玴)2�י�>���*�s��]
��9`8�U(��!G(}�����Ҡ(�̝�\�u��*d]�@αF��?��c������-+���^�4.M�<���g��?�e(|�Ӊ	Fe4l���:��}��[\PZ�����N[��M�&��9�Ιz6�p�pm"�H���F�����{��m�ջ̦s5� `9���e��೸���/ۨpW8m	B�ìTR�*������68����k�S�Q	5���k������L���h�!�\CZI���2,# ��Œ>ݱ����9��f�Y�:N~x��׻�2'����!�+p�@�!ށ�j�� �}�O�g�I��>�Ն�N"J�[����z��{۞��jt�/�UyM��G��~�"���1��N�����X;�����h]p�ʘ�g�U4SR�<CH���N҅���,���3i��%�R`1 �$���M"�Ɛ�K>|��>i8����ߘ�;�'����*%[�* �҇x�9�}�#]����z��2�3É�P� ��؈$�)U'�+pA��i=M�G\���;�2�N�a��Y`���O����e���E�F��|s1��.���7����B�e㎸+��1�����i{0\l�3��������hx͕,�@�u]�������/_�d��&���:����9I�ґY������a��Y!#8Q`d�ޓ��@��I�r�ќsF��R�k����EpmΨHk0��uU��"�6�4�I	�#t:#�*724tn߽���77Cv���1��	0ɔEF
Z̐�Q��5K�;�"#����iv��(���"#�e�$��I ���q�C��6+2�/>�"v=������b!E�&�[]�	�}�b��/����|�͗A{y��m8:bA}��Eཻ���z˓JM�L�9�`"#b�O[�q�,1���)u��������\�S��v�M̩���r��H���Ў��Rͥ��gB ��N&w�!��;�q7�B�(�qH�w�c�v$��c�,�5���o�)�|�m<§�l-�s���������G�@��^�%YjC~�+�d'�UpH�8 Y�<��8X(�� �pO��\�����%^��l~���o񖀓����D��=�e��Y[��MS���>�d�Q5���|NfμL�;�&��-��~�_AISƏ�#H�1Xq��E�ac�������%�|�x�c2)�:�7�Pz�\=<��ڍ����dŌ15�>qѧ��E��ׁ��������M�L�s���R��%7}M�;��A����j�n�^a��'F�"G�]�>QLt�W�e)�Ow��%��;��q3� �6sBE�X[e'<4���U⺌�>�i�6�Ȕ��9��3�P��(2(��hT@�~;X�&5�A�oS��H4t�S�R6*���&r%�^($BE*ro��/��j���;	�~'A�6�dL%�;�Lc���.��v9�)����DWׄhd.�ǝ���Cy�&���܅���A����8�8���,	����W]3oؠ�a�3l=�%d����Ę�-6��|ƴ��3N�	qݐ \؝��y�=�"C�����%n��QǺfv���Q�/k̳���3Ձ�#F���e׃ʊ� �dc�Ɇ^*���c��.1�[yM�0�]�]S�;tSwH���h���^B�pC�J%68	���ۀl�l8�:�ٍD"��b��r���խP�����x�/y��'��40���Uj][�S��h+*�z;�c�]��q2�$C�(7*��i�e��yJoo�$��]f�Vw
���f8O�{�/�&V}�%$ �)	'	�P�v>oA.2?����@L?K�<Kx�����6*�aO^���c�m�=%��(��6�����@�Rѡ'9�U�a<�gM>�0�U��a�I�Mς%���>,���D�w�G��DؙkԴ�|�����$ �g=Ŷ���1f���yC���4ixU���C����۳�����l-��
ݛ��t!hp�P;����_�ں"�B�K^��*#p�����*���P2�����>��/# ����cв7] ��d���{_X��@�Ή��O��N}�IJYUSw栆Dw|Y���W�К$�~��\8F��'ڤ,ܙt8
\��e5��$����z�����;&A�*q�8�� �Em��qφ����X=�;&#��y���E ��X���M�&vmm���7�i �i���)y�R�(li=��uɓ�4� �����MR�	n�jY�^O�^=��,��LA�R�"�g�E���wB2R�0��y�ir��5OF��wZ8(7V�����2O�YI�����):�;np�����Mx������$%��Qn����L�:GYW����ӹ�ٝ,W,\���Q_m�84�P���C�	�,���M�RK�%2R9����m�RǸ�mpFQ���h� ��-�e(*}��7D*ቩ�� 9���*��{���q�{Rs�q�������V8aW!,�$���⻾y�yr(��#p��᧟&�`�;0����a ��{`&���Q�S@���$z�j�[�2t�bϨu������:%�m=ȆI=�'	��|�a�5v$��kg<�d�q����\<G`�A��ljH�Ӻ��Hs���I����D{���5�k���P�'��C��Ω]O#B�{����]��[h�hئ����'a���8}�I��i�H�t�bS`Nк�^�(�M˱
O!f��C���a�T]��`�/	���<�T�oŋ#@�x�d�����>Ep�N��:�u�cy�����Y�|��R�*Kf�.��W���!��e`���w��p���� ��#2��^�[�g��,�ҀjΚZٍ��0��Ԟ��x�EG{-�Y��6���*w!�KK���f�����e�e��#����ct�Ew�ꡌ��a��PX���������If�1�/��ux\�k��	6���i��L�SU�"�(�r��-Cf�ʇ"�!�h������Hh��K󮛳B;K��a|��%'Q��\Y�CJ���&5����ʖ���;�p�y,��r���s�a:h8��N���E�ǆs��I�3n��p���.�gi�I-cW�N�Fp�M5Z�w�q�:��б��Z*?����^�{�{m�,���|�6#5��%�>��ul�"�v�N__�OE[e�����/�*�e,�������US�CŧS��6�ZK�T���/�!D�8��6�s��Nc��������e�!zB5��6ے%l,��T���q��,Y{��yW�M���+�4��rf,S�N�@������-)B�Px'=
��Z�9B���,ߘ�x+��[j�&�^��O�d]��ԯ�D��È��,'�h��Ӂ�C�z��p���xĕ���@���8�u��a�,=�,�ӽ�K��޼��u@�u����	����+	���-�Z���s�t�Տ�6��fS�e@���ﶬyˊ�����T\O��������q��޲$f��;( ��Y�JW��gk�����f~?|��t�5/5�hK%���p+= 5L�LLѠ6
���CY4�y7�?|��ho�X��^u���g��;[���2W���y|��O��oj�	��3E�� ��܃���[]�-V;g�p��;@ਦ�Ms�r2�.5��6��-U�OVY/C��@�]�Z�S FMXx��~'>]i����>��fe�&K���%��OC�nM���
�{�w' ���{��+��Xl.
/\���h�*U��@36GX��s^�1$��9�˴�����TeG�4�:�G�����ɻ-(�����n�}�GȂl�� �e�r{�.!p�}����0��Ha���`,:��ļ6>���%�v�&��&��b-�l(�Ӄ��I�+i��>)Ox�W[���5(J����D�Qd�Z{��(�����3l�����m\/t�����?~_ d��^�d$�W��!�6[v�kA�c���u�~4��n�n"����˯?She�8԰��q��A2��M�Q�|3��'�ظe�V�p�0ƺHD=��Γ��NZ��\�Ǩ����2��;��ǟq�$��pv�tS�j���jcٖ-\���b����t�<�:O��� �﷝�:&���U������慻9�Yk/"���A��G�O�������4�,��#�N<e�z��{�"�6�@ו�_�����T��T(
��i�?𪕸��,/�S���^.(\|4d,sM��yɌ�N�}�$�(Ё��n��o�S�L�?;�I�QG��'5nŋD�����\����P���R
��v;�����Y��s�T���n�x�F1b	�bd�_n~��WQ�Y����Y``�<�z����%*��Q��>�p�0xZx���>�|�����I���������c4��e���"�˟�����x6����θh��k���/�Ͽ�T~�������=�>����qm`��|�l10��5O�|زU�L�T�}e����W�A����57*���?������~�É%`��!�3|P۠B>W������3���٨&��"ړ���%����)�g쿸0R� ����4"F%��x��`�A��Iך���j8�,T����YL�NE�f�h�TI
��8D�ݥ��m�uEw�laPҖc~n7֘���Gkr�0��j��郒��L�ڮ��M]��?�G�@�}��wf�Q������3���2��i<P�>ޘ]=U֪uh/�*X�V�Sg"12�FJLt0��󒁗�W,�/�@�<ʼظ�/kH�m
A���%QB�U<w�h�%,9٥��C�Jg4��&=�P�������;��3�.OϮ��x����2Kټ'���T�  H�x��&���$�?�U o�C&l5�I�|���_|�Edh_m���_}8(7������dG��V0]�9uЧz6�`���m��~��ϣY����+������.\xǀ(pq8aF�6�pJ��!�,�SY���Ѕ����i�j)f�w{?*�A8(�4��xOyu6ga�3E\�q�UǬ��UQ�)�|�QT����B��v�i]�OaQ��R�b�N{�V����7V��U����
�k!�����~1`�=��AՕ�G�'�S�ޢI{Q���ā���d��>��şMݮ��_�������7Q7LK�l8�Y&6ǩ��P�]]GV����!H׀�8�|]8*׎�q����-�~&���S���ʊW��(;䃤�(.AN��{�r�g��b9��:�3!�<2�k�Eh����h.���,�� ȗ��D*��޽6�����c4���a,�����(�d�Q�5��KW��km�š��C̸:��4A4�~(3�C��^_�y� ��@I����/� ��쀋Ҏ�U|���B���wo# _p9�\2o�nd�����L���Q����c����s�1�9��;�3�-뒐�+&<�[T�<xԛ�O?q
h/�¶)�Ȥ�����b[����<T�A�B�?I�ד��MN7#1�x��CCV~�+�ݸ�ɹ�c���Zd�ۚ� �����5�jM`�E@T���/�����^�Yx��O����x~�,��&?Gmh�����hj7����n+uMG�V�	b�9��n�u����EY�45;�K}��@�����M�TǨ̫v����a(�+������
M��J���EAe�9a�p�TY�{\���R�cн���.�{�ۨ�s�|��0����.7��9l��Y]�fP.�]�0��/)���(�_o�:29,�yR']�w���w~�H-�F��)�x���5�Iu���c�r.�Ł����T+�S��=�-���Ki�7�̷=�Cku:��RK[d��(m������~��6���;�Qi��{�d�b�Q=��`���+3\��Е�{��qN��.uk!�{�	u��Z�����&��?�#&���b�~/��>�`���`0|H!�j7�"�o���C�k�u��!>/u.>}�Ďɝ�5�y���UtC_�F��#��ʹ���=}�G`��KT8&�m�jew07��z��{c�gJ�)y�u�� ��:�u�ΰ�:�Fw1X�'�<�l�3Eq��m��[� ��̬���wn�U=�5	�����FW�{'����k�h��Z�XT^�\���|n�y��e�g�kQL�ci����W���Xl�l5 y:��N���Fٱ�Y�W��;m�(�G�B��j'5g����˖������񚇄�]�J��l�������t���;9F =KWx����Z����6�|��mf���jb.{꽎�R��\o@G؎��U�@��Ӊ׿�-ց��;�c�2���6����x�g4�Pz#��?H�
����7�N�� \�nx�<f��s��cZS[�5f��k�'��X�P5�o�|���Y~}6Rq�� ��UҊ��lJ=���Ac���D኶k�!��ϳ�B��ؓg�#>�\�_B����k��L��T
c��O�ǵv�~߃�,NjRE�V8*���y��X^�����tN5��=�a���s����[/��U�c��`��m���Y���Tux�`��9�-J�|A�<(|XdO����8�iK���ԤEsQ�[y#�9��a�2��<�|p!#!aRp�7��R�ĝ�D�Ņ^���+ڌ����q��
D\�ܓ�H�HKL7��5R�Y�I�+_������p<^��J�ԡ��>m�� l�>t��C�^��Ț����;��
�?|���^�ad�UE��a�lt~u�a���g ���+���}��1 Pt���hL`�J�������&���@�/E��]�_���.dgo�3T��R���o"���ߕ���"J�z��}�R�SI�|C06�9G6H �/��!NP�)p�n���60WRs��hئ��5��;�������ot��ܻ����x�XCƌC�����:�����c|F�,���ͯ�i��t$K:�4=���?%�ӏ�	��f� 8J�gh���I'v��1�\�<�CPc���2���N�,���A�3���.�UnoN&�,h'�Yg��1=��x�`~52h�>q���"'���H���l��kD�X�x��b�cK֎L���u	1��`lNt56>�J���3��ZS��"�x�J�(/�Ag�lPۛ&��}�d��L�h�$����<	���i�,����g��G��~��������+N�л�0���+u�_�B�-�B�g�*cB#�0tK��i�M�@:*��: E������7Z��(����}���u���_#;5���lo����a@��A౏G�mSoµ��D'�X0J�%�|ڮ2�fF���z^��Hf�ȉ� ���3����������/.o>��|����g���At��
�>���_N�q�+6g`F�f�_~�EP��%A��.˫�S�NGX�q@a��7|���%�<�;�M���όJ���s����������L������o���E8 �Ò�*�"��ᅍ���$���������NN�?jk��YS{����R@��Y���4Df��z-�U2/J��X�%5��\u��@i�`���ԣ��6:ٸX+�"K2��i�B�E�X9���'�+;%mTCLիK�G�b`�xNz�h e����"ӵ��5�)Us�R$��jX�{$V�y�TbRy�r���2��XϢ���?B,�y2��[t��.#�"�'�3��x��ą����H��ڍ�g�YtӦh����씧|�rkm"�C`Y�f��;u�Bc)�y��O �]l���W׹@c�
�$�ӹf���D�o�	L��/>����F����~-�����= 5��n^<+_��P�"�2Q���=(#��� $��'�&�N�@Yʋ-��)��C�<�2�_~��@5��^����z_���������ٟL�tݮf�*��U���@
�R|�g�X�O��b��`��_�M7�弹'�zv|�Z�u�i��0f����SY�q]�˘͗�g�ЀV�g����������C@78،�#���A��޿-ϟ��%���!n���y��*�q`�'�eF]JzGE�N��(���hL���(T�����!"�h&�j ����8�ٸ�d}35�:�.������S�\q���ׂ"̤e���n6W����'m�7x��G�N��\�:�T6����[�ݶ�9�r}������Ԡk��uf��$W�}���c����N�
��o�_K뛾�-�O�:�EM�0X]����=��Q]<C7;�Ew�=K�ȴ�-z0�
��Y"���2þ�;��R�|�7���X������l��1kQ-����#C�	k��1���@!�a,xȠ���h57��FH�=j!�U�v�{ G���!c���^�޽Du���>f#mɶC<>��uy��M��}g�w3�Nx]��QG�xR����������PA�ߥ��NUK
0�����f�j}t�Xr�l�WB�+-���H��_��۵{ ��������8�^o-�^�V`:U��q�Q
i�;�O��4�!yʆ��O��x�]mB��w���	��s�k)V�
���9S�Aa8��C'LN(D��]�(�k7�K���Ȗ�H�8<�$9��(w��W��=mP=�Õ�f�����0�"XV�=���/��79��F6Fb��ͤ��I�D�����٤�S弝�ǱY��xc'���Vwo���a1*�eI4��_xF-�ƚ�g���V��#&�C�7ǋ�7T�����,�5Me<�(=�G���)r��t~��m��F&u#�b"��eiG^�sΆ�|ox�n�/n��e�[���#��*;�� �lX�[>"���g�2	w㽀���P�xI{�"���ڂbf�\�ic��1�&&�� ����A��XN���[~����>�\�
�v1�nk�}�C�˵�����h�][X�l���P��-A\O|�>���  ��IDATߋ��-�y�]��>���N�'�<�B_��W|��.�m��4�Al��LX�9�:ÿ��5�*sbT3Ͽ� �R�ڄ�^<��[��8uO�)Rw�$E06�㡤h&�����@�����YTU�k�|iN]�u���p_޽[��G�h���A��p�_>�`����%w�f����ɍ�&6�`�����:}Dd�l��e8��.6�i}��>�t�E�f4��J�e��xt8��@�ˎ��H�����ҝp�F�Ө�2-��A�o>�S}����[�Mv'.^����x5�h��bx�ȯ��>K!d6T%�Ha��8U*-<��)sg�)�,:`���Nk�eVVJ�ƃ7Ns҆)^��h/!��[���ܬh aQ��oʷ�|]޼&&
f��b �Ա�C~�Y�zw�|�w��)�|�M����M�[�_~��Ƃ!U��Z��B;�E3�6������F��})����`�vh"}��F�0 �]��e����ʇ��۠9��Fw����m��1�R(S��Y3R����)� ���$��u�x��: �딕\��PSSHdM/*f�5��k���	�ߕ���o	�t'xOɢs��t���Z� MF�u�h�U���Urx;N;��g�;�p>`���N��:^Rk�2���5��о���0\f���D~}=	���Q�)��aZ�e��cK��W������PV/���Ҧ�˚����i�]�KQ>�c�y���	J�WܳO���AJr�"����e��7X]?Ǆ�u"����}��7p��A�f(�,kb=X��7��o#a�<Q��^l7����\ѱvC��SN�-h(]�|��@Ou�g�BQi��5*HA:I���A�����*����8�iZ�S�P�F/�8T�3"p���T6I(ci<�!DD�~j�Ll(@A�߮/�]!��RV�e�?�����y�9�9�z�Ck�ٛ�R���Px���#1X�|8G�q���̑[LR_����v��Ӓ����}r.�c��lJ�e�W�X�$�&�t ���Y(KZ'E����澦fm;*슫Mh fG!��[��� =�d=����N09��r�q؅�8��X�HL��h����}=Mi49�ZW��.�MY.i"�m���i���OA�|r6��1��б.����Ac���=�D;bVY����r��8�@�"��q�>��8���+�@as�R��&���0)t|�k�2��;r�����q�E|�O���32�}�A#��������c��ǂ�� �	Y	��>���o�9&_���f��c#�X��Χ�" ���/�y������U���e�k0�F.��p�h,Ɒ��rR�H�!T��Y`��]�|�YP�����l� J�{͸��R{��f����5d�L~���*úy�(���`�� �#�ZCЍ��C�bd��R9�旆�������O�6Ξ�����y�}��2��!I��O������x�2������<y� �^��u�����?��1=O�.�*�����Y3��Cl�Tx�!�Ɗ�9DY[|v�]{J�ղ��6���K��2��F�X����1���ML0+>��L���:�Y�߽�eN)WǄ0g4l�۵&3�C˅UV�$n��9����Q#�ss@�N�OJ��:8�z�@�|�H���Iٸ��U����eqt	U�=[�l�A¶֍�ccV_�J�<1��1���@�C�����@�#���G�16gC�]�$`��i,lp��&���G'G�W����u-9�Ex�j�q�w��<�C@ WA�:_����K���J_�Z��B��^n��D�(X���
��t���v�Јrv��|Խ�H�h�BX���ͩ�	�g�l�@j�:.HN�E6�VM̀"���M���8,�>I���v�o����J}�x��3B�C�4��e�1����eqt�����Ѧz��~�Kg]��.��Dl�M�]܇���l:�ݟ=�A���r�?0=]'CP� ����I��w�+�m2)��Z���n���.��j8����2St���^\�ģc�����bp�N�S�$��K4d�<��t�{�ntʸ�5��S��j�rֈ9�p�݅~/���LFPɀ��e��
�O�1����ϋf�Em �����c�Oz/�-����ׇ��5/�.G-�r/B�$A�hh^āA�Z�iј(�AP0v
�y�5C��M��`����М YY�	������+Fʷ��jQ3S��=��v�L(�T6�������jϮ>Ns��av▢�t���)����`x�8dH�����==RX"3RfX(;�����������%���:l�b&�>����k��@D���Y���޲��^������ �Qu7�@�(#���=�*��@+���T~����e�(ȏ?�P~�(d󠌕kq����&6��|S�뛬0�8$r����;'��2����������ʅָ��$�oQ��,����n���o���S�S�����o�~��Ͽ�A0)�d�z��p����K���3��u]iK�q�u*�l)�#���$���%��J�kf����`��A��؃�cMF4,`��vأ��W���Z� -V~���[�Ł��HQ�a�hxd�S$${	�Ԅ��z�fDLEIi]��1�&N�����\޷���~�������j:�?�
�d�Υ�"t�B�d���-ܬ��b�7:�σ7HG�3튥�΍�i��i%Ǆ|s쒣:��$���ߧ&��"�-婿xT��1�zz�7J'��}�]�`9_~�6JU��0����~|��82��~��%�n�RY%2l��neI|�^�1pD�H�W���f�JzJ,���i�X�@��h��C63kS6Fq�"<qG�����QLKR�X�a�}{��ɻ�V��}6�Ɖ��2���Q���~-�%��Y�`�*�/�����w	��G�=���_��~�{;��QnS+76�̨��˲�&r$ѓ���� &����={����k�������?_�|���px�},_5A_�s���� *�����AL9WG֞�x�2�՚��`�(�+��O=�5�F�=�tK1���~-O9�ᠱV;@S�隁���J�� Kq��Z�x�u�t���nt.�@8m{��m����Թ��f�����t�6�>)�/��"|{Z\�Z�΋dy¡|��K�U�|��E+�v���#�����Re�hG��jW2+���n���X�婘"����v�Y��d�}ts��U�),r��a��6)F��0��[d?w�F"0h3}�㣰�ƍ�߁b��e-��wDC��N�Eo� �at����x�G���۳�1��<�A��n0EI�%����ܨJ�a�������TR
�;=�1������������[p�[\�\Q����qO��Q�2&dǯ_3�����+���#N��	L���.՘fѰƱ
�x�x�������3��g���ա��_�w���)��u�Ѥ5	ܚS~r��E�|_<nI:����j�'=gU������kv�Ro���&U.s�4��6_���|��=�I;�o*�1r�wÒ�E���/N|�����=�"J�=ଝk�ی�x��JZ��+�%�q�?@?tf��_Ү��H�������z��7�-'|����&A��~��N��x��t���>F�0�@m�@^@�H�ߧ�.�N�)��I��T�-pȓ_u�y17v�����.��(��+}���TP�-н�)F��Ѳ����D�bF��#�[�	-O`�hp�u.����H���xu�_W%�p�f	uu]1�=�H=������ڡ	�##=����Gs6C����\�Rz��!�lD���{��������Cu��g�A�@����������������Ͱ�U�����
��?
�-5��T�APBs@��cڇJU�?�c�z��W�7'�Na����}.@-0��a����Wo5w������BG_�Lf�/E+��;$�u:��
pO�rc�L~^9i��b�����d�w�[j7�2�"�`Fz/і��8���V�E�$����Ie�
�"Fnփ�9�*�؟8h���FV,O2[]7�x��}φ�f�A�v:�1f�U��g����'��l����?��&�*���I�����K�ɥo�0mԯI��&@Y��[�:�,�`㵽�հ��lY�(=V7F�R0�T�:X��K�9UD��X���<��/1Z�w��׻��(WW���� ��l���uJ�&�p*&����o��SJ���gP�y���M�%�h#�c4i����]d�6U,,���F�̾L%�&�̓I��������G ԰ٵ-h��V����@e�_���ypF�Ɂ�vG�1+9����(,��,��V�ml��Y�ڠ�f5'촐8���8����M_,5s�e��ξ'��8��t�2{�Il�G(�o��/�]�U���<D ��>�2�e����v���"4Q��Oe�J#򞹤J*�(��+�����������(<�x��3����.��!�(UY��eb�� 1k�ӏ�Q�$��X�3��b�Yf׼5\T%�-W�����ൟ���S��|���3e,տ�������L]Z�7�?^ ��T�9GlJ�^3ၕ=�������iv�y
�<���,�7i��<f�	������8����?�Yw=�,����?���'���A3��Vc.��Ƥ�N���,��$�S۴���ߕ�U!3 2�㣂ω�2�� G�o�5�73h��|Q:�.���޲�����g��C:��[9u��t(��7���!�l�e]Lu�%u{�Qh�zѽ����DK�W!%xw�<2�'\�y�*&��䲛dwf�>��;mY�a���,�j4]�Ze�C�1���MH��JA��g|�uU�ULg����T#Z��`%������l}!.x*�����U8�v�O�W�c�5�2���A���{�Q�p������UZ3��˔3�[��Lg9��x7��!��|�/j�ӕ�!8= ������N�׭i��s��	��]�&��贸�|B���%��IH�>Q����o�5�_�y���,��Q'>������Od.�E��{�L�]���3]�w�кa��XS��؏9��q�ܐ�I� �ȴ)�a�Tܗc���t.�w�����Pxz��u�'Q��<r� ~��3�"@"P#-G��u������y�Q!�b:׮�>�h2���0˳3K��*`�N~��3"�.z����*ȡ�A0iZ��eb�t_r��t�}v��/ބWՋ�����תV8��'�13M6�J�!lH>d�b�S�@z{'�)����vV�*�6�8������e�.|t�52i�A�'|&@R!xk�2rخ�!���b���7S5�&��8OY�[l;�G���&'�o�ZXE7��	{̒匀���!���K����]�Vλzp�q[m��B<ڬ����{v�\�vP [��gC��&�ux�bĦ>:���F����<�]��~s@+�4��b��f�-�I�k�nS�V����zp-ހ���%n@4$`�L!�ҏb$s-�!�J�A�/fE����|��ӹ����8�y�U����+� ?��j�KMe�W_}2���_ߖߐe|���UF
u�)4,��)Q�2E/r߼�T�{	i�NA4�-{z��e
<D�>�ʌ� ;�ef)֓�o;ZHk�d���!����©��fFhT8���GRW"�R����*Kr�o��!a�\U��pƋ�xY�c���N�K��X"�7yn��g��������}r#-��=�#�<��~��DZ�|+��0n<gFJ��}�}��(���>�8���p�o�鞥tU�EcEp�Z�u*�P{M�H�a!��vD�f�
��A��R!�0��F�$	��s]��a�����"�u	
��c��2΃���i��.I��P3R_/�C"��2���k��u5#M�o]R�q�,���q�T����k�/���=��]TF7�������P<���Z%��fPf�Y)'�]�b�uF��.w��?��å�񔾙�������vgr�@�Es��kk�Ic��[�|S.%���A]ʁ�͚�b����A%�&�.Ơ�ס6�V�������BlZ]��5S��\Ӄ�&q�����t��2�<�m)����Ta�uM�{hJ�I�4����w[��ߣR��w��ML��V�C���l��
� �'|��.�)g�p�>o�Dٍy�C����Ϙ���]��N����D?׃DU|p�%h]S��9�J����m�Z!;�����0u���C��&�t����^L�MբU��Y1{�m�Fs)3�&1�����MMj09� �A�WRЭ���������������E�	3tM�6���&K��֪M�S�6 ^`�Pk�ZkH3F|:����NB�=�X����r�%�L���tJ�F�I��.:��^~�}O����ғ���<>1t��X���g��V����э���ލ�!3/� ��_��KhzFp���� E�l��
.�F)�M�!Sk��`�N�.�@o��ٞ��N�#��������|9ZW�^�!�좊 K�W�x�_����7+��ch��S�@PQ�W[r����Tn�o�ci�W��JI+�暁��������������fv���m\�B�����<���
MC\̛�y��ġx�ֳ��2R�j���G�H���Uф�؀ԙFVgv��Z�f�a'����@/˚��e�ChLM]K�I�a�ks�CY���{����*�޲Wu�c-���8#D����r�贜�d�}~����I�3JR�� VS-u��=j��wc�H���R� ��Y�3,ӝ�c��~���MO77�?ٵwF�6�yZj���f���dB������#>���tb���)f����H���^�u(h�$14�6A>��Ѯ�C��P 1=bn4	gQI�����L���,�u��)@�Q>'Ή�� �E������l݂(g��S*�t�pW�iM�q��'�N�>�)��y�� ;mj{��U��t��z{
y�I�0� �o��m�F,39�tl<��
L0Q��v${����V�8Ȱ	���?��`�i������E{�������[f�h�Dvs])��G�ܜU��b��Kn�_�ɦDS�l�M�˷i�Rg�:���G� %�@�������97iCs�n���V�{gIʍ�y��6��w��3e��������ֺ�a�a���l3���`�6�A�4�e[0��q[���=xP8s���1ى5E��Ks7�}��C�oi�����kVc��t���C���'0��
�����1����E�DJ�˙S�,F���hz�؟���*�c�*�����k�굃f��R?�ʬ�i?�G��!kC�r�[唝�x-�K��X�X����Mau~�vp�ݕ��d�F��*�)�L<�+�=7���dx�#SZՀh�+�1L|�b�p����
Ii��j\y���kg��O��%��i!�\ ����r{�!��Pjڂ�*��9cbE�r�*�D�$�?�! ���q���۸V]��\n��L�����!�o�A#�0���^�0p�C���Wu����]���e|���x�".���gE���`P��Y��Vxj�tͿ�}��V?�{b��ա��7|��*j�<�6�
!����A
{n��y�����0q���J��u����3��s�k�\Q�`L0�"^�)Z�������sm����Xէ1�4TR�.��Zi���L?���i����PoN���(Z{�� S.�H�9g{�����i�����D��H ������xg橖Ķ��u	G��\����g9�ҝ�,Xl�~�rŠ���ͭa��=H�}���w�Y��~4��l��ն��L��T������V�)��h(��-��>�o+�`���i~�L�#��-ʀ���4�1���}nw_���wAm��A��:p����n��]���A_��:p�z��O����F�J�R�M[@C���g/��B�{n����v_
I�iӬ�c��n�)��h�t]�+߷�0�Ȑ'Nt�Χ�����	f�n�z��yx��@@/�Q�Nj�q�l��	j��^9c�������1GF3�j�	+X�����a���'n����^������aIf������g�6h�����9D�K�G6�յw5�I����,Q`�� <Ѐ�;�"ڷHR�g��^f��Uz�X��$ᮚ���i6��4�E�ާG>)�JF�Z���3U!f��a�}H�(H{�o]~�L�פ���z�8b��g�2���Y|u�9|�����M��/�?K�#�f���.K�LC(8������n�2VdG��F3I��R��s=_��d��l+�pp�zHy�c���cmW v�6���Ǹ쭭��o~tȯ8���� 2��B�����W*�8����꓂i��M�����һ���y'���(����fP(�Ϲ�.��5�5)�`�+]i� ��(d��S����lG(�X��@R���!��`-p)�a@�u
LT^�2O|��-D>|�n@�����jaq�kL���M�q�؛�m�Y#"�B-^����*�A���3h��-ᛑO���҄%���I�z8���vQl�ئG�92�
��ì��6������B�Qe(�_�;�V�yټ���pz���c�k��mk��&�Y�O�$���N�b�|DT��1�Ҝpܨ�������0|Ռ��J-(������p(�P	"36�s��et/A�#ձ|���0�>R�σ����97�²�Tq��L�����|���BJ.��f_�npK����g�^L�Ш1p��1��}Lė����Xٸ�c#/�U?�|/�f���:�P�<�!=�&2��xy:(v��o��t!��	�H�49��2��Ha��`j�2�9C���1�:�l��W��l�:�4'�D�������ܘ�����}H3���׌vO��b�G
�m�7&�0�QH�7��k�{iZNp���v>||�������(�L
�#t	���>���l����䁖̎�T��M��������\�a�1W|2i]gañDs��׽h��@�L������<�+�sV�7��x�!~�.cm<6��,�g�_��/����w�r�ػ�N�{ǽ�[Cym����z>m09�V����9~�_X�(��B����Wp��U$�/��� -���L,�=��Y����dB��d7A>�0��Axd]�������)��"��Cܽ_rʄ��w��:���#n4��a�g�!�{�A�3�h�Z���ʴ��{и梲�*{��n��D����{����ՃG�6>Eh�.S.J��c��5]A�&�z{�BW�(�~�_�iXO:��6�	��
�0[wӍ��Ͽ�"����B����M9e��k��繍�a����hfK�	g���>��r+���O� ��ǿ�sBx����S�Lk���n*x?(m����j>���d���U0��)x���Z7x��={�k��J\��V�xh_3�&��v�%������΁����x[�Յ��gۺ{�g�hL{��`u.���2Y+4����K�6���gńɏu/'5RM����լ� ZᲊI?���T�#�S���v�Zb�ɯ����zj��TK��8��Lc�8����9�*GO-E"�z/Z�GC�;��iY��"L�v4P{�iE	�./\�z_,ú�f�I�u�q-<7\'ZtE����28�.C�"f;���£2<�r\s����״R\���������#��h��Zet`I9�%6�����M�𓺉��Y.�4��4j�������%1B���� �G �b�8$�NI���޲��q�B���̝Lf��)N��C����z�n�UNj����(?��}������T*���FMhb<�M�譆J���|>����bB<
C4�t�Ӵ�:a.�~����V�@$\�,Ns����m��9��,�Ln��� �aai��6;Y�������j�u��	�tf/�k�,CMgM=�S�Q�=��"iXm\����:�U�w�R�M�t�Ƅ&�����2�ܶbz�S8$2RߌR��ی�6j�A3�p�xý"P�����.EL�
�G��V�h`���-�H�iF�WzX�Y� �6��^`u�����Z�)��2���A�62��_5Ia��4��^o���R�EYKSI���*c����M�=�0��< ��N�ҟ�.��&`�:MiA C�̍H�W��j堹y����D�얷�5�8�V-�潺���:��a������ut3�����c����c��pR�!����AU@,ϼ�!��6+N(��*U��_����>�ry��}f�2)]�=!�Mﮕ���Y|�`7�Y��9����Km�������:�7WwQS��X��vи�a��{$(�!��� Ty�c��&��_����/Q���HM�*����i���X�d�ܗW�(Cn�!�8�g�����}�,�]�z����2��I���nbܴ4i�o��z�8J�g�G�b����N��vX��4���b��O��C��]b!��FF�����]r$ɑ��{\���
�*���r8�v�����2�yCv7�PH��׺���Y$��9˙藝( 3w35UQQ,�����'~�<O*��S��M�t����͂w���e�m6�f%�O7>D��C�n"X���]���A�n�"3����Ŕ�a���`zʃ��Ʀsu�f�e6vai�ꀳ�̠ź(�3E���
�~
��q;Am�N�,�Հ��L<:�;+��%]ދ��Nl
n���0�,��A\\i��Y&[�SE��Y�b�{Bɿc�#� ~�� ~��r���VT�䍦�y�kŜ�W��j��}�6)M��>&�b��SVU��J�D�\���3k� +w�#�6��k>H����o�0m2/u��QY�-Y"�X���s� `�_�52�A=_�\S��U�c�]]Kg�5ȭY���k;��og�WB?�Ȭzƾt_d�W���&�V*J=S;�4̉
c�����?���v���{�;�Z��(�����Y���T�oN[�,�y��f*O�B�P�Q������C^`(]�OY>pE�`���"��f഍�e�O�"^+�{��H����u�}��hDl4����m�4�_�>U�v��j
Ȑ��	#����;�QH�8�ח)qY��@���.�1
����s
{N��B����r˚��O���/?�İ���Ҳ#�Q�_.T���/=���sP]�}���I�R�t1�d�FgA�V�/w�3PF�r3�Р4��cv���or��,
{�}&� �3u�oDo���Vl%s�f�����,�C��Uԉ��=~��М�*�\�&����f++E#t7d`��$Q;<��͑HL����5*��'~�g�=�'|�/�,K1SХ�ȴ��s�@�ڬv�s̸fk!>^~�x��<SjJ�a�ԝ�	���$�1��R�E����w9v�Pw�X��>;�(H��3�>�N/�R9����|����+�����P��"���!�~���O*�2�E�F��Y�k,�}t�Dit7K dR������m����������0dَ/�8o�������L�N��YE�����	k`40�Y@�! �|/���b�l��'L���s��1��b8`�O$��0GkX��S�o���.�k��ʪS.�C�%V�Y����I�D�� ��̟�����qA���Nѥ�쿼إR�5���$�F�g�T��u�e��T3�P:݈W��۷�۷�Rl��͏�|.4Q� ����$�e-��sc�ڤ�5��斮�s��YT?T�J�=}�Y�1+M4�N��**X�K�#��rۓ�3�|��*���`��yގ��;�O1k��]��!T]^�g�C�\]�(�׉�vo����}�N��:+N��R�tͰvW2�n��=�X�]���@%�Hkc�f�yRu�y�L4:��;�u*��~�'�Z|S���0<��ɦF�U8���jH�{��&q`x�2՟�pqȖ�0�-�o����Ϳp�/뒥I��5�T�̣J���q��@a����W6�~��G,_R��a�#(�W�s�Q���n|�7�ƅ;%�0T� ;?�y��rsL��Ԍ��Κ�����c�ۂ%����_�o⯃W�����5���Ҵ,F�1��`zX�54���֭*�p��������mU���`�8L�y�-��z��!���d���c� %�[��G���@~Q��|n��L��P���ݧ�xm�|�� {Kv�`\�M0p�h�In�U� 5L�=�q6	�t�2t�Н��m�4���15�x���2�U�3��8G&���wXJ]��w�y*�u����̤Bj�s�w+���Z��\·���`��FC�"9ʰc2�����uu|ׁ��P'��0�z�������{��9���<�*�%�g���É�����h.�$�@�i[�b�? EɄ`�E�@�����LQ�+}ɊO�QV�uqs/դ�ۮ�*�*9=K�R��r�$���*~�L�����������	&�d�%7E8b2���z�εs�1�9J�q��{J�q�;�u�$ h૯^�Nde(��x�S�FՇh@���� ��J0��ǁ�<ӲbV%�0�m�m�����kq�]UWJ{�NՃp�"����Q��#��y�0*���B�'뚕��Hp]�������m8��C|u���c�����^Q�����nQ��z�4�@�m3��Sgy�
�;��D9�a�ґz�DV�&���5&q_�;��-;�Tq�R���b��e�.���Jdanژ��L����ו���}����B��������*�KŴ�k�&c��q	��+U4�Ү�U��e�`�y����6���&����6S�oÅ[p�\f�͡��J
��a��hfou�1.�S3�.\P-��5�L�F�Qj�^��app�4P�q�e�#X(�f%L�x���a��L�P�V�u'p]k�~���i�0��[|]lB�~��w�сq����+ΰ�X)�pS������m��S{�
�����d��SO���E��O��9m��Y�������llt��Gܘ�-c�l$�1��<f�!:܋c꾣=��>߅�SnԶ	Q�+aY�Xb�ŕ�>G%�r����
JP?|�gգf��َ�I�u��v��[0�9�sz��p��(VUs�&pe@OB���,at���v)�d��ş[EGwMA8��ȴtؾ̃p���-Ȇ�-����)�°�M�C|g�`HZad�K���d�Jr�m�U ��h_�@6��Ftݷ�E����8�:##��	�̮�nD��U1L��ؕ$hr	��
i����'=�px������C��:�-ʄ�����3N�=�l����Aj�i��ZXHk��C���RͯL��&�s��Z^	S���0�o���J�o߽Uix���s�6,�i&x_]}��>3R��)�Zx���*#�Fj6�i���:4m{ܷ߼�'�?��?��a����'��'~��oۦ��ӧ '�$��=�ŀ�fVt5�i�`�2�e���w��wߕ������g�Pa����Z��c{e!|�?[���EKY�0_���%!0&�L���e���4�+<�|�8Z�"6���5�WF���)�ߐ�撟K���a���/����q���P��}Í}G;�;��]�>��6t��h-�@������|���1�k�i���챌ƩrY���}�����sY�w1��EsP�i)�?ex�A ��vH ��sb��H#˴r?^��̽hyd�\�rB����8�����9Y��ڜHE�=k)Ⱥ����r_�>�_M =�w*��^^��mP����U�?3ԦW�9�Oo��D1���R��_��?��*�*��W�hf�����|�8E�f<��S��%*��S �{	n�4 �������F m�����~@߼�E���U����"H�b$?2�͍��NT���6�\E�l�yьS���}TS���q���9�6o��9�8�0�1�S�p$��0�υ�:�8�lI��;b�k6"����}X"k0�V�����f��{&�a/�k\}����9-*w���
9��$\��Z	�s���2Mi����˟C��/巏����K�n?���G�����F�g��4��{ҾUT��\�`���~�¸��
�Y,XYe�Y������R;��X��C~�&

 �@��@�osp�mRfI�]M��Z�\�UW&�k��TkҬ���^9��l��4��_�=��gi�Ms(#D��d#0����Y�-�ݯi�`rc�����1CĮV��=�������2{�f���Y<���%6X	\�	��a��Z���.��w��w�����ђ�
�<KL���Ҝ|���u�V������XJdbKr��3}u�4^d~�	� �+k��G%CNu�Bxn�)�#H�<�d3Ɂ��#�J���8g��x��/5oN9��6'y��$�e���va�w�9�]s��<$���Ķ���H��P��>�	¤�r�����B���m.&ܗ��M<��|���M����Q	�P�z:�Z������� �Q�=6����MnX]���Qy/L�\Jd�yH�5Ƌ��E3c1���6���p�>�A��b`/p�>)��A�+?��.���\<�7�2ј�{�?Z�8A��p����e�{z���Q�2x���,TYf���)�)�e�
9�D��4<@���`��	�f�H�WZ��j���J�1�����A���Q4���j�ղ�^ex����d)�_Χ[�ߗ��ɬXG��U�1�}�@�`�}}�&��S�|�gO�ipg�-@���@�N�������Z�a��n��>V��x�<[�,(
}��5�s��/WV~��1;;�ݠAYL��(�)�1�hc}�N�m��,c�ͥ���I�d�k��bmH�}�A��ӻ*9�Ċ�Nu�_�2�\=(ܙB2{)ҟ�{b�6ⳌX�3�'����w�6ǭ��?���CI~�j\X��iPcm��x���5@P{����iul?Tzת9n0�m��?���y�]엟%N�)�7��(�RW�&���|��4�&���a���e�� x3��~��Z8.2h�]��]�aߗ���4���F�~	��1�o6B�	���<�1�UJT|9���s�.4V[�ԣ�]TE6��A�n?�,��:�0c�؃l��(����.�;/�AaӏݣDZµ��}�u "|3� �B9lB�=�����H�Q��V�����u��s�U����u(�A�jzw}���������jdm��2˒A��h�Ԍ��{���-rRG�E]ES8���:����a�(e)�N��P<�CԀYD�y\%&��/Vy�ȈQ>,d82�[�%�1�fN9;�@z8�W'����3j��l}�y.�Jji��4���u[�R�77G�kjA���k.���&*w�Dtl����&�w��x�,�����#P��P���H�Rq�Qdof��<1��uf��6�yd�B��m���b�	ҰV�(��˿������|��Q8�OY���`ĳ�w�BAp���D��9IRmb@||T3����]p��bM���4y��I��a ����)�a��ӓ �K4Q��/��n� =Ji��1���o�^���{|ޢ�D��tp�j��ʹ�E=���\�j:o����jU2��.�;5&�]�xo�'�U^�j�-M���F0�
Xe�N���u��nV����jE��$��H�_��.�#⿯����U��73R<O�����:�F��'�`	>}��rIc��]���B�������٥�5�>sT-d`�
l����y�{j��.aUw1&J<��F��Y�d�}\��,!8�M Sm���k��g~����x}�JB\�;�qL_�����Z����2%�'	b�	�&�*M�\��rtq�in*�%\�X���J�Q�\aB_�5�ΕɲY+,7����ǘdy|�ͿN�Z(YZ��Izۯ��/��*��/�J�;1<�>�a;��������m���샎�GeM^mMO�!�y�
6y�lҎ��Zƃ�b[���p ��ݻ�Y?�&��l8�;۫!���5�A����_�� DV��tf��|W��]��ޮ��/c��"�d_��͒{{MU`%'���ǡV��4s"g�]ҏ���ág���2���R��՞�[EU���kl���m�3M��|i~�k��RI�J	�xOIHD�Z7x��$���~}tW~V��7�8�^�^����&�6���a!�>�t*����i#��S��b��O4�7KS�� eQW�!S���������_���Ngv�倫�[#�`�h��o��J��S�$l�_�p���n0�c�0�S.QYV�� b�n(3�([Ks��1���86�m-���%���LY��ڔ��΃��D�eXɠ[�-��=�g& & �h#���NZ.�1Qt���ŽBP���L�������O���筤W#�xv�A�T���f���(zJz��S4w�@ uy�������b~'���S���n=p�A����*2��ۗ$���p��ÇP�*ѐ���N��H�@:���D}e����/�<�*�U�n��֜l5tG]�]'�>�T��EE ��C�Oc��ޑy.���$~��@��Z��@_�ރۛ�7K��6��X*q��	��x����g؍�y��49�Lׁ�ҴL��1PW����9Ú�C��^��
��t���8S�xq�5�e��B�k���kDF�i�{�O<Vb��ɵ{�R�H��K��ݐ�G�(��;̉��Ϯ�'p��X�w�Vz�馌iS�.3R�[<��m�
��gn&�~A����>tQ)N����@>G�9)2�������J{lLa|�E��zJ�C6[dC0I�%Iٚ]�Ӂ�V���<;�ȄrI(��k�*.YV�w<G��ؠ,�3#�F�������?�ݲ���.��4���-(���	-�'f��Z���@��O�JWz�V$����\�F6,��)�.��n'��DPΩ{������'�������}���t�H(4f�܋��i2���@!��*2WR�愸���a��jR:������xb�lF/���T��r��S�5FUoȍE/����.�!?dS�t5����eL�n�}�����������Yk-�?�p
ރ�JV����/�w�ޅt�%t[�!�T���Ͳ\�	���(����/��x��@<�0Q��:�^C,�P�c�-FZ�JPg�Y�!3X�+?v�W�/ty��	=��N!�[�u��͇]t������"5!N@]�]]� ���cF��w�������e]�kԲv��g =�n1қ[b��%��\F�'F 5V�C����9bxP	C��̓��%n��5`|#�=!{
1pY���Kg�5��]����W��n�ajT]�ՙt�������X���Ǟ��B��[&UL�E��,w����?3�y�f��ھ�u�㩻�i���n�}����9�<�Yb ��8p��2(~�	zM��Z
�Ja���
���:��\�g�X~���b��_}���^�Za@�\���7~G�����9��б�Mk��z��*q��ԇ��Jި)���Ͻ׉mOUp���\b������S�-TF�['�RMB����̨�\;�����R��?�q�ӆ��2/�0`�s3Q�����d3��PKƷ�;q�M4�Wz�]�S��d�5t�򺏓G�Y�׾U�7�~��I:���%)No͕+�00WˠSS	���s����áR���w�@�a�s�{�9��L��xt����#���tִU�y�Q4���K���$��R5��8� �SO�Y�SB��ϸ��:B��*�/����2W�-;��jW�,���l\K9�>0��xX�/��*�Hl�����<=^¡u_.5(v���m:�M:���AX��HC���o>�&���0Bl���O%6'���!D �P|�Fm�L��9����>��W�_�y���E���.ɷ��=ƙ�
h�"HB�?�^����M�k��$�� ԇ-�Z��Kt�`2�9�6q(�}�<�x�N���m�a������E����1H�?���T�|W&Kp6�>esNr�C��FJ٢&�����1�l�Dy}a��\p�����>�v�6̂�_��l�?��W�P3S�t��-�Pi������H���*.fRy���i۶_k�i]�Id��>|�'o���|߇c���.���]}�N�o�4;�$�K�\���d)Ԍ��	���5h���1�Z��8�iU��K,��m���,>�5s-F�Z�a�ټx!�%9k�q�]�=9�0��,X;�$��EF��/1��;�����-K`T(	{�AW��)f��k���� !?��^Kf>Ź��S�T҃��)@%j<�$9w��,�b4"�s��lΡ�������w���0��?�(���=+�q���Fe�1w��W[���¸��ޱ����*�:q��G:ǄW�Ȃ9c�˯œm�,�gN�!�d8ĸ��M~:�����v���'ѷ[PG@���
�{f�m �J�!���)��\�8�8D<�[{�k�˩�= p�z�6����@�πr^J��b?_����Ͳ�.�(N�H����y^��IH�c�N���K������%�a��=��	ASN< �>gbe������Á���ki� CPL�����gZ��u���gy�#]�����ȃ�g����eW�AjF�{�h�W7��C*�*�&�K6�y�E[R'ؙ�1�|�t�7��s��'���F����%ʺ��|�^������6>F/�m���{�������#mT��)F�uʌT*T���矸�+޾�}�n���Y08N	vBW����X��V͌��y���`N�))��-�9��߅t������� ��Q�q�`�̔���A/�y=q�p�_o䙆u���!�A
�9��*��#�)k}�w�3 �H͜�)��Y���w��kS��1?�d��8[[���8��Dy��W�_DP�WE0F�����Ge�����/&�N�����&O��������`��+
��:�f�Z8ݨ���b��D���d���S���^�$���4S_�yw��������,�b��)�Y�x~J>�W�a��	��'�I�H\p���)L��Q��9�x�~)V���� �-۟$t� �tb������Z��`��XӿJ���'���Qz!�*8mV�S*NOy������I�T�A���a�b����Ooys넻�}�l�"7��%���[##n�Ag�&�㔂d�g�=����H�7A�3w��ж8��NK�mG�
��%���ڞ_�"ޏj��ı'�5���nn3@Æb]�A��P��خB*���S?����k�Y��C���Þ�8��yW�/5#+a�{�����u*;�UP�J%��>����?�#34�~�����&�?�;��9�h�⿱�����IQ��DQm�Ϝ����۷Qb�x��i�}6x��y�ÎU��~N&�����x�߽{�l��\4�°�Cs���'Zd�3��ɦp�<�Εn���
�2=ixq `��ݮ'��J+x:H�����l&��qU�e�Y��@������hX%�������r�=���,LL\w��l�Y��n���Y�h]���X�vϐ��]��넱��[���σl�+<R�,��b�����'�ˋ�S-cfj.c�-!�'E��OUO'����>;i��N8'��A����HE%Ѣ��s�3���;�v���ob�ׄ+�g��B��'�;e��&ӳ�c��v,�n����=3ҋ|���|XGKX���Jɛp{����^7������C�t^�zC)_t7�U�;$&���gO��i�5�)�$O����#��,3l�GG��`������(�Ⱦ��8(��Ǉ;� �Y����]��"����/�=܏{�b�Ǹ磈��~��������-֬��oY�#CE 7����P=�(�5���.e��bM�bX\c��$���C̦+ F������ .!kc���5Ք�>���ܥ���u���A�����!�c�<º�r���gT�Դ=Z;c��k��]4��;Y�L�H���!��Ӱ��Cb�OOUO����~ga��A?��qSȰ�n�ȫ�+�H���c��j��6����M����vב�Y���fSl)��+G�h6��d�%��&���꺨�y�Jv)%ʩ.|i�7@ٸwv�������� {|��
�9M���;[�bX�m�{�u4�v�	��D�g�wp�MG�_���k|��?��?�	<�\;d��L�,�xf�C��iqSOAZn2Rw~�gzN�MQ��AT"f����n��X-0�x8��l��f��h�Ǜ<�k�?�u=�۱����_P�z,�Gr�m��.Kt��u
�\�2���`J�Z���]���ZwP2n�.88~��G�z�l=+�o�޲�o���=�3d�*E������?F(�fd��k�A��3����U��?��O���%5ǁ�E��z�e�G2�ސ�"��'�<]�L0#��L�%��Ԃ.�\3R�.��--ŵP��\��:�}�@���cc�h0���>ǐ����P��-��㣦��]϶�ց�dÅM��;n�K�.'��:��wŕ�S,%�t�m��U�q*���E0~jL��s[�����������oF�����H� Z�e���9�~A�j:�J}�RԦ����xB�"�SӐm�FbN���58eh+�ݒ7�?�M�<��Ǭ~���^R��(�J8R����g���#m����62 ��92x6G��TƂD��ݜv�����7��y�&�����~6/@Cn�`q�~%�K�Ҽnk��*�i'��@�Q:,�� Z
7�n; �}�K*�)�51�L��#���g5
Un.*�)���t���q��n���?x"e�qQu�q|���:��`4���|U���P�#�}�M,6*Hњ��!&��y/�F�m�O$:��\�:�7���8����ϗ'fy�`��������Exء����c�&����4�LO�\4��߅��3E���6j�c��6Dڧ��8JZ�wY��K\23�H2,{�5�Xdw�ߗ��������DNK���]�o7����������.&��p���R!:��+Ҷ�h�t���:���!���
���䥝�kjۻh1�/2�6�u�[�c�䳙Zp�T���>�Uc�ւ�Ԉy�%�<4�}v�G��RC��h\~��>2��cz�.x��Ң����R�Bɰ"�����c{ &��\R��e���Y&�V�����X��\� �2��ڜ�d���������Y�����_KS'{f�/ev��@�_HN�$��eu3N�1�nw�a���.lc�q�񿔌+O�5u�Р��w���_��9BX��y��gW���Zb).�/;`�><q>����������7�8d�@½�Ͱ����o޲�|p��\��JM�c4"���-��@������A�+Q��X�Ct{�l�\_H���<Q��ٵ��!E{%��9��5�Ws4�P��=�����0N��l%�w� ��b���V�/圛}Y+��,O���4ɇ���	G$)L$�J����3nՅ��\�� ���1q�qʽZ�1j %�wx��X�Ɗ��&�@&̋b�V�r����m ��d)��P�U(��tK��u ��~�]2\��iҸ��������	��i�_�-�k�{�0w���@�2b��齻�%�p4Z���!�Cl�9&5��1g�����RK4y�UӴ�g^���.�-��p���kf@����s#�A'
Eh���m,k
���tj��*o#�����O�>0K�H$6:�&ў �:mL�d��K�m�S���z
���k�`Gn�������;3�Ȇ.Y?{%t}�h��bi	�텙�2сYX��i��r��F�����Y^1��k��w��A��L�������4�/�����
m>�4��Y�;�����m=>U���&�����̵`��=f�_���l"��E5���R�������o����r۱���dY̡��� >� �� ��wwK��?�q �ґ������'��Y])Y�e�bZ�9����A��:���,S[f�z�XlȢ!��zU���z ��)x0���j���{ux0�K�=�RO$�C��vekTF�0O�>n�{"�{��.�_�?�8�hZ3R_/<���646�p�3�ps1��Tlb�����D��4�Y\_m=x*��ҴC�!�7���T���,Qm������<� ����|�L���c�`K%��O�����P7G97�"C	��~����?���/Rf������1�����=���?�q"̘�/^�����_�;�5Gb��0�U�x�Y���X�Os����:N�S4�� ��`w.e���J�!�0�`_(�EFP��J�� K�)޲�`�A��.W�E�5�?7��yAWU�n�5� p�!+7fV������ՐqUÌ��Fx������(P<]���U��`���H7�ͮLHB� �����/Yv�ٲcg�]c�fXf	�^qܻ[6��UG`W���j�Ah��I���^1��ɧiv�X���S�3\-٪��F���Y��Lr��\����C^/Q�
��g�^4�A.5���U�����`�k��Ʃ��W��j,�7U˕t�4�0ph�w�l��re,�v���>W�������]��R$����HG�bA��X"�X w�ҥ��q�� *�@�f��wƁ�T���I����0'��[yG��z�@�3�ee#��:�7��<���>>�JP���ŮK��NڟbZ��vM����[��k�ܮ�;�jb]`�A}��"���6��湌��p�KN�`����w�H�>0��j��1,��#���FԐ�/]bU��BUΣ����~_e�8	�=R<B�ͷ�M��1&*amb�8�&�7c�i��T�����HqN��[9xn�83�\{?;Xj�W/�O�>l��m��5�N�3�]�Q��r$U�1��O�������9L�.���\���J����\��D�j�!e�'M�ʹ�"���kjةkbI�E��)��9�6Y�Z���k! ����N��*>����]Q�i�I�����I��J�(t�.�{��Hi�a����n�������Z����k�Ef�,V�U�&��ϐ2�h�Q5�Z�e�v� +XI���/XG��<�;��Nx������C�� -$��B����'
�;<I�'�ҽ"Fy�g�� 
�lvU4-����ޅ�L�����:_�$�&�k<!Ȗ5G
�ѺyDrs�����[H[Qi2&"�8p=�Z\1!��K��������%^<�b*
�q3���ʄܙ�
@C�pBuH����&iDM�A�D��I��>~T�&�9��V��Ÿ�SQR�B�ㆠ6A�h�����a�� \s�r�MC�mБ��0`
x훯ި���60�C� ��?Q��#e��g2L4�Zb$Yx�'�&���et7����#��jm�Z�G�O�'�N1z#�l0"ၘ�K����O���KZgҶ���goz��l�s�g��s-��5���$�75�w�>� M.���� �am ����NA<-�Ԩ�Z��zb���.E[�������Wx�|ք��
Ho����[v1�q��gbq�ͱA4�x6����Z�4�Zn8��(�MĽ,MW�^'砣lr`#���s�x�����d��j.�x���:�D�b~:������e�@�Ȏ�[��̆��.��7 X�r�7��Q
H(���Ԍ��@
���Nie=�Hi��W3�+��xщ]�:���Y�aWr�3#-�tX��kjQ
��'�aps�s&��[��>^h�@\K�["p��BF��O<^�Щ��mc���4n�>gR��yQ�!&\�����GF���ÿQd�f�����o�|�ꛯx ��NC
2��X3�Q!T��<��*��}IȬ��<*Hh,��a�Z�k�(�Y������G6������2���w�����U�{%8}��q臄�j��N6՞��$��25Mr�AW��LנT��ǫ:�u �D5�����J_�FH_z��H�>[}�}�&ED��R�?�W#�k��Ԗg�̤68�����g���د�H�PEa{u��>Lhr@�6��c]��щ�,6�Z��I�8le���54���|B� z���9T��A~R�u��^�(�ڟ�aQދ%YW"�U���x<���e6w[��+?�224[���n+���x޲���Y��Gt�?*���u�'��q����ڂ���}��Y�y�x�%b��>�9�	xs���p�Qa����l|,�-X|���m���N��Z*��香�l��y����׻��vd铦�X�`�gV���q�Yr|֧U�K�iɔ`��tʵb�̤��~u��Rkfd��(��N���i��_�T�?o�q�NA	Z��#�ȶ��s��a���@,��_ʿ��^�y\�-c���^�ం��=�C>n7��%��!,u��ތ�*��Wt¬)���uS��Z#!����9q�I�����:e��pMq��u��[�"�B�0�P4�;P�!���!ǟ#�;Ӝ�w��X<���Ont������.��%2Y\O�������TT	�l�y?;�/�~<vy-9p��k��p���9�]}���2�8K�A��&�H|��K׽�u +�Ⱦ$6c@Z�ɒ����5,�w#�S47��n6q��H�6N�%AzƖe=n�g�$����h��dC�~x��m�R���!N���
�w[ ݽ߂aP�>�߅���)O���)����N��T���qVQ@@�������[����ɱ��R|]`��H&���ö ���X��N��@=
l.YU]9r�Z��-�Dp�t'��8)㇀���P��-uՔ���/&��a�;pS��&�d�|�C�vp� ��᧟���K�j�ڞP˸����3_	�t%Љ�5�o	���a�fo�z������	���D0�t��q,�?=�~�5iEaC
����_�l����^�|�d>}*�sj��YSm��m��2N|�*đs����e�U��C��q]BT��}B<H��k�L���2�9yv����g����qv>�<������z�!yp�����1A�Oqv��~_��T�':�GOAI���@���X�
`/(�C܈Xꨯ94t����D�2ϳҒ�+���6��	lȿt��(U��`o��>�x���R���|>޶�s���q�⍭w8�p�/,��M��H_�E� x@���k��X���-|���cQ�̞i��ʹ�`NEm�D���R��;D���莛ma@_˧�ч��,)�)��j0������Rw+A�Ң���j����(N�������������w����#x��?�5���m���I?m��@�2O5<+�u��C�XJtL5^jq�\;fp>؞�i�í#���Dռ�$�(�T8ѵ���ϳ����&׶���	��W�x�2���,����4#M7���Tl^��Rv�ʙ-��]\[T(�@z)�����0���H1�
�j���!�MŒ�#;vT�u�H�x�+�e� ��5�L��v?\g$��ll�|��DxP��2� l����C֟����2�SfMID���Su7�p�M//���"���ce��EC�ң,e c<���7������E��]c�S��p8x�	�YO�]�$�9�:Zw��tO�ߠ������J����E��9s�e��I��|L[�uI.�50�n҉6ש�>h� *Kx�H[��Bn���:6X�
57~f��[�!���	7��K���%�޿���C��1�b؇��:�L��E2��(B�3�H�er&[���TT�?`Jf*���G/ �k.��Os�ۦ�~G�Ydu)܏����ۭD<޲��������_��� �F��$ħ���I0���&�>@��9�DֺӔӶ���'fF�(�2�ǘ�Z��|<�����Ĝ�x� d�qؾ�ɒ�Ko\�����G@����>o��->Rĺ� Zm�H;�ñ&X��9�!F��ȂD��/<��[��  ��� +͇�3�]���0F�"������ן�����՛a������EԵ]^��cW>�W�ŋ�+y�77/#�^�<L�h%��2.�΂L*�х���@d��5a��x���X9=���ӂB��2���-@Mg���%)�!& z�|�f�nL���P�,�>��wC	ח�_$8�#�}xM~�3�f�@!�ZE:�%� ]V/�<�O�z�UXm���sZH��v�lܐ Y�1XSs�>�fB`� � M����"�n��M�h��t�b�5�c]3�ﭚ	?�	���_�s"(Y�v�:9e��dv�"|s�Xoד�>���@�ɩ)Z�xm0��(��Ϟb¢���=) "{?���D��b��r�t�N�gf9�4�1=�lE���E�݊�;m�i
+� NC�n?�D�?�4�p/����t^F~NO�A�L��������`zn��(+�~��M����&&��x�ߧC'�9����隳d�.O�,	]�"@ޜ���&�w�}���l�� ��=�$ӷd�C�uRݿgsO��S>�br�I�ٴ���+���N0�c�Y7�| �2s�z���%J�h<�5��bt�5V,x$�/�c��3CU�t_3�uۙ��B��9��f���5:��t�aT���KmƐ�+]�ur��W���{9̊t��nS�H��r��Օ+=�K�#�p�������?�����?���h��
d?��83=i��#8�{77����5���B=���f�r��r�֘XZ��AX�^-MѬ)���2i�(բH!�TXSu.��Z�!:�5SO�FN��Cp���d2�W��]J�����æ��EM����$'HdH���>PY�$�gP���\������(�U8��E#O��
R��6�E�q:\"��R�B��0��-4Q�cO* MXg�e��qrR��s�g�f���\�jaоo�:ݔr�M�.��d�FE��9�q	,� N��/؁G#�7_�w�9~4���Θ<�M29<q:��q��	�h���/^�{��%�ws_get%�N�~���b�HM�5TWf�h83¸�&�j���=�7�p��J@7����*y^�0�*	�5\�q��Ͷ��C��]6|,�"�ʧ���'E��i'��@z��q�_�C	�⪒̼�ꛬi;����Q�N�\�����K1�fS[���	�]�X] ������V��7�\��Z��+���e5�)�>"#�M8�i{
���h�3��3 -q���"
N�@���I�����>�A��3�)�E<�x2+�ʥd�'��Ճe��e�o�dse5�vΛ�� C�5}f}S���9�}�X�+62Jdr
{��"��1�ى�=>e =�8FE@�]6-��W���Q���i��sHd%J���9�@�#�8v1\BukM؃ԣ�hZ��?�x?��k��k����T��!�G}8��I'�- ����gd�>`�׾d�.�-�����3=��"�ӖcV��SP�����ٲ�O��X ����2E�}U����4��N][X��-s��c$遶������XQ�-s&.��b�I���lѦ<-��>wj:EO @�FCy����'e�_]�NF��ɴ�#���F�ā�
�=��5�T��03<$��~a�#c�Z�J�On6>f (�9�G����}f��iFZ�F۵X�e-V��	gz�3��:`���7m�'�\���J�X���ol�Wߡ9kjfMk ��yb��X�4'H���7=�[���?M�ȧ[ٰ*0�a�l!���L�qWҦ��ʉ��}�SbKƎ}�׸�iԗyȊa
:~���}�}V@��s�җ�}�D5s=ĽH#�Q[�0SZ�:R��l���t�w��1�K��������44��:�4��a%��u�{"fU�����-mL�$���9� �4!���sd�͖e�c��Hć=��'�)TD�f �
Vj�S��"!��k6dS��	Kb�����p��l���'�4�x8&%)��W\3@��3|��s�y���M4m�����K�y<���J�L����*.
����y�7�!���5�`b�}�s'f���4���L��ji�'u%'i3��rZ뺣�%F3Ą�i&��U�k��.�6氱�9�<�h6�X�� ���Z'O[@]�!Q7jMha�q�Z�hAz)�saFSG�9-�U�JfP�n|��s��;���)k�V�� ��Z28U {������Z�'S��M`n9��"s��K)���'��L
Ze�K�1��_rI�s\�g�JO0�F�t�C,�����E�;�6m_�x��W��ݓ�� u��r�I&	��0XC�c�k��j߰Y�I��:�dR�m��~#���T-5V��V�S�&>��2Ppr1�e+���v,�jg�bjq�Ptإ�-K���'�%j��Y���?����� ��H5�S�-����9j����縇��;������K�ks]#��f�٤E
ρ� �W��s�&v�'��vR��=�(1�'�)�X���DK}A_��z��K�8�������i�2˝�c�儀��1&��ɇ�U��'Mu�A�r[˜6�Sd��9KM4N�@A�8�����]��}R���5mhhx�mG�D��fJNZD3�MM��I`���a����Ű,~X�g����p����Q)��E��VҲL)�/p��R���g�e��rZ��i��%7��Z�!���Θ<Q?E�Z�,1��N�92��}����49��%1䔶�2F*o3�w�_J��Z��(S�z�&bm����&�Fo��c^3z<�F�8�P�b��� O(`�
�~B'���ǧ�3r��z�xmu�OU��)50L�=e��<�4�������M�l�=��g���f#-�;'�nd��$�������L�,���V8��"��Qe�تy��&��:ց�8ܽ·UU�9�W����6=��{=�*����ʤ�M�P�g �����ߤ� ���� g���Z��NF�������e~�j����`��Y�;NS�Kć �ٸPy�E�#��>���.������x:�G��%�cuB���O�3g�T��5��x�$i�ɒ�*~岕���.$���}�U�d9��.��v��5�σLbV*�sd��F�=��(���F�G<�pI3n���i��P@��i5���|�<����s�
��B�ťi6�r�����~�s��]x�nn�<dOG�:݇o7�=���%3IP�\>�%"vAW�E>�8��G�y��>�Y�D>��0�����8��ۥ��dmM�> �Q�����lin�ԇ(	N�=�í5�&Ɛ��3�լL���q�d����n�fn�����r�����1U�TB�K���P�ܼ�Qҡ��k�	����Jg�������,[�{����3_<�%��}W����f�_mE��_�塹��	TU�������@��q��ε�9J}���p�ׁ_�PGO��YYEw�*�E0�{�f��V�qP�+J�ژ�n�A�U�#:��5��O����eY8��Lh��A_�YY�{I���U�ɧ6����k3d����\����R�\Y���eA`���9��$v7�6->��Vڛ]'u����p�<�L��O�gX�Δ���3_���ǢY��ǧz >��r����P6�.#;�n:��p�G�X�}Y0�ٰ�� �;�9�!����M�{��	�5�^����{��KP�4ذfl�X	G9=��wIu�W(�ә��}��k��k��ϒQ�ĵDv���׵�0���Bɫ\ݸZ�r����6���:SK�Wَ�������Ď�W����.���$|�wS}8@���`zTl�������}���k_+�z�\$_�=A�?��J]h���Hɝ�8�K<l�Y�F$O�<�|13Y�,��Zl �;�<M/cH�B[�0�gw����ύ� YLy8�&1f6�2�����zfxnN�AwB������=��/}<?�4QIk�y��M}�jU����� ����k)�LY���5��C�=f�bgR��V��+�clof��6۵ZF�?��E�1B.����N|�)�<fH�梎��)#�H�����pfe���穝	���	��	�17�����G*3i�*���߇�m����A<�����EXvۀ��X�����f���@�uOQ�h,W';Ձ�	vəxJ��i�^jZkc-D�Ԩ�}�i��J���%�ֶ�v���i��3MO���~�ld9��a�s_��P=>t��Y�|��.��%���CQ��U���¤�����)�G[$�	GEvR�=��+���uio|��J3]�]�]�6t�`N�y��M���
�?74ok��{ ��tY���B'z������� ��1!%r�>ħ=���A�t�C �#��U>f�2<�KdȘ���,J@�,��l?�ot����k�l��*���r��%����NϸWV���!q����(���y��טl�^�v�Ye������>ph�,�)2�%8�]Y-*3����Ů�������Ԅ�ի0�������&Gm��b� Ȫ3�6zS��oYM��j�C������_��0\I����N�Dؤ6���]�.JUi������n��BhИlK4��[�I���V4��C� \b�4��?Ԅ _j-_R����A�>���@[�5��:�l9˞�P�j�WMX�}�1+V/V�#�d�X��Ka��s־��ݖ�3T�'�M0�v�M۶B����#�q���xW7��¶�+e�)��*�0� ���֫���2y���������]͂����D냇_�J2A-���,�m�[-�K��3�j���d���ǃpB�X��j��t>D�%�V:��趒/�������hq$\ �����7E����}~^ә̭�#>CR�b�RR��9S
,cZi]����R��|�ʎ������v�<Dy7g�J�M/�P�Cո�jI�efoq�'�������k�K���4�����
㸡�MD<=���p}���^
)GS9�$�0��-s��v?(��y�3޻���u��u�:�QE��>��މ��_}�-� bx�c�^U�����}��~��0���z���]r}Ծ�*%6tfYό�N!���Ῥ�G<A_ժM��9��Rg�]�@[R{�#�M���o���Ȁ[G��uļ�|����_	�>b�k�v����]���/����,I�U����!���.!/ɻ��J_r1�B��D��\��˚KW�IS*͸%-����&,�D�s�'n���'���������	Y|�SY�3d����0^��rNK�1���U/�r���!��ԃ�ŲZORAx�Ćp4d[��b��e:ܠ�̾�5M�}@�Ϗ9��Nr�@��D�K[���r��������m�/�8�u�����B���Xw�|\GAYR��g暍�׷������	}���"&���u�bYj���7��u{����E)N�aTB��ԻKd�,�k�6)K���t������ͳ��W��>���b�`B�����E�64w�������h����:I���96w1s�1_k�2�ѝb]��3�c?�g]	qo��$*�)�k������9� �áB��T'��]�d���o��m�z���5�����ia<�&��{R��\��]i�9K�dG�Tu�&��}���ܲ�OL��O�!�(;�]�V���s�3�w���RZh�A�xblj���	�X\H�����u�=-�DFl��$2 �1/S�/�w�U��>��J,a;�5}m���� �2�HoU�S��^�fzs
��'m�ؔ>L<�:E����-k8���_�	!�Zm��i��RS�T���P�����\ތTqz�r{/�1�RLZCńT�yy�Li0y��`��^�d�̴;Q����������.���(��99���uB��]�]��a���=BKȸ�%��̆��W�⽒n��Ur�����j�%0쒓b��y�f~�/޼����r�:��V�A!>�0�u[��|�,J2��K(�h�l�
XKf��{�qR��>z
�5�m�p���K�i��nxpd�Ԭ׬4��l9��j�jicbf���h��=�O��&H;Sb"��f��N0]-�q̍��5fܿ(��]Z����xӱ9�Z�d�!�ۜ̉�6$������w�T�P*��vpq��H��>��.����f�ѕ�	��U�.H�u�b�&���Q�n�&S�t��jM=Jd$K4����v�y��)p*<;�������k4{�m�)�'l�I��-~J���+�4��ih#�C�٫;�r������};G9�gp���¤`�k^)�O���tX��<�mY��8(\�\?���LR��B�ʴ�c<W��x�0De������ݾX��)�us�9,G��@�;�@@�ä�5��^�w��F]"�-���*V鵚ڿ����<8��߯߼���*�h��9�u�V}�p͊��`���VL5�]�dB���b�7]��$�,
�AKt��&dP����*FЧm/��ST��.Ka�w��/�/1u���w_���`�ą�w�N�����f��Q�57��ڻ)���)�o>a�G��Q�k�%B	_�Ǉ��ࢻ<��t�!�10���I�'�I�yM2:~�X�(ݠ�'9��2�~1S��F��A ���t͝C��l�����Ѷ,��t��#8B��WF�$���%�gջ(e�	B��MBt4�(��w	�ēG���,�!7+���z���Gv�/�bz��H�ЁF� ����G�mf��OA/k~�קXg�43v���Eb���ٗ��<��pn<_��$�9�ֵ��.���{�f�QƂn*�R�j8���i�N�����o4֦ ��kc �O�W�l��֒��	��Ӏr��9�~�����S��& W��ǚ�A��3�e��T��8x��Vy����D4}hǚ��@���cp���7Z�8R��Y6��=9��!��-��#�mf�\���IQz���Y����Ӈ����kR_�><ijI��g6�@�W����'�T�<��U�>X�2���2����;��}0�_�����ge���>�o�V/p�T�������ЂK�+_���`L&c�&����A�1�'_kOf��'Uo�J+�����;�����2�nw�Oܩ\�"H����O�����B@Ĥ�
��NZ�}t��Hh(F*�'ٶ|���@T%�箛�x�����\tW�H�1�,��u����K��9�r����6qKr;}oDn_�=q�@:Q�ڢӮ@q��g������C�ϐ�l���
l�Ֆ��֙h,� ^9G	}I|�4��,3s 9�j"�z�e5����C�[�W{�n�z�J&H<\|_�z0�����}��R	m�&0`���:�:L�Fa#����w�ԋ3��"��ր?�����}�f�4�SӮ�{��.�}Z��4�M����n�UV�V�u���cy��W?����׆x&,&�'��uA�ơ�c�ׇ�ϴ1������͢��.;���:���HCFjf6Q��>]$�[S9��B��t:���ۖ2���;20�|����R3���6��K�����܎�w��c�\�i6L�>��,T-� 㮕�"�x���Fx�]����,r��p32#��)|���s�U�EӪ����(	�-g��[3��Ȱ���=�(QUr
�R����&�Z�y����I�~7�<�i�����!02�}�s�
Pu�?%�|(G����Ll��L�ko0�D�re��CN�N�)��\��l�́5��b��Oh��E�i-��3�s�$ �N��Ժ�3�0O�쾁��'�1��fܰ�>?03X�~�9��s���(D�������-��G������Xtk�p�ɠ�l0�e����e3�Qq���20�� �%��Q��>�7Y췿s���!�/������c`�*�=?lҞ��T�I�o�-&�C�W�x��|��x�w��]��2��%KQ�WⷂW(es�}n������i��Ff'L�u��t,ns.�����k�.F_dܑ�g΍���)���Ӌ<e�B�*�88�<K�JY�c3`�~�ޟ ���;���#�����Ŀ;#��<F ES�6JS�[��-VmXk���Ă����ײeLS�m�LY�g���w ,V���,\LTV�Q��5BQg�}�� �?D�&lD��N���+�=�u�7^����ˤ�-�}���<�	G��R+���T�C��=� ܚ,U)*�*<��Ly���@��\�����1�����?���8S�O]��댴\em0��+V�ox�����t
��p������GqfZ:S�v!��4�K �s��i�( L��F7�'h:h��&<>�o�T�IK�D>�cz��OvN[�D��٠��̹��V럯&<�宱H�^�B_ת���:���d���T��-J��.!U���N0��9�%N�jג�C�䆎�&����yl��v[٭���ƽ�A�@ʏ�WJ�AP�;#�H��
��yq?�ud��W�>�6yÿS��$=K�	k�8�m<�W�X��s����Qi������Gv��������~���J
��0I��c��=Ž��WQ�H����Ȏ/ղ[�MDh�κH�s�nrŽ�{���@�� fw���;py�l����x}�Nrqh��q�h@N��z�Y����4V;�.n�}1�����y����FZ*m�)��t��#��_e���%�ƨ�N�]��]�%~~��-EV��G�#
�İ���Q�r��@AO�R� �㘤�d��"���z%���{�4�jp-Z,��Rg�e0n��#�����u3����yi������ts��،R,��Y��)u0�ވmAk8d���PM�T���ׁoh�7@)�~��o��7؁w~T�2�K�)i��-�����pC���5B���Ҵ��4������D�a�m	�%���n�>�=]5Mo���t;�ldU�F^��f"մ�ˠ�i#�S�� i�B��op�s��@���k���:�΄I�5�^�<bTW�Ō4��lt��&@�F �~�,���9�=@a�n��V��:��\��a���"����n��pi2�v�F�2��`ָ����1�qi4I�:0��*����7���9���<�ԟ�z��-i����& �������t(�򄌴�����}�<o�`���>3X+�+:���XN��h��.K�3�Pc����N�gn��}���u�L����\ũ4I���p(�P�SV��m�������k��s!�\�-�����P��k�.�B��C���V��:�Vf3%E���(s��:��v�od^�f\C�9�8.���@���<��Tb׀��'��!�Qn�`�,�S x<��r�ğ�j�xz�nK,��.G�{�����T�9�ES��r�)"��/�,��v�,<�C3J{�t���-o�>L����]o)I�M�+6>� ���%'���DԳ�jϮ���K��x�kJ���P�*K�-ģ��/V|;�X�)�#��+������{�J�'7�I�r�jn��]�٩�w�#���X���BIq�"��x �#�^�����
n�ӈu�cֱo2����H}j�bq�V�ť��0s�%)*Õ�PλG��9�,�x��;S�l'/#q�a�u�����@?�C9Y%��oޖo߾-o�~� +n��P�8p�vIO��$�Xl�ۯo����Ş��є�
� F�p<2[Sm
Qm(|N�{����l���O)��e�mS9���9��*	d�nHP�iY3�J��X��bRDYԁټ��	N���ɭ����i����NMm��w,�v��1'4������-���uEM������@�4�b|Qv��rj){^; *|��1��!�z������ꬪ� V7��J���F(�[��gw�O�-�\2�f>��������g�aa���C��gTS)�}��q2�s�n�FN�a�r�*��K<t�39����f<|L������XGD��d߶7  ����/�P�\��zpr��h7�����e��s��=�F�ɏ���V�*Rrd���k>)�&�U*�?>e ��D-�t!s��16K�Z�SK>J��;^�1"e?���%?��N���N68pY��ݻo���,��O�T~����ÿ�������J�ol���N����onI�Ɨ&�\���e������/���"����=\����~u�X�4�1%�6��6į�ICn̪XU7#J_S�hC�]w�ɺ�]td�xnO,�Bvξ�����J����.�<�Y^����>-B�����r~�����)�F��6z'��/X��U
������P��-�kM�߾O&����H��cB{y�/�v��0Y��(��gp?�'��Eը^Ǜ�-�_u��̒U�0�`r��z����ό+��9,+����e�y*�n�KN�m�܈�,ｏ�i��M��PQ[����~����В�Jc(]�awE�/�IC(~���*�'��+AWgT�_��[���<u���
s�����ׄ�6�Fz�G�_��h��e]�N�֛%3�ظِ�������Tl3R4(� ;e?Rt_������<����C�ם5�8�s�S%���~[������������|^�g��2[舾�dHw _mпE �F���o�߼�*�u=d�q�������}P6�Y��x~|N�>���s�*idfE'�a�Ms��E�xEF�4n�N�Q�8�4{�:�ZNN�_1K����� ��~�M��1�ȆFi�Յ �M"~���dvK8l��k@��5�A���jDh�]��w���� ���^m���o�����-�����;#MH)�8�y�.Qj�G���K@s`�%�\��>��3��=>�G���]SN`L!_�ʟ�ڈ�k���le<��җA0O�j�%a#>�]5��t`4;�/?o\_AB��c6�Z��"膫����gz^���/b�Dއ��o�����#�U8 ���ä�8�~���i�W�mZe6a؇��}}�b���L m:�k��2�v���qCJ�!��k*��&	{�bVVM�8�\�Z���A�G�hڟ�� �`w̎Z�E�>�ca��
��%�E|P�Qs��w�8s�9j��D����m�b�D��>��A�q����.�T�;� !���Yb�8�u~�������7�Xa�P ѱd�r����y���%�?��3��j�'L�����^C����5��n���P�����&z:?e���:��4�f�C�3�`� ���cg:�m��!f���<�������@'��2>S6�ǤU���T����I's'�j���<�u��`[h�b9�T7�jp�!a�黨�bͧ��$\v�*Q�:o�F	���2DzM��.
v� �kӹ�p=��l۰M�P�������j���b<s�f|�u�*	�����C`��j���k����������8�����~4��MgƟ�G�wqy��W����_yTt�tF=玕�;���-?r��ty��*������/:���"4�������F�I�w�h:��
Ej4�mʳF.&Y0��`�Opf��φ�ۆ��͛��W_QG3�{*��(�ǒ����j*�Ρ��,�8%���b��;'y_j�4���>}ܾ~�w��>I�>�ָ�=<����`J�	n�IӇ�KW�ǫ?�̂��\X��1��@ ���,��sL�AK�)����^���z�Ce ��½����Ӣ�%�(��
;�����;N��r�8�*ԍ���"���ƷѓS��)ֶ���q�.(3�l�D�dC�+��#�}D���^�뚴��1g���G�a{Ox��|T&s �+�p5{����t��Y�����Am�u��q&�N��P�:&>K<��������J���C���Fh4u�Ŕ�m�s\��T|�6�pM�t�{w��r��=��X�����z��T�3�v8�S��8���K��)���G���~�RJ��O��v^��k��3�R2;B����%��5� ��z�p�5����x-��#^=	�Ѩ���;�t���3W���M���1�~7r|ᐉ"����{��c����V�o�2�ZS^�x��7��%?z1ne��-�}�J<���]������PO1]�@��>j�QrW1c^��蕉`ڑ'MܱD0�8�����o�F����C����`�BN,j���������>$��N�Cn�{�q;�)A~[Θ�a/�P���=Ҋ�2f0e,*:k��뜳�����/^�~Lѽ�Fu��}���;C���%S0�h���Qih��(����U��m����u� �������)������.�L�t��Kx�1	�[����^������sׅ:��b�mZS3U��Y�b_�Ȗ�V�8-��]<��<�#E�;S�E^&@l(m�6)K�Q��(��	O㙊X�w�|7�X��6]��d��X�]Wv�Ӯf�_��ͪ�����@fGMJ�S��Q�T�J� �����p���r�񲛨��a��E߭������)ѹ�-��"h h��ق)��� ��sH�1��bs���V�2�TRpk�aC��cŔV���Q��/DC����v�댷�%�����YRŏ�O͸��ۤJ!�����!�_Ra:��].�t~���<����%��nAb��rV�_c�-���.�����z�uz��lN�S�t����sj��}Nj��U�Ÿ�h�L�9�A��"HM����fx�)��	��Q��v��1#%�T(�%�\���E�|`p�窻��KdT�[첔�]��P��"�Z��#�i��E��{Uk�f���	�i�5���]:;�c?�ڴ\��x<Z����\X?v
�t��Ӎ�!��5�^�������*��?N\�)�`�Ch�l��a��?��G#��eWϛ�<�8z��)Q����gv�%ˣ5�o$����v�����KM���ؑ�)���7p�J�UGM�!�YQ,�g�g�'|G�R)��b[���Yz<'h#h\��nu|���p��G @�v�mޭ��$7��N���ٌAg{�wT)�  �8�|�F�d��ap�rd?�Oل!�Li���4qU��v\�C6ָ�l(!X"[j �����i(O/�x�BE�큀�n9qm�_V=[�O��
z���~ `��
�����0 �^��0K����0���4���􉃑�����<��Aa���wI���A�`��C(�K��ݴ����uêr���� d��S��Ug&%,�x=2;_�9�����k�e�?+���`7�B�~gP��?�QJQ��>�j���G����I!��s`��Mx��JE���?&�;����4�8��G�`�4�>Y��
[G�4�C�v���5�ڃ���P@�zT�k ->��/jҜ�%	��P������L�����
Q�\-�m�a�J��&'�Z�Z������bQ��"��5�}t
��#����b�XPq�.y��9��x^��O/^�S#J��MⷃrOLid@��)o���Ǔ��^�1SEKN�Gooz;������_���g�fIC��|0��)O]�֪���ߡ�:Ӫ���'6N�o[vv����	��Au����ߥm��l7N舕�*d9e`���H�M���l��sy��W� �p�|����G�5���±Yiǎ�L�� C�nf��kbY��E<�ʴkH��&?������^ۑ$I��9	�Y���|�=���s�av�{���d]TD�,�Y3}�E�hdeA���TEEE�I<`"����{W�)[	�p��fe\��1>Hj:	�ȡq�7���6�&��xs[5.��ʾ0�l��6��4�*�w��I��B0��0�#e�� �EQ4�D���>���~ q�AЄ�O+���^C%�����3+�R;8��$���+W���>��(j*Ji�S�F�H[���$��i�d���&#5��&��OOt�����J�I87��f}���.Ū�t���U�O����
���	��VX��j������~�瑪���T���%.:������綉����[����g��G�s�)26H(iFpCѵ�N��c���?%O����f�a��Y�.�/��Ϣ��=�A�M�^�y����y��u��!]J�GZ�Θ�hF!�{�ρ���w�i�m2\ |����]g�is����������oݳ��#�.���(�I׊�# ���`�s���	M����Q����:�Jպ1"�<�����L���x]&S��:�kř���.;��^���j�*�p�܍�P#<6��9�L)���$�4�Yt�4�:)J�g=#Af�;ds��߬�N�P+��o߄���h�n{�!�3\362�H$�u͌o�s���Ѕ���*�Z�������~��>�m�0�(�?���9�Z=w����i�E�V־f�K�`�ʣ|3���m\D��r0mJ�8a�鶄).O��'Mκ.k�P������� i5b�8/sf
�(AAA�.�'[����_�?GG�%۾z�����Jט���NǰP޲�(b2�Z��Z��%	���>�e�mWv�3�A��^�LnE]Rak�s�Į�X��3�v����S �ۥxC��cg�$�9>�P_p�B0C�A�4��)C�]?D��f6RN�=�FdT M|߇�K��LX&��:��+��I鹣u�*�e-o׺�Kut��&ˡ��gb=5Sv/�'z�T�w��W�s��{��V4�>�*(Kǐ���0��=g �
X؝�H��r��:�ߗM�֡�%*�\���_�z�����D��������~��]�;���w���C�T��~�)��ł����d�H���7�XQ��k��C:
W�x0�2��4���?�5_C��,���bX������˷m��w��#���0��_��`��}嬕��������"�I���"�X/��J��74n��[+�3�[[�a�M��'1�}tH�-�y�(*��)/A�(QR۹��+hz/�'�a ����t�n,|<U`<��M>���dJR吶�)N��$7v=e��Fz�ṑ�r��$4R�)�"���Y�9����YZ��/������~��i��c� � (�@K����3�Ev��e�����������E�$ϵ�:sn�z���d�'ݎ̓�m纫��ns�N�*;�-�.i�?e����@A�v��E��WT�Ᏻx�����Q��=��~��(2����^#W�=�9\Ʒ��A7��2U���^�w�Ux��^��	bD�=X
����
P�2��;&�29����x~���4<U���Y"*�!3�6a��h��}�r*��]�? q>aUYL֋ l����Φ��
�5��ן6����d������	L��1f�"�˺��ҷ%��E�����:ɗ��2]��s�s?��WYs�4�HwU4�6�w��"^�i4�>&H�8����L-R���#���Iʟ�S�xGe�#�43��&f�Z~N� �T�?�]���9��3@X��j�ݼ���R�R�x�˅A�WCd������uL��v �q8?�z�l���iE��?�O:i[�	��0�~Ն�^+g�q�y�|��rQ�#K�,�7i��03cp�>w�K�T�gD�s��`�i�iu7�����0��Z!�Avǥ�ݘJ;�N���n�t��M[�g8�$'dr��쁅�'4�l�;����\o�}4tx��om6�Q�:��fo~�JGS��ÊJ�3�a���p��>�L4|����6�WV�z㸓��tZ)�Rj�i�hаy��O���ǽ|x�X���*�Is�N�
�������������ĭo�o�ݟ��5�&0�F.d��g��e�ܓQ%ox[���M�	�ߚ���+V�!�%"M�|�)�fS~��0����1�b�$U�c�,W���S>DAJz��#���|�n4��㩋 �<@��S+VX�c]כNe�g�y����g���H�>d�v��&lU��zr!��z:wWU!���4=�90�)}���EҬ��/w���w��ZI*������5�c݀���ԯ<�f���UU�J	?����1�a�ǥf���u���۔�F��^т���5\�yn6��冩\����~�L��.2?sC�l*yOz�u��,c�lDU��!>SCi��T��I#\K6g�e�Z��}D ��	�
�t�E���w}�_Mi
f���l��7$v�jx���E�;56���1m:9I����V�}���\y`�~��ݖ������/��,r�nu%c�I��4�̹�J�n�H�\�_dnFw��RT��}���Q��Yu'��\�Gz��v3�!΀��j2�����?G7?�z�<l��wt</(!.q����Yt��~>�~�/Ȍ%�wo��F��>|z���pO
��}�e��ɛ�>R��!���t[t�_8�	퀟~��|�����>mY�p�2.Cfj��I�� ��ipwO �&3;�$����v�AYB�ߟ5.�L��a<`��d�k^�	|�,�JP�
�zj�Ѫ�9/� X���N
jr���:�mo���ܓ@~a�Χ�>�4AS�>+wVG�|'\��3*�K��w��.2{\S�N��� v���V���|����t4S���� ���$[�������kx�륑b�B����f��t>�A��+�V4:�9Z*Wqr֥]
)ĝ�2�AJ�ˊR��2m���27�ێ�r�$ׯB��m��n'2�ei�˲ˇ���u��f����F�*�jb�C�� ୕6����7]�x�Ncl���	�ޕ��**�Oe���P2����Q�
�r�U3|�P`Q����u:(����C�g�I�����R�Yv�(���@�_�i8Xp�M�Aĭ5+F4��I:���U�;���������Rf���80e���ݩ�3	��Ӽ�����A���xN4�v���������~�Y*� )F<�Ɇ�/~σ��E)֌�KWՒ�p��Ț ��5@��>�:���
&�t��c��qϑ��?ż?�w���*C�Y��� �{�PL)�q;;+b�E'��8:�۽���������\��OSn�N��"bd��C�F��z,���u�h�5bZ�����>��xx%�7U��b�Y=�e1�p��H�棓���U�h6�e+�j���;������gM,U���R}�����ƭR���2�Z!|�_�W]{㤼�~!Χ ���3RO��,]�����P}�o>�_gQJ\ގ��"�̥�n}�,�+�2H��0 ���#;��]Ⱦ��r�y�;��I�S~���q����l��ö��ȱܝ������_��������-t���S̶�D�x���e�����D����a�<.����>q�9><LA�U^!���e��>q#AAW?�8���_9��,#����&n�I"& �k s��v�k^�v�$�t����fU�c]O�Fp��u/û/_�D��t�l���Q�y�8{R|�Y�nZ;x��*[��sMB6��%�w��jz�U
8�?~�����;YĦ���'������`~��4��Y��+5�����LoB�� W�*Np�IJ��߄�Q��s�f'��A5��C���6��q����&�Ki�3W�Ff�s�����z�����,÷(�~��9�yW`�Y*����	H����xb��VUk��u���$:-N�,{is��g��� �C`��u��������v^}}��t���i�����^*��g^9���`0J��b��@�@�Zm�ٽ�����qm���%��v�R��L��X#���=������
Iw[f�>(J��7��r�y����t-��?�ٿ�������q+}q�8������ز����s�r�5 ��4O��b�<�/���%��%_̾Cc@��h����������c%�&Nhl���c���;lȤ�������>��
D�I����v���x�X�O�yhFV&\oi0��dY���[�U�`�d��"2w�!Sqc����=)���2�ޝ�o?�Wٺ��
ci_�XLA��o�&�:/�m�qؘ���~�g��2�@za?�FnW٪��h���^���楸d�h��R�_$��wc���X��������$�N<lb_��V1:�f��r]p��c��d8ßL;�n�jw��B�>�M�D�X*�?�����,`9^ja$꯺7�-Zj~ږ������@�'���-�f]nL�B���SdDA��eDH�5���I3؝>�*���'�_�!Q��j�BD>�J'-��M`�M�A�ԲNc(�G���顜� 5<�z�����
#��54�@Ei�I������?�������@����	S���9߿��F>��2NRL*ɞ6�lD��T��yfs
_�8x�_>�2ﰯ�t�F9渗��A
�,��%��EI��?���*��Kf���s�N�B,����߱�F�����Q��s�C���1Q��L���h@�(׮Q��g]��ڇiov�]y�U������}&[���	U�����Wr���m�n�����1 R7���+�v�eiܔ�1�3]Ū`��c�-��0{_ҋ<1,�yN��h:��t>�b�����2y���Ƹ�{��A}����h
�{u�8�i�:�}��
=�<�g���[�{[k�LB��k��j�ۃ}l2��V��j۪ +�7�^�����zţ?ID�=}���Z���n՚��&���'{�_(;��ဠ9�oِ�����p�Y�j@](���5ښ��=7��N�K�"w��83��ih5��=Cl`��&x�S�T,� ����΅�¦aa"�B�r��?����Q~���#�3&��?���N��ӝJ�O�s;�#��I����{MNu����>]ʗ�)`�о\Y`�(^��1��턗�.z��;~��~�B���
�K`��}����|�Yq�C
��!�q�B����5>72L01�R/ ����p8�s��_,Gyj�WC��`����5r����V�G�7iM�^� �wp(9��Sn]� v\G�925'9��J���fs��[��3����y|���Ý�	T���fw֪(J"����]H�R�T�����8�v�� �����3��?<�G 
r� �`�������;�#���GN�u�c�?N]v���T�m�/��Y�$��l6c����k�k�����2��v�$1%ߎ��Q_���TiT.��o���eb��5�Mp�DM��$e�
//�lV%�d�x�������q<��K:<x��
���:V�کXz��6f��<��aBaJ0[��d��((ːaOe�扌�ܫ��uCS������"��b�x�e�wЄ�]:�t8
�!4�\����(c�|�\�-�]�_]�U�����!)���=�E�/75,�vz��%1�� /&0�-[9C�s	�'�x��|�#FN�7$��|�j#�K37zm�^����1l0l�;���n���u���ρ�Rq���lҠ�k���;e���7w�|tŢ&�e'B���V���,<� ���*�C����矻,�I._�`m�r�!N��j�a5��K���;��E9�\S�|� 5Q��Lz�ES}�/�;\^�Z��hG��g��9�MoI�I�޽
����O��R�j�[��1�#��J�-^ږ��U$� �����?SK{Kx�KJ_�S��,}�8��1N�A��y��O�I��1[�O>9kK��;��5 ��&� L�󲞢���w����UD6��u�,�����D�C�����q#��B��~x`Ge	0V3J��g)�ܔ���&��`�nz\����}ϭ|O����.�9�+]1�X��@��^D�
B=���-"3�˺ُ���AW2��x(���ii�����E���8�/k\я��iv�K��r��e*)O�0wq]@$�ߛ��k!�޲J��R{�9gq<�Կ��c�lb3_<��^e���EpQ�}��;��tȍ=�I����6�����h���I!���Y��@DJ1n��D�$^�*L�1��X�]��v��#l�)�1��u�:R�֤�x��|D�(�k�)��5}��0���:�� .q|�O���j��*f���߮�op�6�d�����u�ɝ3g>9J����Õ��@�6�g��ȟ;i��1Ƿ���(�<c��%�A�k̆Ƹ-���'���X����5�=��~��tK ޼Z�5\N�"��-*�w͘�sv�q�7ŵ!�����اǓQ� @�uX�Z;�x�uK��+��$� �'����lӞ�T�y�2���sX�O�u0gP�����a����I�'}k#�X����:�n��d�ꮿmd�Y�h:��r���i��ف�@Y�/)�LݓC�"S��w����O���V/M6�d��;���~ps��JN������8�Y�@7ub{F0��E4nD�i2-��ݐ����H~4)v�hss�͉%������CX|�PBa�.�R�{T滫Mb�x.9��r�B:)yJ�Q�+B���kb��U��>�-X�����lTe�m��v��{�=�_Mi_;e�K@�xe��Dn7�pӀ��.��D+��{��r��t?��=��au� ���n���!?P��H�U�B�ˎ��E�Y����ɑ���4/���9At���U�Hi��t&���Gzm�����o����b��CRu띑��D�ׁ5�vl�[k	��x~,~tϱ!�]��U���d��9M�X!P��^e`ڏGy�Y`m �ڰ���N�wC�8��)��Z[׍Y��8L�h!����&��۽�T���v����1�	���N�A�4Y5$�g�*,kN��������<	ϔfC����A��̒]�9,���c�O����4�Fʠ�!�k�2�{�T��~4�i�*3��+kf��i�Y�Y���B�������N�9�1Xdy}�q"���SjkT��9�6�r��f�QU�xq�����L߳jܺ�e���_�������[?�d���ԔnU)_��i��%���h�����EtG8Č���z:��ۈ7V�d+�4&`����rf�5�i�;I����7~h\w�,:��q���U�x��otI���c۱sF1���xXn0�8eE���G���^�$���3�Jf�MY͵[C�=��&v?�C/`�9���¾{���l�E���f�$L��h|uူ�g�(:�p��9��թ9��w��c}ob��4���s����q'Z�-�������1\7�T���k�Y���)3�~H��,ӋԾ��S��(�1�N�R~����s��'.e��$"���I�ρ�B(���#���hN�w:%�M���U�g;ꖵ����c����g�~)�߯�z�QF��������3�mЇ-]��Fų�X��%��	ۍ�l���zm�R1�g3�!$U��˾Jا4��ϑ���b�S�)�f��*����Ds�8i}����WN�V�Vк�ʚ2e�Vc,N����}|Rs<rigNy�ԓO!n�P ��?�:��h�&5���j �ɿ_�=jr�1���Ԣ��s�L�%g�$�9);�n�0X�I��᱄��y�;�A#�&薜 �b�UË�*C<�J�'��s���m��I����-��~���~JQ���	��Z)����Մ#����{(�ј���:�["�YS���M Q5��\�fk�u����K��,~���7�3h����d����s�^��_q3sȩ>D�˜TVH����gp��� um0�R��3��+� .�q7����ϋ���զ�&L<�Z��X�p,��0/�c�ሻ���>k9O�ܪ��yni_A=\Ki�Q�+���5�q���g�g�;��#0�pR��W��l[,���\Ҏ{M YYo���z��g_�0�5��Q��e�����#.�g����f}�ƥ�5.]�$�*ߣP���c��J�ͰWL�8mY�5&��ǐ��S�N��9�"�hC=����[�7���#0��Jn�m��yf@�˝F[���E�S���Ox��	;�|�yzƻ<������"P����e�^� `�I%[	n��0!ٹ� �Q�S%�%�������Zf�����R�"])��[ m�l�=���~��(��ձ��c��*��C�kpIn�{��^��Y��>df������9��b�3�Uv�Ywj��^����OQ{<vE�&�*�\u���RXyִ��,�s<(#��(dy_<Y�,��8#�B`��}� C\�
P�H<�		e�P�z��j��)�tzIA+�ה��
~��&����A�CP?�D�Xx5m��������ϙ,�Z�W�Z"����Ƕ[UK������0���� �Iy#�Kro�cNR_�e(W��9��]���q�As�P@u���µ%R�sTzU%k[~/�hsS�{`�#ۂb�U΢�d=����
�K|������w˜�;�sd����"����Y�f�`^��/�=��E:����2.�NU���p���%��ך�#3�Qx�;Ü���'oķŭ�d]��Lu1��Dդ\�2�v��8x2�i�-�m� ����IK�ɵ�4w���R��gUV�V5�`�u�Њ�p�G�����l�X�����k.�^3���x����s��Kg�r���`�M@�N�+��+ENju٣��)]�d)2�yN�Ӳ�G0逨\�'R�0�4#Q(f��s��Y��Sy�0[3�*�I��e����/5#��"��η	U�!v��?}+�&����m��s�~��xRlRg�~��`ĲT7|�#��8Ҫӛ����SF�|Y_5Ub���!����<E������X��yMQ�g���-���"������K���Lx_)���$�x������tn6����p�Ӳ���&��	|��jY�o5t��vF�g0#�Nk�t�Y����hF�`^{�02�P��᪦����Zf���1\ K
d�1����U�,[d���}�J�`�|G�]�6.x����bD�����qp-�9{	g�Ti�!2eWf�_v���J#���3h`v;�`�=���7�k��]�Ed��2�*^����~���R�2G����+9+;F�I�Y���.V�wr��q�e�i����#����j�Qv��H�����g��NE$T��§^ι�>��a�É�T�Ⱥ�|��f1�zOy�8�7+�zo�؛��U`4����D���ƞ���n�,��l�՗I�P�!�9�q�WJ-���kD���<�T�����Sr�4i����t&�!���� ��9�����c����Z��׿� �J�5�ٌG�PJ����)t��ۣp�o�l��M��_C�Σt�@z�pσJի��3�T���L�`�x��4�����"���T&J*�1�Y!��+������jS�2U?�w����Ỹ;q���տ�����R����sL���KY^�h�\E��|6��r�*���`z��Ń!��@�&z�l�,��}�-n���6�}TD:d��FP.�Yr��,�S1Z��G�Z��l����:Q��	��,��a/w�52I���+��.�a�� �����:}
k��-����y��0��`�3>&D��^��u�Ux�l�<x}`��F�k�S������π�l�.����<�e��Ȏ�<�k�2OH�����n?׬6GD+U�[!���\�k��}��8����m������y�b~�rS�s����`�]x��9^j�`�jv�,�ܼ�� v3i�l�_`CU�b�C�=���+���?���g�����B�m��MCΰ��o��Z�����H��熒�D
�x�oZ������zs��zyvw1+�6�YaY����lr^���7e�^��?��s��OP���?~/��;�@/ �4���UF:P�g��%Fp��|�}��o����������Y��j2 �B��������VV��N'7	H����yϗ�e��i�>�L��2�o��:D�b6X�e>Z*Ek�S�3:�b`��2����E�2�]��[e��Xr�[��PX�����Sv1A$�mdj��_2pO�9�$�F�i�H��m,�=�k� =`հ$b��5�L8c���H��#������/����1?w	M�_� �ۥ_t��y��w���:#5��b����Ig�HE�Ǫ������ϩM�8��Χd��\,�唋�V
���3�Lk��U��Dpnn\Xa�x)Z������)�i��<��� bG�=p$��4_���%-��x�]./1{��K<������TTHoE7�#d��A�u���6,dʰ�L��6�_�=�}��1g�B�˚�
���ݹ@�p�t�C��8H�U�l�Χ����i˸?��,!ܶ����_~�F�R.�w]�bZ���u�EN���>��������My�?n%p�%����9�`~�B� �	Y������C�-Hu�,���!���ch����;��C��޴��TY���Ҽ��������A7H�
�YҒd�@��f��.�1���2�^�~�6�ٴjEj&��-Q�+;[��XK�0y5�Maz���{R&��u�'�G%;l���KX`�#���T���G$��)��2���u���)��]�;��ܴ�. .(o��B+m�A��lJ��p\x�]/C��+�#�0^���I5����/<7��Fm�����-s;�V��=�*P��%�e�� b�\�_ҵ�����&n8Ɖ!�.������l9��@*�(��zg������@
�P4�5�6��@ ��P�0��)�it+w�@�����@�,��ᰋ���D�}z��|���x��c�����P
N�݀	bAl7~ �|�Hs� �Tt����Rg�c�@�Yٛ�2g�J���L	bDHQ޸���m�T�<w��9�<G0mC�]��q����u�>K\L�HF�v+^<S@��s�y�OUd�?|�v�0ᩤ�?������~;T�	�s�V�C����1�&ͱ���C���H�.1�ET!|�@�����vZ��ԭ骡�[�﬍���cC��qX�w�D�hL�#�O	T�'��I�Kxl:X���˵	�Pe]�po�F�k�p ͉�yJ�'])I�+������xO���)�E��I�N��Y�7W�h
_��}���i�����v��#���%m�9�A�r�d���ҹ6��y�"�ax�mٰM�b(�/,��f��?���0�kd���z��7W1h��k3 ��vpd�ù��7�0����Z_g���.��T=�։�f�w`q!~ S��!���ٮWEsJ�%��\�q���i�`�/6A7�QR|���ȓ���Jz�ة?D����Q���:
��?A:��q_���Hˢ@z��Yi4��]���=�xB{�3K$���ve{?�بo�Ǜf��u��=���Kd��J�|+{�E��#2>*4f#�T.P���_b�g�"��{�-�sN���������ݛ���o?�_~�%����e�J��P,O�w?lY�����e����\�,tQ����=3�`G�i�NT����ɡ��Ʀ8��hL�M���
Ń!��P�
:�JM���|��lh��e��p�ʢ�cj>*��tU��NR������I�W�Ʃ�d�!9��f��A���r������:������MG\�@�U��.�*7
|�\f���?G �����~�C5A�_� .s��1�Y��gZU̪����tFe�L�u�r��1W
��1,���K���N������
����2/�V�k�֜����fiW�&�_RN"r+���a��1�׾�!�E��Z��^��3�}9t{��Z``k M�9ۢ��O�8V��U2E$�/���B�׌�)1��0#f{�R�aVJ��52�lܲ�~.(�q���Nwߨ)7Qd#���ۅT��}n(��E	�R�����A���AGEَ)�>����v���b�=�0q�0��� ��rB�+y¸.���ٰ�#�)�ˋ��z.��3s��Ɇ�Y`*D&SzQ�(��Lf�i��wrKg�œIb�>2���R��@����IsE��Z��@�a��ö�ͅo��|����K�`#X*�t� sO1ߴ�f��p�C�U�u2W:O��S�����t��X�a6�6�+
�%���T9ᮻ�T� ��z��\^����������I�li�.m��t%7o�ʼ�ғ�n�Ĭ�i��ÈC�R2��L��y~1�YH���9�:�}��ݫ����Xitb����F mh"q=�������G�O�*�щ�'�a�r�Ɩ:���B*�G:c�\SkjN�,!���x�#��	wՄIX�vUs�+]^`��Q�~�=�Xt��XA�u)��ꋄhDG�� ���m�~ز�-#3�ֶ��M4Gc����\īj	���M���[C� �
���We�3g����N^Q�p�������|Z@d76���S]�6.z�K
;�ň#���~W<�v����I4�7�����϶rt�끳X7A���jd���SS+�m��I���1�PWXgi��Nxݕ�ƺ�94�w+6�V!hS���8k�+@`�UM�����'���*z2�)6�����u�N&����Fgw4q�i��!��|����LV3ȯ�&�Q�<��٢�p��ݨ�A�h�}"˽�� I��\Y&�]V�QJ���>zO�XhV�5������5�vm|�[��E}�E�6����B$�G�[�4��b��j'��8*�N��Ȧ�7?K����+x�m8w�cZc�B�H̕�����6A�X�)�����<
]>��	Z�[ E0�.���!�,�ycdn{?w�&w�_���� ��1�����{��	��;Z#pw���#���$>�z�\�(E�l!��e��vˊ���+
,kB�B"��]4x�����J�8��LꤞԵ��SBϪ]1?�P��I4tǭO���1��K8l��$}Nz�(^���E^�]�_�*́���[
N;��jvZ�����l��/��θ� N1ɷ��j�ʪ��fk��R�JMO�PW�ig��)cx:3�`D�F�d�%��W�=����Ƭ���w�|XG"�4_�o+�5��1L�8���J���8C��OXo�zp4�	�WN�圿iJR	{�g`A4)�w�A�1/��z5�sDc���
k6�U�n�j���&�5���������˟|ys�jX�@3����M��]'��I�6D	��ڵw�� P�m�ՙ�/���9D@��������DYLV�ܮ�0���AW7�73R
#�lt�h��ib-!)�$i=d��fM~��-�~��j��l�>���.&x���(�	�#>P����ޅ�ɞ�Y�@|X|y��ml�"C�6	^):S�mُ���y��3�}jL���A�2$_��C �+<p8a�6 x1l�����+��2�8�Tn�t���ͅ,���*��r�
�;���#-]KM���Oڮ?I�م����,���\�� 9�o���0�f�v��k�J�,�Kt�cd��?��~��?�Ϳ�����2���m�Z���@�4JcV@\c��G9=�W�_q����v�qo\e�y��t3���_~�6�ω�����x*qQ�{�‥"�Kz���A��;�WU0\�)���e�zE�G�A �)�gS�BY�ĞZwU�|�/�VFʘK�`̕�t���.[eD�$ �
�������K��BG'��,s&=��m�Zb�v��CʾA�l�EJ�1�h��K>��W��=?��̿q� �/W�c��w�52�T��>Pc�� t�S�+o\Y�geūI͐^J:� z��\���2L���#�(?&އ��-+-�1A���E�C� =JY@N���z%T�>��zK{���H�*�M�`V�j̢�s���7o�^� �.�n�e.Ehv
���(�����s����2~��46#Z�.Ӌf�`[��y(�Fv'��֠5I�)���b�jt��e|�Q�Z�۔����r1��)��`?�*X��:k�n��y���7��ؽeC!hc�Ú��G಺�ؽP�p�Y1X�&���>C�Mq��*uR�=���U��׳��rjhqe*�m˜ڧK{��3�d�5�5����i���W���IG?��Z��	���`��y� ϟ��lS�^s�XLෝϧb)��S���QX+��2s�\��i���l�9��R�Y��T�&40�G�B?n��xZ�r��l��wq�z��,�R��h������j��C@|�]r��d�ұ�|��$e��.��cjf�>�V�LO*���p��x�Yc��̎Q����O[F�Kd|o� \�1��i�|�{�U��4���NЕ  0��)P��&g��@yﲊ���NG��AΘ��!v-��)��,XDgb��x��t���¬L�fUvJ��p���;؍'P���U���zI�	��!`��5�����v���xp��=�E�!hz���}J��}x|E�U�c�j;�%)�	m�}�$�ۭY�ǜ/
�s�?~.2������+(a��P0c[v�7l��&@�=�(ziӆ��X���?���U#�[��EW|N��������6|��𙥾*�K>�SMi���(܀���}�~��������,|:�cf0|m�\c\����[������1��X�A�X��腦X�^n����D
��pнfnxt;�[��[O���zI��X�jF�S����MbOuV��$�=�c�����<����H��D�A)�	��i�OR!��l&������
�������l?�p�:#�,p{�B1���sՠ�uh�0��*���:��cl%�����^�Hyd�ߘ�57w84ws6D�Vc&(��6#u�R��,O�u]m�}�8X��նoH)�@�������ޕJk"}M��'���D��"E��]^���n��>�oX�7|��u#KPe�(���=M �&�vs��~%��r���*9�Y*`F�{�Ā���wx.��e��<���[z�U3� 1���{��FL��t��x�T�p�}�`�ç�U���k�K(����)e��VP�2Ҹ�-F�OZ����en��'v���� �R�ڣ�5/��,�T�(;�2w�L��g������ ZJ��D�g�Kӫ�6���]I^!3��|	��Ҙ���$x�6��8u�{.#0� ̅�z�]��ϫ$�z
���-�#r��Y��펢��j+��d�c>�'�l2I���nh2ɾA�x�=qo~хSW��'��%�Ʒ*�)M�&����8��"��#���M�kۘ���(�e�:�du�j<6���Q��;���+u�M��x���4�ډ�1g�}k�W	�G��i�9�tc��^��k�V��?S�}�ܜ��v�,=�f͢���A�����и�)D�9'L��(ɯ6���Ӑ6-~�kI��k�t+696�srO�P5�������y���}72������>_�Z����:���o2T<�4�j4����W��(����F���N���t�w������&>\ȬM	�{�ڮ�&5� ;i҂3�T��ԅ6�R���R�r6�SBh8}~�T%� ���&::��g�z��(�I�>�Ɉ���I���.�AC�^P#=d��fC	����2�9f����1�Ȝ�F�}�~�~+��`��0]>�� ���0"}��`2����niқt�_Euri�6��g�&NI⦏=絙� P����g��g��+�r�c�VI�{�����${����(�W���C3�)�;�7c`��'�R�}b�Weie]�˼�`p�fT?��l��t洔U��
8g8
&��z�ϟ3{���5��@���;]KŒ����S5{?P$bax����~���N���������ON�{���{+��>�7Δ#k�R������MFm�V�V�شDd���e����V۠�J��y[�4[�M"o�B�����3F~M�8]��������ec7�7ʬc����@�M�g��4ik��3�7>���2q�љ2@�,�9�PV+�W��+�6?o6Ƀ6�?� �#�����$lt��;w��r�D����kE���<R�=����i�BzpL�&ş�ՙ|���^�ԥ�E>Ձ 6V(m���/P�~����S!��}��{�]�8�	%�[G\Ϡ�|�Xln��}qx����0�s���kmcH��9������F8�>,>/"��^N��)�.���[���=�\~�����������r͌�M�
b�v�C��(���s�@��I��rƾh���P�M�Q���ߞ�*}'�0�Z��uκ\�H�b,��o��rfz��@Z�+��M�����^�,����� �Iez�x�c\�Y����I{Sr�C�{6Ogz7��p6j?0c�9N�} �c�#�,�!^�ą����4?�W�6��F�|��5lW��>��O�m�&�����Z�(L ��(�:;)�{� d���ɻ��_3Rlk~" b
�⹫�^Z�ūʒݼ�����h�t�I�=��[I� ���?�?��#�L��x7�{/�4���[q<ǻw�#3���c�72N�f���;��E �&��N�����H��(���f&Vf6���� �&�_�a@� ����X�x�UR�k����1M�O�w��E{���AY��X��H�tFc\�L�
`�|�/l�D6�����#��e�{�J� $����ֻ�V������5����#�c����Լ`�����ß'��}1F�k��x��9$�.����ɰ-v�1I��#���l	��_<>ݪ�R���5��2�D���S7� e�O���1�cik<��`zS��ͼ�Y��V��i9��y�Q}�����u����A����!�:����TJ����;X�`�`���T%*�G������2Rܨ�@qڮ+2p�h����ė��i�9(jDm���$	��z &��ɬ�N�Bo��t�Su������5קYybrt��U�c�:�i|T�+*˧�'(�o�<mCa��e���M)��4��K��D�,<�kʷiA]m���MA������<jgB��˹|��$�EߝP^
C���yxf����>o�������~8vnω�?-��B�g��Bpz����-?jы���_g�Y�w�}n$d�>��Ŋ���w���҆��o���p"��p�M6�e4�J����ް��p&����0�.�� �!6+��(�l[�,�5Fj��~�.���B;�(j�$i<�Yp�!��U<s�:Ġ��Ȑ�|��@{���(�=f��e�d����ʎ�8h(U	3�h���2�)�B|�AS�c~�M�H{`XSɸ!��ԫ�)D��,v����q?�*{��>�M��'�ph@�|�U���V6��d���C1�k��s]^��7]�t�����K�iy�����A`ۂfH}�l�AsIV�{��-�zۤ+�~[��d,^oy�������%��7�sP�E3�l�v�I��*)R�C��\lz�����&�<C�2F�w̎߼��?[jYh�jp�ԙ!:Ѝ�͠[�lΙm�/�{�N��DЬ����)4�"d���O���R�A�I�7u	��Gᰩ*#z��N`K[f6�.45X�0a�����x�����%2z�&L1�����놛�v_�|9��}���u�A	v�G�3����W~�V�$�3�44�[�]�� ���u�Mm�A!6���5>'�~�u�2��^�b=Q���;&��EJ�n !��(�q��c��`��t?�z|1X�n�U��t�<�4N⸛q�	u��-�2e��J��c �Ѹa��tE��㬾3�Vr~�O�f�X]7ϱ�^�YF[�p���c�\j ��"&dz�&����.|ä��L�?�J��@�u��sOYd��V�/�����&���"k��iT��ƫƓcnU�#�\�6�}T��7X+�7��n5=��䦄�y;�M�݋0�����$�j�ƓLݘ���'{)�1�B<�����=��O_e�s4Xp�� 7=�ٲtuD���w[���w�>�������#�g� ��ec�(_pS��=AdDc�1'�$fM?��d�Yo" 2���(j��lK�y�5��Ev''�hF���^D�:���8��.I��?=��T��Y��(pL�0�B�]� μ�W�����'/3��v0���Қ�sQ���,~��2R��&��9���(��4��[E�����?g0x����Q�0r�	��#�x�(��َ�9>R�b�^�y�M�������+krp��Yރ �/}m���}`�P��3�v�W1��gg�n&��~"������5fK��A{�\��q�}��	#��/����pd�q�b�s�����ӑ-����+��(m͗!V�%�:�XL�D�oe����w0]o�O%#��S���%�F�_[��v�}��S��h:���Uz8		6���҂�]��(nDJsb��ǔ��@<�Z�ܺЏ@��'����]�����6����-��)+]���;�?F�>t�*� ��nv'���5������Q�13��9W����#{��f)X��)P�M�R'n���Z�%�O��wH�K<g��gȡ�B�#8(�c"K����8f�Oa=��q�{\�=K�c=(4�JW�%J�#U��RWao�*4|͹x�O$���^-���g�FYflN[֖B5��4S�%���������j���ԤX��x���R�d!�P2�C;��� ��u3�{Ҹ�����C��%�E�ks��Y�g���D[T�sW)���D�b#��L��t��j�y+�R��?G\��V��?{k���qX/�8���ZI[b��?7���0�M��=�.K��{�l�Q^0N�-q5�DIe�j�� Y��J�^s��D���S#N�AΘ8��d<�}����փ,%&iO�?�����=K<!T��q� ��)��>:܀�ep�2k����������D`�u<_�jw$�u`�猦�0#���}F`3�{��b+cQ�T�D��ƪ�m;D�4���@.��9*K
{<�i9+��m|6b��j��u�)�U�U��D��,1�)N��i��y:�s��if�m�e�	�wr�)�0��ɑ�R���Ig[WPI���[+<ί��(1;rG��t�<�ʤ1�w=��>f��g�"�{]q�A�@�lg�#ѽL%bf�i1+���O}бVA�},��U�ö�x���"��]h����E�4JF�G�8���Q�&�D�rM�c4L1H���
m5�Ӻ�=`�e_
E.�Ӥ��P'O�\���76����M)[�í8�/6�l�3u�r]�Xmi�}�zj�6�+�,g�8�������5�p֚�n��Vw��CҢZ��^��|oƷ�����5d�A�lt������
����hm��W�(N��7ǜ@��)������C|��x�V��<|I��U��ڭ�y8؟���h]�D��â*����Fm�^K�XS/I:M�DǛs�g��Ĩh�3)� �x�p�:����P~`�68��p�ʪMx�cm�w޽{G�Y��˒���׫�)C���
������T�Z�":�J�t��=џ`p�ش�@K�>�G�{y�/�&��M�"�j��l�����2k�]�ʒ~(Ց��Cf~}��a"\v�븫��y�e2�V^�5i��`�ǿ?=���l�E�u��\�����V��� �aٙӄ�.>/ /04޿�7Ɵ�NZ�Cb�d+�%&�rm���}��-��L�����x'�F�`BuK�sHpc�*I����$̜X|��.�J����	�\�Wͦ�+�R�,cl&��9�T�{�]4��YVtn ��h,.��f �w��PZV/�d}���A��5�N ��ǔ���VѶڒ0*�`򶅳�@G�3�o�f�L�"L�DAiBz0��L0U��%��x�xmtÂw��H�e�4E��92\���#^�\)&	6�9��s���v��6����;��%q֮���}�um�Q�Ly�V^ e
4\�OŘ�x�_��	�� 1p�L�2�|1������g�M�M ��X�� \��/OdMi�]�����U�"��ԎY}s�ǽÅ�ld��������;L�8� ��f��Z1m�;ƚg��L�YR�U��������x���F��YP��Bf��	���y��������`I]��z�fX��STd�ځ"�!�A��=�q?2��z��9��àY���+�J�E��ۯ�T��+��� )�=G�A�K�Qp�ȸ%�"|���k�\n����S����zE����L��͊J�qiB��|ب���<�������/7�vX��d>��������w����fn`�����։὘�KU%|]eÁ���"�C ozmP9�x<�x��q��~�L�T�َQ��I�f��}����SLو�~�Rlv�=��猪C�Z�L�a��l���� ��� �k*���P�S�"���u�������%�c/.&����>�>*Z��ucJ��BWt��!���:��[��b�6�����q��]/�!)���2{�	��~����,l,�+�QEM��`����V��\�szoF��k�5M�MB���# Ws�f��C8�	B�r�xf@EjL�#)��a��������U�ͨ��`��p�p�0��'��R4n_(�XJ��1���L�� \��I����IpCi�* 1��^$\�mV�n.*���賒��u�Ʌ��+�>T"���}�D�#��۰^K��0��SZ7a4���շ���?�*,��fM��s���	a���b	���F~���>��N��]i���]���T;粖<��^�Bn!6jb�����-����tb)l	�(w��G�*m�ÉO���8����{l�]�_�ŤqB<_t��C%oG U�0���c��{������6�'ܼ\�1yt>i��}-��ذmS���Q���i�V�|U���S�)���&��jD:S25+��+E���!�V:�J��R��m�4�����F3)�OTosʌe"�5��'��4�vV�
�=L;e�+���}<al���~�C�	���"p�3-5��>h?$|��۟NɅ�ʭ���x��eפ�]������t+P ݿ�%ۃ�iנ��AA�JU�m0��J�p �p+�VȹO�P�{��[��H \c���}�;M�տ��d�?e�m*����G�V#�)�o���#c\��}�r���Ԅ�z��<06�<e2j�mN܋��wS~��@c9f���FV�$�v�ϣ�)O���\�O��1�}�H��`LC ����v[��.F�{��-!��[���d.	E��!���K<�.�C�ɰ���h)�^Ʊ��鿡?e`Rv��=��x��q���{�ciu8fi��XZE_+/���Iݜ�����2DI}U���.e��G  �N�����,*1�k���BZ�HN�&�` ���w>N����pH�典�ul�&s%����1_<0<�M��L̎�����Oze)#�ӟ��#���؈�c��a���>���t+X�����%���bkl���ݒT����;pƞiF���}��V�y���x���up}����+�~�������^���uS�n�k��Kl��س�J��������^�������N�Q����zpz"�;Sd��X�N`���������h��hS�XZ��6+]o���l��'����v���X<sݐn��R�O&���ߤ�Ku�n�3 ���k>������	��%��i��z���S}lbA�yL�G��q���ze�?1��*�����b�\���Z��7���H�u�ϦHj�~K6E��̛j-�]Ԥ��>cJ�����w����oݨ%Oxz3I�|�*d!��n�{/���~��FoW�W6<	�j�!��]�Փ��_n4Fv�W�ǇIL%�����b!�J;�D����L��ǽ�w�U���FsBTQ�`���˥w�P�Cs�y��\}ש�P��RN.�S�D�F}��	�8�4�bv��y(�	��'�	5�9�eC�O8-�$���wM�hYd��=d(ёǥ}ߛO��)��o_ߢ4k�\��U�kڃ]x>��i{>~4N�8&��S_��#�8��T�Ab�)����SG.�S��1վd7�⯵���`$���a񺝞ٵ�c����k"��3�[}=_�]���c�rO�YsP0���(N�>��3+���)���ՉY![�L|��{�c�Z ;�0K��o|lR9��T�k�μ:׽�H͍�P�!�q��|R���=�؝4�p��El����x>���C�büX��㺄p7�IL��sC�6�12#W 9�L_o���z���w���cB>��&�����F���[�6��"��z����O}�Z�b��2֋��yp7zo̮��z_�ه�P�L.�vX--J��E��@�a����3���m�s�*���5ýw��d�ě�A%��*.ܿ�=�
���jư��ʣhm��KMZ`&Zo���@g��.��}�=37��U�>sғI�)�����Yw�������^�3�֩��5���f��U�������im�'��=	�*9�B?���E�9�pM�]��_���bFAw��.@y�����ǆ���v����-4�H8�F��(�]$��xlԧ��T>���I��X��4�X��{*O"n_�^��sl2��¾�6����Z���MS,ED����ݨ`��B1�O"���QSC�KC��`�w��I-ߖf�kk�&��@5��Ȟ���X
�/�&�8r���l�x�t΃��1�7_A���s;��1S퇍�C��ȵ��F��B1q[MҸ�3����=-Ό�!I��D%�zP�}��Mڱ��w/GL����F�+'	gB�SrINE36Nو:����d��'m�&X~�?<�]z�_�lk������P� &�kA
R�?
��=�4��	���j����h����8��_Ͷ'�4�k���I��8�R����S�L�tU������kM3~�4(��d��v$������7��T�6�.�=&'P���{��E�H�@�Ы<��~�,g��A�29-.�=͑	�cX��z��]�4:0~���~+��Q���	SG�����^i|��7rU������9S�N�0S̔�45���;���.<qcQ�'r��΍�K��԰��zV�������*��Z�u�e��Mðy6w$Y�?7I'�n�A�������E�x��}p;�l�ϋ�x��Ld���� �{F� ��O�ʯ��z����G��`�� lr�{Џ�	7��K�ӎ��02������$]/t��{�֏]Ј��M�.���D3� �D�@�.�W�ŀƔ��*���{���5���Уows͜i1���ݮ�)JY~���6�)��/̸1��@2!�W;ER�hD�lՐS�ɡ�&L�j���Q*D��C�y��,�кj,���G�!XK����51m�(�(j?e��� ����W�}m���JqbJ�S٥d�R��/^�甓:a{���s��n�#d!nE�ĩ�]��B�
\/LT�cɮ������>���Y��{�H�pZ���h��f���=nA��1�v�_b�b������GPy�n����PUq���Vd�x�!tX��L/=4=���rJ~溊:ӑ�o^WY�z?Un7��z�An�K��>G����Ex;�Н�E	8�&��s��~cנ/lЃ	��k��;���=6�:xO��~/�ZX��8���m��SfTlz����$[��]�2tj���j��v(�w�^8������6�#�&��t�Q�����>.%�,"NZ��!�Ϩzt�^���\Z��K&nf�B�0ɔ㥄�(ޣ���$���"L����P��8��<t(��J0,�ܶ?��;��A�3��59�.ߣ1�����Y�$B��.qO�ڥK���Y�7�E�3V��/�N[S�ȁإy���&��Z~ ��f�{3�c��� M�pw�n���ȸ:�J���|�~q��^�װ'�PkQG7��;y���t"��q.Ҹ�p�02��  ��IDAT���~ FFX�v�Tו�N���;e3�SG�Z���cz$�B��!H�g����c�
6Ps���!D�\\��!�҇�o�,&I�ɻ�tE.*/[К̄!����	(�k��&��ǃ����H3��;݇��.�a��y,�?������"VMH�����MIT���CmԤMĶ�Tx���m����௎
��s�K
���cN���}��=���� ��C��cα3�Y��N$^Y��\c�{��`Q��9��5fs���!JT�d7|y�߂!� T���?	V"�f5�����7����"���˥����B�9��y���$�N�w{Q��4�R}x���A+*��q�s��{��1�<���R���^����9Ox��P�L>r4� Q����.��[+;3n�κ�3G�C�F�"yE�}��U�WEV	m�.�u�E�H}��:�6Ğ�^���ʭ������I�h:��H-�onr<,l3��̖%U�������ę3构q l��,��j��h%��M7_`=�W������	�Q@f����{FFzO��I�2Ә��2Q�:���s��#����h=����O:j��I���Z�z��m�����>K3S:�>8��e��G�#�
!�z7�[�o�k������P�rז�[R ��}��I��|���U�Yd�[���w������ ���6$����ӏ��[Ъ�������ߛ*"�"sX�EYG:On�E�郦�P"V�0x��5���~���}��W������C�0tQ�XY���g�������S�%���;����iԗXK����=���oNuTREfR@ΰ�����A�8��^B�L����R8��	���5����a~Z��>�8��Y�(.RI"G{[�{R�&{X�BV�=��4ޖ�E�y�];fasO��&��x�>o�<�2�ه����2�{�{�V�%�H'eA{�%��}��8�q}���=�|@��}�עnh��T/WfU�z��d]k��R���3�I�ϏN�1u���N`���I�/�$�v}�N������D�>�s�+ �&�~T�PܽA�=.��k�٘S4��jDP���.�%P��k��Ut�,q��I�ӹ��@�Q�:��	3��v'JLbq:ÇI@���xe��e����q��C�s�-o+�ʤ�[���.�N������Tӿ��������Z������n"~�*(�w�O7D�� ��{��*�%No"���=ߕ�=6�$^�E�����t��ڮc�{�m= s�񅪨nd2A��~�&]%{��l"�V����%����sm��n%]���}9���=TA���7�j���٢�O��-R���_�4p�y��d�t���0XH�S��.<3�⾆�����ہ_�e�y۠{�}Ϸ��{t�E�����}�����GZ���Q��0X���o ��A�7C{�J�]E"?�Bj��S�W{�JИVMU��Ҁ���Y`��)U�]��;Z�h,!��Nz�̢Q�# X��ٹ'u���\c/<U�;�j�A3�^b<�c��ox!�:p����C��exo,��d><��&s��q�T��<	�%c`�bF gss��Z)�زD�ObN���"�R�����������Yq?�����Ӏ޼݂�{*�G�f�M���,nB��u8�bY|/��1^g^���B�`�*F'��-����e�O�p䵛d�r���$��#��F\G)���-N4���T�9��F��t�s��u�N�ֶ�4����y,���U]��٤�8�EzH	�3�_������3��R�I�*%��"k�~�����g��n��X�����OټTCj/�6���$7rsŔ���P����uyн�i����6o�_��W_U�$�u�ɛ/�BϜȥ�x9�4�"gP�E���9�(&^�}�t�W iZ��ɴ�]�ى�dUn�=��d̘JD#(=W�%m2�Ȑ�ϋ�86�8�P�)�e�ۜ:�T~�2�ԝO4?l��v��3 �������V�q �&-eI�ҳ�����ۛ��En��PG1��F մ�ˇ-�~��r�5�(�� Ư�&e�Ĥ�!��xMd�?��c\���-�|8f�&D-�C�r�zpg����ChGqQ���Y4(�Ϗ��A��Pħϟ4Eӑ�V�214�{e-�i�Sgp�B]Kt_~��i8,�`�/�=/��ܐ�i����UE6�ʲ�'>��k�6BpY��"G�7Ҹ�J�oS��ڰ^3a�	I5���iQ.���M|�*����9q3^��7�ii�`,\�^|��s�}�7T&�z�,�j��6�v�bĚ��n�o��Ϥ�V�
���3ES�*�%gS��_ߦ?��n�Hk��^�a�8*�A<��jx���>����z�����7N�����c�1|w��g�?W�,��]3�iI�kv��s&�_�9��~؉- ��xϡ���T;/��Ӑ�� �$�ǝbd��V���<�	O�!���<R6S��GP�Pj�M^�bAc|ũ�]%�!�^�On�I~���G��)���1K F��a��A��R���:6EEH���o?�����X�K����U<�l����{�&p�J�IG� :������!��K�j�Aɕ�9ѡ+-C=T���{m����e|���@�F��2�r�\��Gubj4��M)b8-tg�C�/�e~(��]rH[��6#]$'�*#�M�gV�I���s�X*�������+�^JWkm�����=�4WP�L4�Yq|�~m���1��4�U����C�7���&!�����+�L\kp)h������H�|�_%�Miπ�㆒�ã�\�p�`����Ė��
G�J��/x�4���ο�[����2�w�⟕��4�i^�q[h�eq�X���x��58~^��T=	e�tOh�@�C�ng��Η>()y����3O0�Ud���:������e˴h�6��Q8g�Kn.�}�Ic![���p��I��t:�[Ui̱��Eb���[�;���6��� �`^��^�I� �_:v�*��r�'����M����
�p8_��V��wR�Bf��X���h6����Uv��<�,�jP۳j�I��SW]�E2u���Uk^�c�>X�x�ƽ�6�w�d/�z(��f�;�*�3�z����t���n�P������̀��4V&N2H�"q�t�-D$�^����V�y Q�/�jp̢3�}�8ܤ�`�Ι(t'"�b�A5�=Uyм.k6jo�A�[m��0�+p%��=�:��Ԡ�5�a�뫔���W�M��^��&�T�kv���BI���d�K� ��˳�O�)o���)MB��W�';��AYj�u]��.��@-���ށt]S���A�3=Ɔ@���~��c�l�@|~�8QF8dp�_�Ƃ��,�Nq���1� ��\�������9z��39Eǒg��lA�[��M�Ͽ���q�\���XRpj���N���eI<u@�#kj�PA�o诵$�:9�ީiP���tj/�"瓲l����Fr�].]]P[F��4�Ϛ����u��^�f��$/rugP�'^'XԔ���8lp$�B1�}6��3���v
�_70�&��<�r,v.g^MTc�8rdp�5��qe�,7�_X����b���@�l�(�����S+SG.nm��s�F��D|v�K�)�n/4����g��S
�X]�M�j���f����n��hN�9�Vշe�dfT㭗O�cI����J����H[�������Qݔ�]��6��+>�N�}��n��k�d�^�#�;�c��[��cS��$��f�{X,{Uhշz�o��T���H|�����_"=�-F����^�T�3R�,Ъ�>@�	�� �AJ@�� �\В%���� ���݋��� M	���ৗ��g�W���xݾ	�4�õl9y<)^B	=����H�3X�i���@�]\+o��)N�I\/��u`������膚i���j��޽��#���'��d��.Ӿ��KþډSP��Ģ��U�t��-Ɨ�����L��ɲ�F���T���mv %s���� �.P�LU�=y�]C�p�T/4��P�1!�� ���4����w��^�-�_2<f�J�p���&}�e�T��z ,��:��z�m�Z�a��/F����F���x����1�s���k���Ag���gcL1ǉZ�ދ�l^sv�o2�.$���8�5����7=�����Ϛ���Ж�U��H@w �~<.�B��V��͂䉸�\p�:~�.fQyj��O�X���t���o�z� 4�� ���ł&�@����Ʃ�U�-�1g���G�����1��t��F״�'8J>7i>�Qx|$Q�J�K��9�l�PK�0�&Jh��߹�n���Xx.˝Ӵ�&���gE B%
Y[���'2�7o��T�DiR 7U3��J<�����*�uo�'�3��qXj���)2��uv�=�rqW�b��i�X�\	%7����a�����)�˕�YA5<b�?��E>�����0b<�S�ڎ��j�QKYV;Q���(kn��X���9H�.���"�Y��kЯ�A�^2uA�C�W��
��!�f@$U	���$�x��vKY�ػkr8����鑭�<������=�o�T�J�&����u¹6��\�R��f��?��&ʋ�S��^+�pA0Zf��5������R�%��x�+4����2`䥃��&�_�6���<Ź�i�0�_wM9��7 ����b�rOy�����/�)���ܘ�5���sR��Φ��Ά�AԜ��P1,opv!r1����R��0km��(/K#d����=D	�&��&>_l��������xN+�L�|�Y�r����m5�[t`	� ������O?���xt�q�;;�I��~�F܏?�T~��/�V6�>R��|f�EY6�>������t�z��z����u��]�Oݽ�R~�2E����Z ���K�l�Qٰ�I�y�����a`��`�Rv�����:�Y#�9��_5�i>�${*�K���ƽ}�was���s�У�YMމ}�5��lYtߨ=��F��lχ×�V<�Q�=�Z�=�)�@C%L�IQ4?ڇT)�w~{ 2�f��{n.����WM~|q�켴)�_}��͎��jm����\�Γ�TVU���R{�I����2=�7���h2'E�R���eZ'�[6�v���3�K�Y��˩ ��^Ԅ��F��@��P]
����m����`����@ ş#� �n���E�n�3�<�s����vBʥ�ׯ��UZݺT�j����%������=]��>�5dSg���Ɵ��v"����O��H$~���K���#����В�8�E#EUu��@S,�����I�wI��zD�H����<"{��n���K��pannC��Q3�c�/�M��y���쭾E�j���X��書�����FLCJJ\���.�P����l؎F� Cܫ���y�ۉF�s���p9�[���dw��bMN��]��c��T�)(Z���)Y������0�{W�ik�Wһ�"��b׫*��"J�)Ӷ<U֜��d��Q�:�����'��;R{8�%g�s(�&�s{^$�s�^ԁ��:���*_8�{�:�n2sk�!���:���43*d���{-�b&�']���X�Mvz�m�h�.x�4����H'5~�Pە�0��5����}����{�,p�~�1���\/�OU�Sx[��U��#��g�#ɓq�g!p���dMuEq̅����x��q;����q�G�tU��Pz�CR<����m1"2rj��:+�ł\�j�ԩQ����ny���Ƒ�!��:kR��BMI��IVG_��^^�z3��Q��|���1.�_�����.���x�T�Rn�&-����M�B��Ïq��Ui*'b��\�������Q!�K���E�qрE��*Jk���%��c��v�Y��0w�E4y�b&�bU��¸�[�+�긝���E>��2��ܜ��
���2�����:�bFض�NGr�q���M�[$HRD���C�ȣ���q*^1
n�>�ױ),0��~Q����z.�E �L�[g߄Ae3öWz�}N菮��Ҭ iN�a)��ئ:(��AT�J��ƞSF}.%����I��1yY�l��K�(����y���V���g)-�K����>�
'u�w��C<�&�xB%���q�.�M��rC�ի��ȬHx,DC��8=&���M�M���(���2�h�,g�;�⨅��]yI���{�W?蘙F��#2Hsb
�nc�RἚX����|�b�$�D�����������C�E�.�V���#���=C��2h�OԽ�� ��!<s:��wG>�ė#mq~3��%}B5!_�D�tg����7۽��r�4�Q|SD*g��
��3�M��q����ؤ�^"¹P5��L@#�q��y4xv� u]F.����d�.n^���b�1ԩ�{��UB;a��	�U�?���@�G��!�z.<b�~;�i�-�6�L���+���b�{��g:~�#!��	��
w5W+1=�Z�Fg���	!W�K؎�I�����~)�_�zB��t7�3����]�n��Y��>:�X06�/8�Wڇ����TV5���V���&�����Z��'����5�x�F>����K�K��UEt���m �`,r������lH���t٘���G����m��eAj�Q�>S�|�1t���j8���j����t�)qG�I�~ئ^F8���8���15q�(q[U��^|���OS|Ϗ?|�.��xhhP���F�Ψt �O��=�>	F	BD��)���T�Ksh�r�8qt��6���ȧ���6׍�;Rl���8Dҏ�r��` ��A��3�F��ad`H9ǇT��.jJ��>J㔢�t*q�V[�S���a
skH��?��:݄3!A��:��קa�1f�Ӏ���f�gCٜ�72�o�{�{C��n1�b��u��QH�H��b���KNw���x�=6�ջ��h��X�5��64���p8��P��b,%�ʵu˥	�|�yb_��7�QҔ�L��i/>F�"���K��D�2�p�/]U�/I5���U,��l�دړZD���ìt�E����Z�ٻ���#_Z�O����͈ʘ�`�Cm��E�7JD�q ����EG�iΛ-�2��� y�R��[q�Fc�@�uR=%����؜��������7ٻ%m�|���4��#Jp7/��}
(ț��/��P��zu�!����~�����ϱ8!�3���nd��ėc69�=���b�$ҪgU�W�k����!��yC,���)^�ϴ�'�Ց#*��戔��F�l�؆��!���ځ�3^�+�v��xm�˯,�mQ�Ku���xG#r��ԟmOJ�ǡ*iݤq)�E+:�hKn#Ү]W\o�g��dHQ�CD
����.x�0�fv�Z���y*\C#��4'��x���H����	��ރ��#��P�Z�lA����掛 nl4��ب��,�g!w.�=j��|r��כ#����9|t˹��\��+(
(��'s��}�deT<}8"4�%��'7[X5.��E�=f���ڷ]Dj������ x��
�����TzHМt���x��:��]�u�ޘ�-ʓ�t=[��1�Ϯ�1��DǦ*�0��s�QX�چZ�m��Tg7)�4�N�T�+1ψ�o�ݽ�XY�?
���9���p�zѻ\,&,��(��9;1��x���<��B���.��:�$,\$�2Y����hWV�� �1�{&<I�3"�R�A���bӓL��l���wq!��`q*"�HS%~��yI�n�������O�o4����%뒚��G��v��Oc�0���\0XU� ���x�Ւb����#N����@������EG��Tih6n$0U�5�k)����i��#���O[\�ް_��h<�
&�䭶R|	�Z�0�\o׌�L�_f��I#T�	�wӂ�T�"�x�u��m��T�:�v�1P�=a��Ep�Z����V2i�V	�{��q�ZcZ���!]�g�@1i[EY�H�"w}��7�5أb�G��iN�+������D��?y��kg�犏YN�i��T�� �;%�peRم0H�� �"�
���aR��[����c/؈��fK]:	���N���!��~��>����\a4H��M�>���ؔ��,o���w�q)�w0��f�ӆ���Ť�Q�%�b��dt�*n����ES�[� p�,����7�J�{�60,��3=&m.R/�d�Y��e�qY<�kz����F��sMo�0�j����~ۮ�#goVw��0S�}\G\P�8η��� ��"���8�T��w����v�^�������ޒƧ�na@���x�Y����{����=v�yFu�ӡỐ�9c�u���Ң0j��P_6Q�Q��]b~M���4�tC�� �}�1M<p=�=Vj�^��2�ل��4����ޘjG1�v��m�Sk���u�T2��\�������J?0����!�/�ע�T}V���3�~|\%�z5智+4���,T\X�������W�"����JjD>����|0��O�֜�b��ԕhHQ {�N����Jx������0�2���CL�m�4n��9�������$!e��Pm��5@��;�<Wj�S�Vt�6q��QRͲ�wgQ�]�lZ�5��� =+d��<���M���Gn Ec<����Z��#����Y�A�F�rM��Y��jG�k��G�jޫ�k��v��G/Lz��xn��\`�kQ 0C�%Sv���M�U�|����c�9�����F�tϖ^;�0��{Q�lHq�WuW��1��}��Ga�l�ը���B�B�x�b'�(�f�D�U���1��@���c��=����p����+q�9qP^�UtAgY���䗛!����d�^���tO'�;V ��� f�k-�i'`A�P�Z�Y�ON�׈"Ӷ�dc�L�%��=տ�3*�1λ��|�'��ִ̍���R}b�^�]���M-�(��$�m#^/�n���t�r��C`J0Z,L�W&\�)�%��JW�G�A���D���T�P=z�&��!�������W���@�h7��X�
���v/9��������p��|n\�P
#K\w>"R�7谰E3������=�7mBwO-�ȃ�t>���Fy�S!� Z{&C���L�|�齎��i䐨/����"$U�Y����3�����xT�a�?&�� ����-�����^S/��5�@
�5�j�0dt�h�gJ�W�_���j���.w��3K�*����K�+�{�F��8b�V�"7�圆�:
����G����	5Z|u�����g�ܢZ�'�O��]��"�ahF� [�=f搆����#�'Z�o�#-Md�*��G��p��Ӎ
R\?A��iD[9I�$�"��[����eڿ<1��x�c�9�֛��2�BG�nѢ2	��&s1�r�����̋{".�~ࠍ Z�B�̂G%�ՠ�\m5�!g�����g{����4PQ���^&�	��n��{3�k=(�J�ǄoĸDUu�L�R�����#����#a/B7{���^�*�V���-k7�� t)���j�R@��O(�˛�*uI(��hV-MՕQ����2^޹/�;~Wj:�G4l��nv.�������_o�c��X/)1�h�8��`�#��;���3�i+�T��bl��?)����㘱����J�&S��yK�]9v���*�&N*����e�N�A���z��K�}�~�ߜ� #���k�߉��h}��z���m�cP�=����uk�rܲ���>+�5�Q�N'M,�`c�A=�7�훫�̖�5�f�ĝ��V�b��r9Ĺ��FѷT%)��D��[⥶��cj_�8�hY�%�np%��{QO��EE�=����QXt��Ţ>��Ӑ�ct������Ά���T��T�$Rc�{.�B�FA��q��t��
�
q�ٶE<Z~KQ�hL��HF*䉞�k�L��J#�eH�����LV��f��CO�4C��Q��.����M���Q�#GS�
Et��"1�{r����Z��x�"H���,Cڕ���p]
+���Ǜ�����O�6{�4ε�d����N�[R�zeF��T����EE��O4��!�4�����6b!^J5�{5C��#�d��3�̼�������ib&��&�$���_8읱��kD��H����:�6֟&��ʐ�]���=����vkBa�׵Tc�jM˷1i�U�hU����|��b/��Ŏ�-��k��@e*[��u�C]�D�lU='���}Y|Ԗ�?�F�����ڜw�Q�?q��L�vU!�ѠN�4�%�~ȋ��/eh�������v�P�(%��Q�"���h,E�Z�����rtH;����Z|�=���t.>����S!A��.fD�+�*�ָt
�"ƬH�;�Cr*	w�}o���Y���n��
��b�����x��Um͓R�t%�
��%�Ʀ����A����� ��RQ�:[�q�%�r��"+s��q�7�.֪��Z+5B���s�G���Ql��i�^xN"�S~U!�����k�����K�4F4i�gj��;-R}�T�Ņ��։E ffu��;�R�C�_��MF�c5��+�3S�
 �b��� ��%=���\�VS�`�DC����Y�!��Pä!t�9Y��0pVW�����?iY)!�}�����.��J�U-fQ4��۔U�n��v������o��I�����1P��>YOcZ�b��i<��[K��`){�v��/F�g�M	�O^�SGeWi��tGQ�aH���Q몍��P�=��A�k�ۭ�����+e�.+|KIɱ�iQ>׊�0Re8&ٷ���̇�@L���Mek�Z�`�t��&��-�<G��zӺuiR`S�zu��;�J�5Rfij�wu-Ɍ�`����VQ�J�6�5F�����tV��I�Ѻ�Οm)C*i�Pt�����6�!�'�?;��y��ȹ�V�E�OO��<�`�b�"ϕ�ٹ��zLc�%��Nc�[���	~���(�RA�#P���р��0
��A�]��#�^%�la���_O� �o!l�; 6uc�Q���Ɛ�<9AƲ4s���6-��.�(�,�Z\S��RP�>)��
��w���b���?��il����Y��b��hѲ2�4�ջ�S�j��6��\�Pz�=~y	��E�L��=ON�G`��?�@`92�~�tK�����`�n�B�Y�M*=đ�]5�7��t��?�g�rArc�� j�ӚOv����4a(
@o<�3�MK�xȔφ�Y^���|!P��P���f��+���Y����*�⚖���\Y�ݶ��aX%*A<0"I:�5&W#�!�����Nfe윘����HqUl�� �PU����e�d:���#K���h�=��_�vP�ԟ"J<����4Gh��󪢌��E]����A���Ǡ�qr�C����*�qO =�C	����zd 1d�w�a���`M�ym��g��4�د�<�M�K5#�}�in�QI~�I����YMɑ~�|����u�"�	�2fc��*�Lxh�D��*���{�bl?|]=6:��q�}h�#��\�[ո�^7ʘXM�=�Q�huʩ�f�E*�P�KG�?*��ڊ�t�aa��!������Z@��ϐ�i?I��`��|�8�X��\��nP?S��ȸF���W �A��h�y]�9���;�9*�9��.����5���s��^ڝ���g�%��"+���D axb]�:�u%�9�ms�<Ε����KyAҪ\�m�1���)b�[�*\����H��Q��3���kZ�_�L@*���%���*ve]��n�(9y8{�������6�] �n婳�������LS��w��A>FpfH\�(�>���M�1��~�8t���]g�_Y�[��WR��s�#r傒��.t#F��7_l�zqi|O(�mN�bڿgt�jn�ⶸ���0�j~����aL��(`V䏾}e�1\kr��}�(�ef5F��>�K��c�\~j�M{ �XF�ɚT� w�:��U�э�8��~g��{�J��ߏ�8ztd�n�&0y���S؛�ӏ���аYXؠ�A��
P���5��W�gbj���^�*�ö0̡�
��pocCG�ŞC����G����q�/T��zV�b��"�&�T����횿��ƦȢGH~ 7c-n�Ԯ�;1� b��ո!�����P��0Nq���]4I�U����:!�.q�e ԂGd4�W�a��݌�]sJI�5F���&,m�[�����*�Ltw��^(��u����>6]>��O����jjp�J%/v�����*b��BG�fEة�����̏�BT�D��F�,��c��{�"��BX��Rt��1��'���}�'����g�)�jUJF��L��I��6�X���zl�;��?ӽ�� Χg��d&mй�3�-��R���`v��$Ak������,R�^'��撲a�ZI�J7�P,6��wT�
7(�71rz����ܲ��[Kt�`;6�suT��/[�AZKQ
���$��s�7L1X_��u�����C�%r���׬���V
��>�*��c�Ɗ���j@�۟xCq��r�W�kaHQ,�1�Tp�� /O�5�O��x؎���٧K��N2��؀7��]WG��(��Tx�~�r3Bcy���b�ޓ�uM1��:O(�S����9n�rn9�$v��`}��s@�"۝	��]���m���)Y���Q�u"��&(;=�ӯ��R�?���Ջ�>�G������>~��H���5y��ً���5��C�7�o���t���9�����U`��-�~�ɶ۹=�"��r�B]�9ڬxq̈́�u��K��*����9�b`y�8/�/���ð6ƍ���b@⺿/��1�wռu�X��N�u�������'XȄ�.��
�L�(�R+�U�����G�����1��C�Ȕ�N_ �l�H��V�d�s��ZF�#gjT���_1���X��\y�����`6�ǵ��&>��L���b�z�q���%�0��H�lI���3T��|��z�x/e�թAD�Q���K�F���C�[v|CbB�Ȝ8_ø������zT���J���젇�rU��I�"���Շ��,��y�yDF���x�BC:o�eݜ��?!�s�8����0�QRܭ�X3H�����8�I��ݜ�V��T(R��00>�Rۄ�4Y�&�օ�:%e��-����.�B�"�E���g��x�+�Ό�c
��"7�Q틞=c��7G>����ǆ�
cs/E�I�h=^��ub�Զ��DGˊz_U�6Í{���\?z�Ȋ���z�X��Ѩ��|�7���E�'�]F� ���E�0$��������ߌ�*"�W�p�<�:�ѫ.R��,÷��V�d�a���s9~�1�������A#�R��I���!�~��T�MWٛ��ɬv�����Q�n_�^�����+nk5�� ���X.� 3���n� ��Y�2��M�ƇjH��[�x���D�5��'U by�޾(���>z�;F���:�[�r�:"��xzu�ġ*��s��0�l
h0�a�x��ɐ�ۿ�!�.�)RJ�l�!�Ȳ��cbD�l�\�H��Érf�3��,7B q-Ðn絎���g��?+_|�y�h
j�j/���
�������B�Y�]F���34J�'�%ƪf��*U�K�ԭ�)�*�t���:����/�3S�eɓ���*á�uL'آG�͞�񬍓��E�0�[`=�f�a������Fd#���b:H�����A��=�7fƗ���X�ZL�q�H8�/���=7�|O��U814N��Q\�!0��Q�Z�,?��$n\��������,>�1�x�*U�IDj��$�YY�1f�7��k�ݶ��gV� �ŗ�>E����8�O>�����G�E��o��v3���z���j��X��Kc��U4�#r�W��Y;�ʇ�����䨑�TcagEI��Z����V�!7=�ڛ`O�ș��ۈ|����-����.+QY�xވ�^��{�Oh�fZ�M6�8NŤ��0�FąBJ�h�B֢J�{�=�@��@��Zn(O�Ņ4��4Lg�⭳GSD'����M���[���+)�S���#���Z�H�u��WQ�����R}ިU�k��9�wM���b���F�hT�%��{c���������]J�A��Y�1��H1
Og<Τ��b�����6���;hin�m8��#�����y:"m?�}b�*r`سǌԶYv����3p��g\�C�Fj�ZE����&3T"����L��CK�3�4���&�s|I�K{�W�m;�c=B�@�N�(�_Fu��*�kA�l8N�wNѝk�m�s��y�y��~sԐA	;�Z�k#GÛ�H�&����M���������W�����џ�w���wk)���[=�񖩥/�m��!�͈Uf4�����!"N�kR�'�o!���EvD����=͎J��X,��Rq<��j���$2�hIS��0V%��e�.$��Hr��G�ؔ��e͛��Ѱ1,W�*�*��v ZI��s�"�3B
�]y�s�d�9�9�8C	��B_�~U`�G�i�cl�(�D��G`Dq��Aϧ�xWGq���.�,�x�T��X��ɧ�s�8�qG�v�P{ū���ciLh�v]D�ky����f�^�1$q��7�4��;�}T��\#ϧ���1C�x�Z���oN��#Z �hQ�vj��R���!�T:'���W���6�\�H��j\Qz��5�+�R�jV�G0K��O��1��9)��|ּ*�m�yqm���s��l���d�=��b������k�sٰsME!������S2�v���i?���DFu-��7skL�)|kҎ���sW��4�	:�����s�S����;	+��	��:t�K92���Srn���z��nN��^΅�<f�ex�����l{�c�%�v	QL�z���aC�E�E���I����F��-�F��k��쮣)'��������{f^c<����xs�F�w����9f�GFpc_+���E�����(Nݟ8n9",��14��<u�]dl�UY����	!t��ɛ{���,��an`�>�fzmdd�u�J��}n����ê�h�8Ҙ�e9��a�$\v�X;5"�۔�R��
_C�!��0�#����߶�0+bZ3[1��c��tMD�\�S@^�Ͽ�"DU(}	�Q:w8�I�-�����Sߦt�� )��V�Pf�o�%�@%�nQ���Y,��,�T)9;0���1*0��=����E1�5�#)i�tp}�e�QJ:��ݹ%4����t?zAՊ�>2u�Z#�**�)�Ǎ��&�1��'�ψ��A����7^���0}:�811�4%%�ZZ�Zշ�(��K�@Q~:3x���l}T�`��]�e��I��o
%c�#�f����~v��F�Cu6���t���f�ɑ�R�z�A`�6���6-�C���<wG�����~c*����r�Sbp�<Iͽ�F}��j���b.� �A���FʅG@���̭�5$yȪ�}q�Jӭ��M�(V0C�ǖ�]y_8O�z�SgQ��<��iM���~
C���h�Pd��$t3翳��XqlY�N��o��H��f@Sە�&�$�'_�lL[��N���X��U~��b��ߥf���L03�={��J���z�3���,�ͩ	1g�jL�X�^���������oǊ�k���F�%K�l��uf�O��ZϽ�xj��|aR��n�޽�}����e��D�W��,�0!E�6��&���l��Y,��u����p�(��FR!RZ�MF�����!��19�v�'��宖��9h�"#V,��~��NA5j΢L��{�g�u��7C�,�Y̢d��L��9���i͋��Ϟ���)���{�5מ��u�@���-�Aao]k{cF�p����l��_h�Q�¹����y ��C��وn:�L�)72�mhmB�����"�#�PF��5.uMb�\�<!�q/?��siL\�aX�/�q�~�i���(���������$ֶj��2����H�RG�G����#�#�ߌ3^y]��u�P������y��ߨ���#�*F���Q�%u�s-�{�}�Ԭ�"zҔ6b�_t>6O��^��%�k�"�����e���"/���V�r��)Ys� v�~a�Z/���-�]��6�iD]�O���u3/�]t:��=��~�)���J4��.��b1)�`��>%զ����\,1�$:�п�{:�������q-e���Jy�E�ݤ˅��^��{�1�Y��"=HvܰBʛ�^J��מY��+\WU�!�|�ѳ�4��يF^�?�A�X�&$�[U�9?�Ƶ�,�l�V-���R/+�ہ�|+&��.������ǿX_��0�f�pNW:ɘw����������䀻��!��s�n7g?�Ϗ�D��O?��gB�g�kQ��*��.|��>q:eO���!fh!b=�Ё�x�6�*rͭ���5�4��ocr@F�����crfE*�D�6��d��9�2�*�y��MD����c*��.�$�#��]~S#Ns�B��\ǻ���R�*�6~�Aָ�OL�hG�~����F�n�&n8���m�# پ��]ҨN3'�F�R(x�=�ܐ�2�-��Ze�h�fXP#�'��jPCZ#Ҷ�^1=��݅JC����r��P��?چJ�3"�C��t]�X4m��-qQ�1�S'�h��[�4�qqM��s�Q���H�ZU�����e���f�\��-�1�FT��H��l��� �*��?�k�H�v�Uo�ⰻ497X�rϐ�1���e���w)�|I��5��#f	���<k�֢~��#!c[�ٌ�?������#x�����~�*��6�Yت�/��~��7��}�)��M/_���,��������!u	*���k��ǟ�w�}W�����Q�X�0z�#蠞�n���4҆��߶�����_�X��p�@���V�h�t�S�v�sD�f��Ԉ�U��yg�h*drˈ�w	��2�D%��& 2ѹ�k�\I�����CHT?��d-iHT��P`���)���/�e��N��Y��5"e p�ʔ��H�nn-���qF�Ci�O�xV�t�گ�OQۦֈ��W����}������E"�&0�#�R�f�2A�YR��I�Ե���!�G	l��ז�����,U������]��x6���^dbbMA~��co�����-N��e������<�!fZ�ac�Zz�ƫ�=�ړ���;e�x����^~�S��Tٰ���W��%@���	�"F>3btj�����" gʔ�S)�4�q�@Ȇq��_8]Rs���?g���Xޤ��8:��H[]��u��L���L���>R_�aP��q�����w׻r�g?��ry�BS�s�;��9�-d40>��%"ݟ�I�)�JX�X�Q�ߢB�*8(1�繖.W�g�q��������lǉ����I�p��̸�V�u��	p�?#��3�*�l\��9�V�;�����y��T1�4r����*�ߨ���:�aDb���~X�UU��ΐ֌����L[d�����J���e���T���	+1B?"Zl?k�I-�i�l-�AQ�(C3�Ȣj<p$��Lk׵n*�ox�7�HYawʍ!lå���Q�R���Ðj�X�H�7�M^��KP+��s��� �]S%��W"
?�b�'�22�!���X	�R�q%8����I�x�°t`�Zf��R��=�Ǯz��pԽ��,�° E���fHM�	��3���3\+`�A{ꚬ�:Ud
G��/?����O�.�ѝ�h���)`�p�f:6�{E�B�#�hup8D����b���l��L�
cX?�p�A=px�b]!���Sh ��1��_�`ǋpQ��/!��9��c����f�.ځ�����,91���Yu^�`�<���fAA˪���,;B%���?A��+�a%�u�U�9⡝���:vP'�L��Ei���u2�֙0��ua[tpp5[���J8�#��ΠVL�v&��&����D�{`����faV)�]���'1ӎ�)+n<;fYX(Jiz�V2Q�ww���%�<k���0�b��!�ڈ40���!�Ξ=St��~��W�\Шd��y2jTD�p`���R�xđ}�_�׈T��RQ�H{���Fb�ӆ��ōj��y�E��������ѯ1<o<�;ص-�O�<���m�.�K*7yl��$�cS�(���8��-���T0R�~��t�����(j�F��8�2���E3�Uq���}��q5��Xܺ���w��}Q����-��2R;��ݴ���K; ��/?Ә"��:x���kn4ڛaH1�.�^�FJ�0�5
����.i,]d,2�Kp���82�q�j�m�p���pU|�ڜ�U���1����JF�Z?����#8��A�:�T��R�LݳBX|���������o�}U�8��]��.?�+O&��R���K���_����OF��Z�6m��{ѯ�-�j�I`>��!��lW�:Ŕ���*=�O���9�&8��0�B�?��R+�A��"N+�������=��	r,�X��F�R4���J�nr�Z7���n#x�%��6!=e�0�㚴&W���Λ���!+�,M�5��IJ���{<ߧ%`[<).�ϛ1�1x�B���Q�ڼ����Vr����0���)>�BP`F����Fט�L6GKn�L�)�:\�v�i�Ny]�lH-��@i="�(�m�.�	��%��R[$��Au�*�h���Q����J9���6G��u~|G�6���O��l�
��`_��`��W���p�l!6.��9/�)���� 9��A�|iD_�Aǡja�X5�G�����J�5�f��o��ВU�k�ƀ@m�è�]j�1���\�2%G^���0�Uk�����:�f�{L�<1ޙ��ʍ5��|�裭�si���B��-�4��je��-�U��U���z���hχ�����\܋7\]�1�d[��7�*����N,%S|SX\�J�vf�׵')cDM�g�M�ֻ��A_hU_DsQt�墬Us�4��N�ƯN��vE}���N�۹j�wѽtU�8^Հ��_�1�|���~�Ba�1�~�(�U䧼'չ`S�h����9���J�O[Z��8��T�bʉ∧���ZII+%#�Z,�(�c�V 3��u����?㘀��s�Nu�"�I��VӒ����IBK�~��mctw�~o����GQ؁����SFMД�S
� ¾��H��)��8����"K�ɕ��x�?�~��e�)�/�c3�y���'9,Ns�t@�ևJٲ����m���H�$�w<F1k��zn��ґ���,�7�E�Mg�]�e�"jդ�M8�v��<�X�6w��=�F�{q�"�&�49��KNeVl�u�U)UX]ɷ���c�|�f���3une=�iȌ�/�wY;�y��\*N��9���E��B�J�ż�~�<R*pj���9Qqo���YԚ(���<�K ��j��n�Mq�0�仆^L���;��N�Y�+Z����5Ҳ����n�,����٭
[,��8/�qτ! ���E��`R�ƭ�ś�e_df`�4F~0.x�S��f���l�M1=s�Z�N�g8�F�̎�V\��oRg��Pr|�m���嫯��w�r��謺'QY�bK�2���#5v���ǟ�:"B;D;������+�l���o׸Ơ)Eg��Qb�2�^�W�܎�6<�5�o�H������{'>s�b�y�WICj9K��vP�5�?ѣT��ȬG�	�r	︍�t�^unžOYj�� κ�z6�,;�m��,��\�UEw��9�C��;x�?1����C#{p��W>b*��!�!ጦ�վg�k/w�[�Šy��R�ة�D��I�?�"R��x���K��S	�4�98�*���Įޕ�w�aH��T�F�5ʀ{�C�L���L���R͎�I�$4c�meշ�I7@��\J��PĪ�"RG"BD��2e�u=���s�I�H��.��5PG�\q�Q 
8�w~�Rߤ�o<���*���6"��\P�/[�X�
W������(y����YE,��co�kq3:5+��Z���F��5-hK�����P��G+�v,���~�Q�lL���j%�Ћ#RЩ~�"�I]җ/C���?��vD�Q&�|���h5���f��G�3�:��L���,�7����l�uAΙQ�&_8�j!x�>������2�ttPD���3����f��mW��D�9h�_��})����1�n�n6�������mՠ������V�������4ŷ�"~P�㍴+z4���E
��f��wHc��M�~@�4�ۅ�[,E������+�Y��b��[�1�6�JI���*��3�;���������T�D��>D���t!�)��@�S��#T�J�8�kj$�˸�fH��0PQL"��*g��K|W���c�h��-��0r�<�z�v���D��Q��S��Oʖ<�#<p�F�>3Ԕ©<0�S�P�KR{��Y�����f�5����%����(C�� ���\��j���{��Zώ�c���nxꨮ ���|�(�s8\��h�s�~)��[$
c
�j#���sf"2i�,��L*��Q����D
�zU�f1�t8�SJ��]�&Vg��jƌ���cJ(���Ԙ�O��e`q�L�"��`�:/�ǵ��4s�j��⼮Yl��Hv��4V�wz9sVm}/�fI[� wm��Z�j<�:���/��XR?��;.�=tv���;�R�As3Y]E��ZS+hlܭ�@�ń�I�D��#E����m�7
,��UD�ہ^7�c�,�w%SsM�r���%��ԧ��jU��C��4ҁNE��"����-�rH��7�9�"i,BN0��>S�"E���1]�=�ʏ�����I��C���w���6��H����T�z�����!�D��;ҟv��b�K����^<�7�����Kuv2Cٷ+cX����c��l����=����A��}�E���Q��/�^����������B�C*D�hU7�V0����A�
l���'F��b$ƒ�7yDf�x)��5��j\\��RKw�~-�������o���~�`cn>�m2��Q�M�[?me�����r.�=v���"�
��gh�Z���]n����Ұ8ڡe��3�[mh�l�	wM$�ϩ��G� �ZB��7F�uO˭q'S�<�����x^�����.L
鮕Lk���+� 3R|��p˛�g����h2���nz`p1WF_É�U�M��N��C���>f+��؍��M�<��@-`]�����6bGT�"	6��;��b�<��Q(�L�Xo~܊�_.�0�G�I��p�TuĵŦ��OU_O�ާ��sxn+��{ދ�^'�aH�����E�C�f� C)l��oK�6�R*v���&~ٌ���=Ry��CΟ"�|3f�)>��\�^�C�	F�J��V�R���>�~B+���__�����g��_~���l�i���kyP�N�����Z8�s��i�tq����Q��y�����'�.}�2~�1�H�7b�$"s��-;����$�J��~�z���]ُ~�9e#A��q>r��.�k�A^�X��{���<׌�]V��;#�G�y�b�>��{���q�/�;(gj`且�H��aulC�3�'�ߪ�Юf�c�Ac���GF�^�<�򇏮��!m�T̓F�߁�����ɔj�Y��8��V�(�Hznn�E�M��Ж�T�:~׭�����GsgЪ��M~S��g�u������R�"�]X�q�7t��u푯�|8�!!��ל�c��c�'�܁*���b���6)� �,�h#���M�o� ����"�E	�W8��������cEC���ﭰ�o�2WxL	haB�����p�u)�L~��8��@����a/�BY6vB�~��w�~[���W�O?)�~�Iy���a�ax�	��޽[�ea���|�}F���<Ρ�tٮ�� �}\��Q����~��1k�ш�e�k��g�30p�0�)3��bOrD\wz�yJSR�JWS[ޫ}T��u]��M��xL����gqe�9f����F���#�#EVM����(��+�j@0)2���$����2���Ň[#���Dv6��1B�("]��8�/� ��w�A��6Þ���49��|X�%�_��,5����3)˅4��M'�50��EV��"=�Y8�Cj�q��/_��"����Q�!�O=^��f��WE�D��b�g� z�w#�ñA.���X�$����@��i��(Ea��G��ǏH�x`�ww�D�m�RLU~RRlHG`�6<���͸|��7[���f�87<�l��S���rj��ӺVt�C�`H�7SfDh���KtH+z��5�:[��~�ڛ���)���+G憌(��et[W�����z]�w���w�bT�q�P��)�B�n�}'um��9*{&���v��~��wq�Xk��ʛ��d3���pA��������:�)�?k�Fu�ն�5��f��s�����<�$V��,Jj*�
Q�ҽV/�G��Y}6�[��1]<%1�N�!5vV]�!�P�C:�	�۱Z.)��7S,������2�E{��E���Zc�=<�5v�R���� m�q�b%���Э�w]Y�aµ|�0���/cs�Z�
�����n���XtMG_=_\� ���B@e���ZT��ٖjw�B�
����ia o"�������`�KV�=���P� ��[� �!��[c�*j����h���nf ZB�%|~��X�a�tn��g��uI����mH��v�h
��+�(��?ޫ�g�Xa���BV1���F������-��.!�c�m�AYC��*h%e�i�]��>�y�O��6�5���G�ڃ�^p;��G ��h�I�r*x��͈�M���$Ļ��)���{�D4��﴾���F�����~�Eekc����g5�QlSAqgH-�oԁ�ŸٴP�I�a��rf��_��h�05��
���N�u����.j"�)�4�v܃2*g�C_U�n�*p=}��W	�6��k�B�b^��J8��d�P�b��|�\q�t�]kEL[8@V�F�MTZ?w�dH��Qh���jL��K���Un��H]�"�A�1<2>�#. .N��
O\�EUwa$g��2-{T�'g;�E1���56<��04�C�.Q�6I�Q�%��$�E�璚���;E��=;�@��H��=�3E��j�D�|���)SO��;U��E�����Y���l�r���k5����j٬V�_C��믿N��)f�+"�!ϱ�������f�	�)
.��@b��!N�6���3�Ӄ��^Ʃ����q��6"5(�F}�NF��eu���T?�Yѯ�������)Y8�c\?�8kEP2Z�{���HD��}_�Y�yH��Aw�we�h��((�Q��'c���(��p�y�ax�n�����Ѱz��m
#�᎒����U�8**5��Ա�(���A��"��� ϐ��.p]���G�I��x.X��cX�d�0��^GWᯑ���S���30˥�u��J#�iH�$���hC;V#�bOO�S�`�c ��i4ԡx���Յ35)���,n!��W�����}8GUn��E`�
�\���J4�Z��=�|�ߣ�Y�������HU���Ű�Z�-��nu����HK�W�H�7=��a�(�E;�5�|�;F��V��Fv�?/1DMv��%(���?#�}��Щ|�I?� "�
#�s3�������(.�}�
��� pX�#,ցf|Ϥ.�Y�����ҍ��y����6�ǽB;�� �������I r�p����^m�����]F�2�V ��燓�!P�������oU\�(�ir������+�;�)�ݳg���)��fd:�Y���-�]i�&2�g���H�׼?�����'���ܰo��])�}����.�5�y��ٜܺn����v�������kd���;��h���}Z�b6�Z��0*mO���ȥ婢�7�"b�q=̅��I�޽��Z8��g9�x�p6Y��4 �?g�%�i���� GDq`t�s�Ũ�N$TĹ�������0=nț:~�'=�15x�����pA;Q�"�3N���K�<d�psUU􍶘��:���~�N���/���*��Y5�;�bRt�(>�$[䅈�_~+��y�m�g!:��?}Q>�����g��1���]֥D}Rj�i��`oOd8���T��������1�ch/�j���g�ך�~Uƭ�-��Xa�pJ�?�T�9��+D���r��I�0��0���sQ�p�/23���i\$�H�f�[^��	t�g���I�ݵ�Aj�����*���#G��NC��fԦO3C�� F��\(#�@�_����Ogk�2D=��	~��z�7(Ԩs�&ѳ�Z��FN�۱6�Êך/O�{��њj�5rP��]����хQ�.u�@[|�b}M�ۂU[ds�Ŧ����Laj#R����\��'�l�1Ń#%.ۉ�'='7q�۸كZ��%���
�I��c~�ma=f�y��hm߿1=\|`��B$�6�!)S�w�g�釒��{]�3�]�����S���ļ�ۂ�9r��@ŊyJ�uRw�H�U��2��ϊ�%�(�)`L�h���;��k�#�kQ�䩙�[��z��Aq��_�-� <E"�fSM\ģ��p.�-�f+�G$�_D1J{��{�yu�̄�J�8����1��ᜧ[�*X��WC
����}h�C	��}���O~��g�p��)�
0Fo?��PdY���}��8W\�y��^���W�b�A����Ґ&才��ms��������q���u,�-��:���F�BJm�.�?}Z�X
�,K�d�K,eB���>#�Z�b�GQM��i��କ5����P��ݎ%�Rg$'��}�z��U�S�̼w��a�#ڲv��0~a��m���}S�Z��Q���h-�����(�M�u�,
)��=ᵀCa޽���WQ)�ᩔ���mh~k�BZ�Eަ��*g8U9�:���ߞ� Y��o��z�����cl��*gB͹`�b �c�I�2�e���W]CCO����^lIu�����b	xaL�|�ȅ�tv3��������y'�8<�fvJ���a�@��~|>8�0.��>ތ�ˏ^��mE���3qa���,Z�h��[����	r�s�MF&�o焨�$<�x]�_���9����C��W��?DA���p�V���y���KS0�9��rt�}� �gk6�ZgcX�7~g��ؓ��k>�5��)�]�Y���8V	M~x8V=�
��Ұ��͛ ����mw��N��ɤ1)�:��*��0ɦZ�]ک�4'6��9�V9*/[~���������~�X	�>�NrIj�M$|��,�,�1jŐ���Y$lb�=�������:F!6�sQ�t�s�C�*Z� 
7dL+Lqu�:ra�(婎�����(���K��M��Ɉ`�s�.��-��B��IF��鄽�{�ݝ��k�%'g����(61JY����Nf��=��bn>'DIP��1�5*ˈp��ӗ��-�E
jL�aloM��[C
m�P�~�q-o��]Ch1Ez�h����E~����+��4��=�
op�f�P���{�p+rAvS7�\t/A&0n���8����7ߊ�L��~G�y��9��6�|]�؎����p0�_o�	�'84���(,m��NG��<;�j���nǪLt��
�YFq���4�=~j$٬@Z��Oc�7�ǞSe��F���Ŵ�[�Mf�XZ�v֠���<���u�T�5Z��
��p����4Y�Zo�u4�����<q�	�Q���oXF,rd�����Q��nY3nl���!���rj��۝Rt.�~�,�ʂ��V�S���q�47�-A���;ElY��lH1�BF�M)�,2p�MQ&�����_�UR�s2%ޤBQYӐ�cd�~?�B�>QfayQ�ע�nW1��tÈ.�:�+n�2�=�R(��16�5oy-)��+�eE݄�,	*w%ǳx\oܗy�E
�+�NH�q��n����2�6#�oa(����,b�M�Gډ����_��Fq�Π�[$����-`�����9@.�CP]�������F
�����\)����z%�0�?G���m�����o��pR{c�p�,؍ZC5j�I��v{�t`������8o�m��'����"A�)��J� �DjL��x���,kٍ�� �O-CQ�Swvڝ���A�;H�?� v>������
�����0���l|�گ�h{��#[�+V�r��mr��i1�>�5��4��]��1V%q�?2��E���h�Nw$U�NC�	��C�3��8zUF�4cφ���şm[��4KZ��ݲW����93�ѹ4e(�^4QӋ'���d��R䈮�0�3�i��#�,i5�N�Fb?�\E[�<�5�>wW�������$(�k洖�֚��Mx���QR��3u�fα!�s�63"B,�����sbఒ�|�RGp46^p5�Y�*��B
�]�Aw��Et��)����>	�g%/�%]U+*h8Z�w�p�p�	-��Àa�w�H���ϿG���P� �t����w-S�(�)p:�;i>W8ZEWpވ>��~����V�����$� �kP��.ڤ�a.�{�(�F�z�T�u������m��L��~�yD���֠�Y�׮����>8bme'Yp��DO�KN�u�ü�Q���)���l��{R:�1a&�/j;��3�d��vk��$�ڳE�����},jIe��r�����Ol�fs��*V���T��G�	Y���)k/s��#�t�+5��҈f/�M��]�9��"Z�=�O&��5����%c]:�%�e �Ɇ�!�:�a�z<4���E�?�MC:�M>hV���FZ~��bʅ��-��u�%k�e�"�6j�ƈ��Ն�3��W�:U�يo��`ҔX|� �uX����	NsUgg�A�cA��(�=��K�ԙ6��R�k��*T�_}DJ����M�޲��d
\�U��Gr��!:B�;�Y ���y�r��]���{��q���RC���F�H�9��oX@�Z��'|�駟�?��O����ߢ�t�Us:	bՇ4<���0��M��ѭ�k:*C����/��	��}ܯ����q&LP/�����:�<z�˺/X\[�
�O����B=����Zh���d�m�� m��)���UЌu�����p��9M%+܆�ܮ�����Ų�xM�Z_<�&ܼ��l�@��^Ly.�X�=��ir��u��|;� ۜ�zl���`�۸�c�����<��?�K���v�!m�����Βa'А|���W��x���&<܂����.������{����F����Z������Ѩ7�uM���^��~�U���80��B�w]m�6C�����ٳ�R���Jg��Q�gMk(H�̌Z�ʫ�#�͢�+v����w��	�����L���:b/��V��*���:��m��0�䍲�m��A�ĺ�9��Ȣ�҈��3i�D��A��zyK�!:�%�򀽻t��X�)�=��E���_����d�RBT�9��Y��J�����vD�塚c�7��;�5�
�<�� xZgw:��b�W>5��X���u�,^kc�[�=Ũ�f��t�*W%N�/0�9�Y9�B T�$���;��=�u������e���5%�B�`,yE����ȸl4�����:���!�tۂH.�m�^;�����z�If�m�NMqs�:��\U��}�#���R��s|q���������4ྯ��o�Eԡw���w�F�W��h!�A�ޒ'5v�4*�E�u���=��7�s������֙L��Q�NY��8�����C���{��n��D�FZ2v���X���NllG]X4G]2�"�[ve�!QSz��#�80���ֿ��aЂ<�Q���A��W��Ғj�.Ϥ��~"r�{�V֗"��s��|T$���+<8�jt�����)���J���F����8�G�̓]�k�(��>ݢ�?o�(i�}��^��wa����0~�M�]�� �c���"���!����t�m��Y?�:�8\�����~P�����k�߯���b�u�wY�΂ ~8<�#��Τ|o��x�B3�5a
���k�~����%s�f���6M�Wërxq�(޴3\c��j����a� �ܨ�w�/�)ǚ�cp�F�i�U_u��o\�;�t���t^�'F�N��c�L�KkPK�s[2BuJY�����額A.�\��y,@���>�{7��RqJ�\v'G����}��fE�璋��e\��w;.�"�o��I�#l��I�G�1�$���x��O~P�.�M$b��:M��Β���&\ґ9��+#��Ė�%�Q,���%�@�dBZ��Hk��?d���+UJ���/������Q�gn��3��J��iR���/u,�"�x���+��뺃(��6��®S]qn���ۺ�X&�)=��o��-��X5.k�R��$U�A4�;�k^R��m����hG�$�m&���δ�K\WXd����6^�Q�t�#�;Q{l$KW�_����ډF7��c�����/Ű���-�����JZ�
ծ�X���jT�0�g�]M��{�U�>��3��2Z�>,q����C�
�.��d�L��������z�����t�Ր�A$�q�`5��@�<�T?���h5!��!����2�6���J{yA/l� 8͸��\���Vꗁ��Kꔍ��+�FaQ��.�Q�uO3����x
L��Ȗ�\k��U �Ŧ6)��Qo��q{_햺��ޅ��۵�E��G9��~]�R9E?8�����1VZ���@_�D�+�_V�S���T_�y
��@�P���\+�+|\>���0\�Hm@�T��*B�u(��z4���a�W��*����,@K�ߨ�Nv�Q̈�>��s������崻IgV���Q��������va�q��bJà��hi�|��wuV"�_S�
߇H:&�n�8F���(�QU�2�9��fu��a�%��'r��u�m��|.��8L�pc���%N��;�"b�^������!�ac��3�!���g����!u����9rV�3{#��yN��=$;�T.�	�������Ycs���i�;�4�M��vȸ@`���.5��xK�;	h��nS�|�ۅ���Q���%

�4�У?���Qh�5�!�hy���]��H��E1���R�7	O+��)$��<:�����ңN�t���!��`���"B�N�:mOA��0>.�#�ш�ψ������.���?S	݆O��g�}��@�1�:���"��)�!sc�3`\���?�?m�.�� �s�.)MŤ�2h4���ӭ27�V�Ҭs�ݶL��Zz��v%��sD�������
B0�X?�/�T��X;�/0eD����K!%�EL���g�!F:>���17�4	�X�4�m�FF�
�0ϐO;[K��g%����7;砗0~L�����@��3�\��Qo�ڣ>Z���F�������p8�u.ָ>}��X���լ��!��p}�ɾ��CR3tP\�1+9��މ��ة'&���I�k��F��9S�]��U�j z��T��E�9�֌���e4ZJ�6��!����S��r־� ]q)]S�Q�)�_��C`���hVM7��Kc�ܜ�ٺ0�o���~z�������X6���n���n�G%�l(�s�9����)o�jS�C�,�6
aH�������^����w��/�����c��1x�Q~wL�i2���hFx��an/�v0 ��ҿ��/Q�7��s6�7��נ�E���X����mV�,��J9��c�����E�1tn3DW5e���>x�72��H�h��t��i
��gwv���tO}�03=���)~���èk��<Bpb�p��,D���ʑ��Y?"ړWj8���.����E�tI��4��$�<��ru6��P��p����z�b��,b��o�uDCzK�8 ���D�0�_|�����V��gʐ��Y)�1�5l�#8ړ��(K͝��}���Zkt]+�Q3xm������F�������m��ɢ�	�K�T��M�s*�,�R�I�"+U��SϿ.�+��T��:�t
h垵iGe�ʒ��nw�����j�2���]6(�$��k�s�[�5��cG4�݃�t��nt��G��*�3��l��4
ÕS��V�5�s�l�Jc�}t����`��gI���R��5k��tJ���GN�|��]��Gt/�.�s\���8�b��3#�y��mW$�Nɏ�`]w����I�hs�~V�I�>�I��v٭�l��9���]��،(�\K�:���H{U���G߭�r��Q��F�*�I��R�ȹ���q���2�*���Q�t�k~�<F���%�D�;LB$׆v�OoѦlu�U��M�R?L��P��{\��`�����|/�����x�Á��̵�`������ZS�r�ܖ�N���5����K�����\ܡf65��ĪQ�*s�Ͷ�A����=U�{W�z���2�/�]D#v�H`��;t*���86����(�4"�4���ÐD|O���n�]j�L�5�����97?6��U3Ut��)kױ�Pp��ʵ��hI�x��	g���X%�.�N,�����Cj��0��������y��_��fI g�e�TD����e�M�$���9��>Ȉ:�+k��(��MU��Xx�͘[�(Q������?��d&���01��\����ET��k��񘥦��ӳ���h	�H���B;mН����ls��%��^�����k�[:&;W�!�;������b0ju��Xv�'�H��B�!�/�9�4Z�Y�C��]�c�&I\����>�!rV7*�<XTAJ[�E�(P�	L�A��z\<V��^�r��%�B���"�J����F������}$�z�/����x}�ٔ��<�'f�W��N,Θw<q~6�}l^c}�����.�� �jA�'}D�x��VcY|���
�n���ے�tA���0�N�p<���5h�R�xh�ȡ�Lה�s
R�~��0=X�Y�e��v5�_Oݞ�#"SA�1�3?�zJ��#�"�5hvT���T�
�VP|��˟���)�G����?]I���ގ�=9����7#��' ;ߦYƠTgx��(�{�9��
̈��z66�L�ɱ���!ź�J=)�Eݹ��T���,�hk
�;.ˠ숑:>�tj����3��h�����be�WN��H�5��U�9Z�I$�W�M��-D��s}��t5+@&@�F���p۱��}���퉨�ڶ�c����͕\ٵ�$��J����`Q��)��j�'�������y/Z�*#�NbG<W��q��	��l���:���}�e~bH�DX<u��d�[T�>܊Hk�i���̋i���Z���U���	-*��p�"u�y�i{[��'OAcPuӂN��k�J昆����;FFE.刦��07��T�,����{1o�otzϓYw��J<����J�T��˟7X-iAk*����B��,yE���O5��0~'�,J�FcĒW���L.��Q ��B|J��lpd�`)Rj��55�Y��yi*"6d�n(g!�q誂�e�~��(䬔�����rS��k���/��(4���x�~��>5��ˣ�vh)�H�J���Zi)�_��q�Rg;-�0N���A����Zm��1)���k%��q=K�� :O��Yb�oGqa���cmj����y?�7� x�h^��V���t���|&������~�I�v 1]�8�^�*/�]�o�J#M�c�w�������iIE(z��6Ga�S���J��b�(PSMk�|/�Ջ�d,������ǻ.M�3H��s��o}K�H�����~7Ym�ۅ�5m��Q��꠮{E^-�LX��I5t�O}Wv*�2���+�ۧ�C�F��1$�ȁ�pd&�tgʈ�c�1-��NQ����/C�������[�9h(J���/��R�ԩ-���ߡ ��H�_b2'����g����[���uI��}��t
���B�8�����R���v~�y*�c-�hBa3NbuT+�@�NLqCs�l�W�GN%^m��F�W�i�}j��u���i�G7WZ\��Qc��(j}�>>�(�ПP�F�R������U�@���T��p5&\�{.p��~��7G�<֡�x.W�$"�Y�:�1v[����^Ȅ�O-��\[c� �]��s��DDG��U����wh��I�3�Wu�2ݗ`<r1?��;{o3��)�{l�#���w_c=1�J���� ���Na���R��E���蜹v�=&Q�0�Uu��i�q�v8��N�ya�m�g��a��	���d���ت�o:�n���)�?��,�ZT�	w[%ѽԈ
\�"Bx�HQ�q9�8q��a�葑��=�ד�h|����e3WnC#ԝ���Wl�ܾ��K�{B���U��;ӈ_/��hBw���!��ڦ�}x�M�Z���?ǽ�����r�!��*m��yW��k-4F�*�t=#�ܫ]�g��F���/����o�OY`r���͚ɸg�pL0�6�������W�\�`H�V�8�5�M��c纇:���A���Ru�K�'�n�s�{~<O	�$�#����b�0�j<:ʖ[fgf~�8o�e�ƃ�:�ҨK����d�,��eۦۯwV�T����ڐV��ũiQ?��R]<B<fy��������!m�`��_���I����d���$C�����x���HQl�c�8�C�Ԉ��R�|ʈ�T"�.��o���,�h|00�Rv'eٽ{�E�p��4 bV�Ų��A��[��7�V�a%�=���>�C��$�"Z]aV���X>�;�,��97,���r��F|7�5���1��t(��r՛��/2���_�ߏ��ׯ?ۢQV�?�{��-�P���������:��[\꣨��/�3;{Ta�J_E0����Xv/��t�<2{�(V0Cv�dD*#6P� kz������#M^oM
��F�G���x���T�b�S��>!'!����ӑ���Fx�;v�5C�]Ȋ�k(����*ϔ�������%�r�(�6h��*�`g�����2�+��{����ω�{���E<�x]o��_a_��O�y�>��l���^؄�z��R5�35_��PZ	ZM9ǵ���X!�]j.��	|�.��.��P����_D�t�b4��Ԑ�A��!n�u)�Z�A��WsJ�
'2��E.���"��fQՑ�1��9ӳ�b�����y{]Ǌ�e�ےF�8Y{1S��@ ܑN��w]v�DBE!V�ORf*�K�϶��(���H���{n&8%��0ڦ�v��a@`</Ѳ9��"F������4-<}j��p�2��C���[u�C����a�=�x�j�:x�0h:���a���/�����Y���5H�PA5
D九CU�Z�Da	�Q���,)���\��Uųz��N��8vDs8�A?c�H>6v�3W29�i�U���f�L("��"��oa�~F�>�Q��ШRtܭ�S�rJ�!�J:��d���,�u��X�IYՐ�xy!C-�]*��X/�0�p���LH�65�֘�C��M�[2^�	�c��q�ޚ4�m��#��T�="B��O�̟�V�>qU�;��n�,45Xl�*�"]à�����v�Q�\����ESDI�i9M��u Į�j^����?$�}�F��	x9��\TI=t������h��-�<Cp��NB��9�d�ZS�X�w��1d��k�91Ǽ��W���d8��D`lB��x,?x3J:$�5Ƽ��.��t�������bRxg,��#�h�(
E�����QFJ*1�|�V<��9�6��˚�����I[���,)"��c�mH-���榉�}O�:#O��Y���3'<p���ypG�����E��D[lz�qF�iD�px8��3�<�a���9��\�EE��)�O.�\�q��UǱ1	s�1�H������OֆM�J��8����G�A3�I57��&��z4f6��T�6HW�A$��L8{�W��g_����Q��	�RL��~l���ר��JV�N8���ħl*������*,
T���T�rڽL�k��!E�-����!�U<I+��3U�c�=��⁛���"��iG��`�ys7�+pו�ô�Ò����@=�(�b���2�K����T����&Fz,��"b���{��Ҧ��XFW�|�ICz͡y����zS���k[Ȝtz ��D J�z��<RD�5�3�s�t^a�bX�VC���v]����#�<q�0��P�b�[��Ɛ5K�ف�g&��s��'eNYxd���\Ӗ�����������q��-������ÐZ��$��7"Rd;6�7�Z�kK�DT��=�/\�Y�r�юV�f�WE��]�Zz��e�<4$�?F4���4[��ɐ���+�x�~���\c���͠���Q�|\�s�-��pB�CR�'�r���4�Jb�}�tp�@CBQ�Ђ��q<ƽ��5���^��׼v�,m�<"�JSG��Cl8����Gۛ��q$IW �%�<=���?l�ݙn�$�@U�infQ$u�ՃEudFx�����{i��$���sׯ�@�.��COX�Ar��$���_��
��_e�]��ᒅ�n���Yz<4�7qQ���)+	9+�Y/K�TK������7���w7�\��fٞ����Ξ�Ln�1i���b��U��n7ǖu�"�)>#wA&;���-�,_I�6��ⶄU���*f�5A����D�L��=˙��$�����=Đ/�|����4T���ĜA;X�#~~��`�U��盤���c6{ч�TkrKOSU�7_�YpFಡ�?ݱ#�꺇�{fa,%#C���'TP������St���F�B݆ڟ��c�^����U�z�;`�y�*�>�;jOV)���<}!t_[I7��m�:S��r)ל�1Eύ;�ќ4�_���=E�G�O�nz��!���)�{j=�$M�=׫3��z���>��Z�~W�Q��� �ܾ�:7��hwz��^b�ۍ�7�����_�w�k_�t05�:�MF7PO�f��LE"�
�5Q�8V���e�����+��H�E���� [A��<����t�m������Ae?�h@U@�?S�98����N���7�|ZA��K�����cF��Z��p9�[�v���ߐ^�
�t"��zY�Jڧ�$�5�2��1��z��?���R�Q��R�.6̓#��^�
���]�+�/m���;���i�{�Ԗ�kv���k�i-����R�(��Z��,L5��"ؿD�j>/��sՑ�tU�>�A\r����:U(��Kzv٨ժDE�1���}���Z�7���I�K�Nl�jc��^����E9v�]~2ஂ�d_o���W�����ӧAw�(J�8�p��!�Xw'�N:�P��}�n�\Is�Ţ2{:�brp�CԦ�)�Mܳ�Z�c;n���$ǁ/� vƜ�p�I1�VtH���5�&w�	��7����kM�w�I�m�Ѓ���'Q�Vaa�Y������8�YN!��1nJ4�����!J��*�j��+SMR��3A�:�9pyy����K\h˩#��a�ün��G�V�]g�����rw��*��i-R-�n�7�=�X�*�I��i~�7	��Ԟ�#���$M��l����r�F&���.���G l��9��;y��0��2��2j�<�!��%D?���YS]�mv/�=1]�Q�F���h�!8B���鲳`W(�4�B�������S`��^6/d����ŚƵ�e�>O���M*��%�Z�pbhM^��+����sM'98|Y�ĺ�hs4��'��&�=LQ9��^������E�������*ؤ� �� �� �ɥ�z�����1�W��� �v�#f���@���ҐO���^Ģ��V'O+�V��t�m�=���,�tCg��m��!�'�]����h�}���o�Fr��}r��s�|\���L�n8͓�#dCX�������������o�dF����x�;ix`�I���ʎ�������ÿ��K\���F�����-�S��SE:�<{u��B�K�Y��u������I����f-��yR}6v�OќB)�(�uI6�f ?�L�jy�k@�O�!�k�n��-�t�*@{���
��l��a(^=�{h�(G��3#��G��C��3!Cw!�&q@=9-4d�G��$�`H�;���gZ�|f���b�[���f'v����"e*MJ�^//�)@mKd���'�d�]Ng�`f���P{8�rP�
�2�Yn���� ��|B�QS]�T{m'DD�����堄�d��Z��.K�k��	d��fCC������������a�����7��;��%�
�t@E�set� Ȫ��s��|b��'Ɗ�$��������2u��'
�7�)gk�l?&��,r߾��J��&���2��Ϳ�����+����[���-cq	vp�Ml<i��>�R�"�u���wఠ��������3�ƠjQɃ��2��֘ePbp�bb�������g�Pcv}\�f\��F�W݅v�N3PK��S9�j����@Yj��X�Y��7KG�&s� ����#�"me��`bv�57�-�Ɲ�#���yF/�ezA��B��ћ�d78���V9҃^�Ճ�r4���rZ�3C9iZ-Wc��16*J?�ǍƤ�*8õ���(��N�"(���:=��I8 ���/���N.����@�sS�[�o�'b��Ab,�x�ֿ�&#��2�}�z�������C.�6��O|~�����I��#�V�t�}{NћC�z�������Z���0�):��Ԥ���]��\��舲�!�����p�Pu5)����XݽrV�}�:�h�*fCZA�4m.M$[��.�j�xʟ��3Jv_`��κ��<����[��.�BC<&Q��=���:�!�;Jz�zn�0���6:�o��y�vdM�xP&�I�\B�$��؄Ѕl8h����ufP9$��R�9�i��;i�����C|G�(3Y�m-�6��GM� ���L4Up��uks��YF�"�����$J#�~�̏�)�Y(� �\¿I5�)6�Sl�
C�Y@\�p�<������Qaʟ᪬sTv�����A)��Z��)���,8������h�5���BU��7>�ǒX3�*h1�P�8m�u�jz�v�fp�(	F�����O��},���5��{~��h���D'S���uh�P�S��r5�g�E#�d ��{�w�_��!SĎ
��"��	�������
�]��k�X�ȫxn)u:��N����i+JN����sw 'm��Ϧ��]��k��N\\)׆�iV���7+Q�ǣ�ߐ����W��:��Az�vus�k��"�?<�wCI�쩠�r�F�R1G=SL@�;�I��\HY>���-�6�GTL��ׅ	j��\h�D&��T��猍���X/>w%�.�$�H8�ZE�y��K�@�����{��8�{�Μ�>�x�d�^��~�46&Kύf譵YR%����?�Z�&�#���c���E����C�øn޿o��G� ����0I��$([%�8���P�����p>~��(�0����%�7?EC�Sy��w"������_����*�5����~����im�J ߼?>��qGU$���<�Lz�C<�C�0W%#0�	Av�	�Q�9�m{�r��;x_����ϟc�j�	A�f���G9�:I|�����X�
$R�j�1�n���>�}�uP�8т�ҟ>=��xo8�pXұ��`Ҡ�5�0^/�Go���F�^瘘�0a�=�}��碵�S�0��[l4��ju>Mk���l;#�$�MY��ɫ�^�x�ke����w)/��
�8^eñ�z�H:�c�W������Q�i/*M:��@ܳ(-k���I�\b2���K�[��qҌ�׈���Kx�<�^U�����Wf�F�DE��k-���v�1�`M�'c����5؊�u�ȼ �ahW�K�3E͓P����\��#�k=�ѯ��Җ�N99Уt�Jt�\].N�a/��1샑M!���	����Qvɸ.�PT] @�u��X#�{�z*�Ѐ���h����Fc�Âd�x��P�w]8�rg�?b�J�O�M�u���:�����?
Yt����90�y���}P��}��9�i"�5�W�
rm1 �,��@��w����M"�>Ή�r"���������Qd��y��O������9އ\"�o���I��?�(2a������KH?š��A���f�M�����}ܶ1���A��䃄Vnӵ���W��*�i���0���
H�T�����G�`W��+K��k-�/'*�ʦ�#ַ,�R��6f��|������m̮��4x��ã���@�A��b���o�5�}��B����EA���ZCЃ��,���7�v���"B6��g��V��ܗ�0�lQ:z��"�<�΁x�S��t".�.8���� ��6r�,�l�]��s�QS"H�r�� 1�¹�{~�A�v{��e�nI��\@�����MA�Q�]#��ks YB)Q^�xsd�����9>J���q��(��u���T.�1��^�����R����#�b����M��Ƿ���G'��Z(���&���G�VO�J�2h8����>���,?��kc@���[�W�e�	Ki7/���P^V���>V<��L�C�e�0����X~��;�ϟ^i�c����8��m���Ĳs��Ʊ��:����.�~�6�H�>{v�cp"���<$������q\���qd�x\d�q�1�z.ဨ�x���ஜ/MϢ�_G��&Lr�dlg)v����z����3�k���҆��)q�_�?�l���DT���7�+u��&5��.
��6*g�ݾ�#�f����<�Ήz��d�5�i%w�����N��Pl�Aafr����t��M�$(^G��}��F9-��R��jx͛�uIk)
���6i{��)+
�"p�s(���s"��i4�LD�z�Öt"���¨�T��ކ|�U�O1�ݕ8<^� q[.�T�G ��U��׽U��Ɔ��4�X����N�)�2Q�������t���,�oH_?F0����3�&���h3|�h������E�1�V�����Lm���A�]���^"�}]��E �H�P"C �k�Z>��%��g��X�� ��� ZĽ��w�����a����JTS�I�Gq/������1_��ܷ�AΚj�3i�3�8�=JR;��J8M�b�E�Z�k0O��8��tן��9�n�u61�zyu�\��s+��f�����q8a�]�& ��/���@�ʱ�7�dwL�hY;���9W u�� s�I�^��gB*�@ϻ�~e��6YR��J��[42��;N���m8����Y�^4	7�\���frt��D]e�]d]���;/2��"�F1%t�EH�Љ�M��s��{��뚳���`(�_�I�A�ڳK@����|�G�6�ͳ�ЀO���͗�ٳ��N+��*>��W���5����c�|w|�3�!��CK����-$�@�ڢL��A�!X��#3zz<EF4��g���4�YjH�P�6�f�(9�m�p0$pH]`>}
�A����gpoH�zzzZ���Ncઠ�m�ff��4�T��'�7����/�	�ϟ�˻�~����4�2���5������xo;`�ȑ�a��������~(03BFZ�C�����=�@LӞ�ȅ/ܛ�;�Jg]oǚ����t���XC�g���M/Yu(s�D��FjV��X�rTz���l��N�])��X� ��}ߘ�ڀT�'.u_b�����Y�E�1�!�g���Ω����zY���4�N��N�ά׍w��j!fKm�֌��%v������5�Ly����{!2@a�������<����F�]�8���C���qȔH2*���D�.#���.��i���ZF�.�
ϰb�F�L��=�i���D�P���'u�%���E��ڙ3�cgg.bdQ��cr�(,��-���+�	�^��W�ϛT��Ӎ�#�\\�l��fA�9{�Y-�����A�E�?�|Ytd�ȓ� �m��lݪ�!�R��'e��I�O�t�y����Yu�	���&XP{?2Øk7���z�oR'�2c�'���*����h�@D΢vE`����/X�`8s�Pƶ]���s=�������sw�<��9b����[��቗P*�4Fv�l���1֋3y�q�I�
�1&����Ou��� Iȝ�߱6@g{~f�fyʃ���M�̓�b����AL��Ǟ��^z��E�-���vS���+v 㾭�ڴٴ.k�4u�`k��d��Kh7��EV���qm�(�lu�� �L���|��!�N�V�Q�� ��[�@b(�֨֊����7����dvϠe�p�<�;�&�O3������N: N}ʾ�l �K	�r��N8 M�2�cw�����SC�h�$�CM���S��u�v��[���6������{��[�6���f*11�o]�[���
��ѭ�MG��YJ���Q�l�����q�:`��B��48�륈�9�%�?��Oy�c<1�"eL9�t<��f�82�z�`�yB���)�Z�g��Ee����^�
	!-L�I��l����ŭ�E��D�9�f�]�)����׌���L	x9\X�w�38:f���ؤ��I�}/%OYŁrҰAY��O�
��a '
�#x��VѴ��D��!5�?�R�nFl���f��(�W�V]�m3���M!��F��Y}����y�������Z�>�߇��'/ٱ$�TдH�J&9�V�|���G�{���?�[����ԋvc�h[�Y�	ߜ�s΋�bw��47(�����B�˼
nZ��!#m�Ѹ�lt;�c�.Q��L �:�(qv�C�9,��:��Z�0���,��!PY�|���>��q�'g��5�K^h/�b&�e�p�#hE��j £�\�ө��i�.阞Y�2R`y��u�(wH�-
�2R�U-�=~��1I:�T�I4�S<�cp\��x!���ۏ�!�@���~����u\W��m�m�ue���@J��W��{�P1ե	�5���ag���Y�f����˨ό���C���,�d�葝O·�~{e�$�[�7o�i����\]��P���އ%�����mHL;�A�+!���z�`�)��ک罸�@sוR���kC�o�F#;bʟw��U��E�Ӏ5@�^�p}N�Ep(���$V��vB��cÖ�C�����?��A�>��Q�GG���s�w�E�RS�=Pݧ(p~��U�Ө~%-*�g	~t2��������HsZ�� ���)�2+,�1�G���EK�?'U�����]JB&ʏ'l©�"��z��/�v#+�N�(^�R��S;��5H�A.��x����&jZ[r5�f��,Ѕ.��+I��,b� �Mg����B�Sf�=�j�<@Mu�F��4��C
���M4��ؕ�F�3��妃U��ڠ.�m���XJ����pd�H��e�u��H4������5�;XV>3�Q��E�A����kN�W+p�Lԝjg�س��}5c�k�m톅�����@�e�Y�$�֫��^���#56��N�%R��o�@�����;��ٱ���-�b����<j?@����y튣-p�|؅�^�5�SOy"�k���~�K���Z1��l6�@���b\�ӆʠ���7(�gG���g#�i��oc��u�"Et�y $�T6���YV6�"��}��i�D`e�{ٚM*Ŧ��d{S*E�� ն�iVԬbu`��C2e�)�/�S<;��^�Ag�r]���P����@�g ��"��ɩ���Q<�v��)+�D�-��PI�C'�G	��Y{��G���:�2��|zJ򼗨qPܓ���u -f`qz���fxC��K]�J��U���d���ꉁ���Gُ��<���%�r������򗫺��T���$y�t��j��dO�)��vZ���!qH��Uƹ�W�e�IRZ�0��<�	�a�����W�w@Q�۞�d�h��Zn������(�V>q`k�ٍg��9�}���At�x����*���/��Y4������u����Z
��x�rs�Y���͘J:}�VGPA�~�<1��βXG���yNT�@����+��=y�\7�n�
:[��Ak�3��Rf�x(p�eS����Le�S��4t�%q�:�ϸ4�閥�3� ����)�*ŵ��̦��3S���Ag�L�&�����sy>�'8��z�E�b�e��H/1�s8&��2�&g�P��|�@�=?Jo��1��A��x/�J��ׯ�����D�}��9p��Z���)s6�\Γ�>�ߡ�8��r��2����`�x����p=qDl�ęnM&��D�EA���_����ս�oyy�,����Pl�TI�#�)�u�v<��QA<̗gk�.�[���&��L��6�$~�A-�N�E}�T���*�܅M����IX�*F�C��-� ��b��� ���Ӎ��Kǆs&'}�rG�|?��O1���-(��L�?����0���:Q2����tk����w:�}/ޤR(T�vnD�xx�}�H��ٳܳz_{��vF:@����c�M��]���(�}8@:����ܺYT���M��K��"��Yw�/w�tSFjm�^��m��@fO�������x�d!����M0�)2��כ&ep�%/����c��ڙ�Rc�1Y����2�~�����E��w��V�"40�?����X/(��;�ie�a���n|t]fQ�?��~��j������g��T�JT1v�{��拌��Z^8ʫ,ބ�<Ħ1��K����E ��XN�H��Ǣ&!}w�����)����?�/:D.z���� ���ݓub�q��JQw���:X�ڥ�gJ�i��j��JJ1{&�:�O���A��R{��Ą@��k�5�?���m�-��F��"��z�MNc��_Gį��� ��Գ�1gt֔��iW;�E4�Q�ZX�I�-��&뛆�S ڠ(� ��) �E��>7���k�qRZKf���dBD��v�TWf �tƯ���?���1OS�Lv$i|>Kpa������:�gv�դ�@��_��)��U�#����#F�48�\�]��?��l~��H"�^)׆�2���U��1ˍ�zzb@l癱�0�
n���~F����X!��w>H�ً={���{#��b��.&+��h>a�}�v)�SWXx,�.B�A���+���w�0H& 6�����:��P¿}���{+�����uVy���[����8i�b?ZfQA.��:�/�=�/��N9�΁���l:d-�iv����kH|�b�����=�P�g���c���@8�4�[c��]/�t�T��{�԰�ޜod	���"��Tc��=a�[�w�L��ke���� `�58��E�G�����{��ߍ��;$���{7�콦ٝ>�f���&�7�l<�	��}���Cn���\�q�^��o�(`��]���F@�SY� �˸�����b�:0����x�v-��73
�9�<ˣ��%>��A�`AK{e˶���l��%�X�F#p]լ��9�1�[��Y��*�8�j|�Q�hp ��cZX�1,>h�A�f(uC���%Ki�.�+�������� M ��qm0s��?�ԟI4;�^���_�J���b�G�X��9�����}C���������=�c��|&���q�,����I~���di�2kF>iGRײ�B45	~_�`�`��cTdNڢ�dt��f�³|��D�(��/̽n�K�\]
����M�[7Gs���t�t��Vj�/u:r�(��Ȱ���H�{��4�>�f���b��V���%����X�+Q-��I8i�i
��B�����%����X��K�m�>�d3��)�S֪m	6LMׯ�2#�� �U��e��JXx��G��x���
)�|J�Z,wO�M�9��M��6f�4U&��i�A�<vC�Wף��YQ�����Bdիl�䅮�;Q�wkx�[�x�tVĶ�4(��iu�  !��o�������'�4��tV�Gf1X���p�7<��+�;����1��?���as���߄;���V������Z�1=q>~Y��jV���	��93(�}�>Є�
V�8$ı��� (�i�w��k���ӎ�{��)���y��90@`[�ەk��������fN�5)����*�#^/��cr�)����SB6uϲ�������p��"�[��UMKq2��0�4�Q�H�Cp����T�2�#<ΐ�T��CvQ��MUK7��y�X���d�o����/]���>�BAu�%��%�48���ڹ�KzH�/��[�����;��=�[S��}(� e�4��O�ւ	�����5��:�U�)i5�TU�M�pY�7���t�[<����H��S;�M�����}�p�j]���'v1Mb�S���i7�Ry�6��P9�p��"�{��l�
����Q�`�*}~~as�~[�w�8�!nR��s�ĩb�\�ul6H{��_�o�mN�0!:;��q����.D�q���Ø~`���ld��\e4dN��ŦH@C����3�|�D�0�>���Mc�^31n(̝�2���U��V��1(�|z�u"����o7lOE�|oN*M�Zi�b8fO�t�,3�:�V�#yP� ���b�w{���oѕjC�ƌ/g�I�� ^�2�4=�4��	��mKHq���
������^̓�w�y�i��T�Z�����S������_��^�m�:��u��	�ߒ�]37(ğ3�jbx0:�~=!���)J�SLEt9�L�^�i7���o���B���<�a�{�h$��Jadv������ )�>Ȑm9ι���5�N,-��Pv{͸	��	�W�=b荻����x�uEP��`�������X��Մ�?<=
Ҙ3�<�#�,n/����8=��o� �v�q���9�u���hx �GV��v6���J@J6K��-%�kB��9P����i��;��A�J& z_+�u�"�?�߹�<^k���y&�T�7�d�+�v��T�Ǝ��k{��!x3��^�Ǯ8�����s�M~��b
�>�0�K^<�Aέ�g�=o)GB��Ps�|S%E�ʸ��3f��M�/ga�� �aί�F
��8��ޜ�G�i��?�9�{.�X�t�����F�"�ޕ���&�6�Ѷ�7��[�֓����ds�䲰9T2���^¢d�M�2d�����o�����>	�\7I�ֳ�u
9��\Oݦ�o7)3
`'��}vm�Ɨ��V�H�ͅ����nI��x��3�c���k��4'�z6�u ݄)35���ծ�%u)Wa�fT���!���~�v~<�n�U���9����\�߾��Wo*��ש�IXup��L�)����qN�<C9��8W��X��w���9�g�������pQ��nuܷ�@�D���R�z)[M�E8��)�~� ��[��?����� �
�l�1�@�j�M�A��]���̫�#p�~xT�q���mP���U��QJSn�ڕ�^W���;�y�G@��$�}��л�^m��t#�!� [N\��-��)0r%���=ǟO		���R��u�i�U��P#���9��������x|�#m�h�rs�48gt
u��PX�C^,�ͳ��������a'�L$�Q�|�]��L`le���-q�%����d��'d��j��V�F�Ӱ��qk��'H���JQOzK��e��ϧ30wC���A��D�����Y� �i'�5M�����.��\�_��$�6����D;��d��!K�E�����gI�]�^��I��a�������l�8h���x�Ȫ������-y'�k~/�24����X\^��?���O+��>_kC�nV
c6��u�O�q����A�F��J����Y����.G�V�=u�4��|1�
���fp���)���G�u����2{��㯒�NL���ł9��cO�*5ĵ�|��ʰ9�B�o���pH"�l�cvO*��¸���'���Wٞ#p�6�Ȟp��\W��)!�1���C��ڑ��EAT��lp�&�C��v��o�2��mjN͍:Ԡ� /�3G���T�����������a�SK^P���I�.`�
��B��\T2+����LRC�`0�Z�=\�����9N��T��Y��jC<����H�H�ͻ�!�j�l������B�r��tv�;��Ҷe�V��G���T�L���z̊��ޑ	�>P�>�	�\5F��N�̳�~ȞVM\��_/��[���X)��*�7�+�ݕ�˪XνuD������|�߻zp������M��_��څ�W:���Z�`��h0AC �5�����J��vCf���T����8��hm�|_���T�e<���`@FMqh��w�K[��-/%�E:!�RR���:½�=O���?V?C����^[Bk�<��^��1���k���.z9{&�/����u��'��E�ON5AR����C���)O��M�ʕv�1*&"�)x�)�S���IrA��6v���<e��`C��Ħ��ER����s��GM&���"�������fT��R�GׁԓV>4��٢2�U���j@���q���	Xg �U�zu>q��^)U�^�qx�\)��������M�Xg�x���J �Q��]����%V�+Ǜ?��1/	����5�Q(�G6H��i�̌��Db<O�{�Hm��뷪���vS٧��v�@35x�}�V*�t��(?W'���qi�5/T�����+-aH)���a�M6	�{�F���s�NU�o�4`0�kɷ���m�lD2�0މ0�8�,�=k#hE�{ӠΞ��6�����HF��މ�'�t7���pz�d���Ғ��j�1�I
�����v�#����	�������\3Ҍ�y�kǯ�f�f�ܰU����c���B�l�A&N���~�D�CNk�B�`G<jZ
4�.�A=)���h�\q/�Q����(AcE*�]��tgW�c@^�sm0���Jڔ�I�y����G��
��u���USP%��a� �i���J �Ҧԍ�l�p�\M5�7������T�������>׀	�Z��:�)����� o:��>�lF��u��GPb}�"�x�')�b�uW�~�����%a�P��B>D���b7-���.�<�^BԼ���3����%�T��##�J�*���3�|fL�a���A��:.�g������h@���9+����eAZx.POJ`pHU�j���k����M\��㘦�̲.BI>d���}:S����O����d �0A�a]-C��Z��F�����F���O��/m����i�u�a�W��,�\D^H��Dƹ�m�;)�HE�I��i'��<i֜���TP O�Jpv��cg��ݙ�����rn�����kL	3�7v���<�BMĀd���(%he;(&&Z����ߋ�����"�����`s�.2�ۜ�Vˇ~�e���������'MѾ��K��	_��q�T��p�2��iL�P>�RL2��:�����r9�st&�����bdM�����9d�.):����Y����`�!���'w��9��<_4���q՛h�I3��).O�h[��g~��w�	��-e���{���וz��!��k�M8p�^/}�mVڮC߫d�d�(�>zQ׼�|�C��:�ͭ\�Y��<�����uO���S)�7�ЍF�gK��xc�{����s�<����&�&�%l�+� �'wi�O���[�?����W�)�ea�|��9qb#<pAѨ	L6�.��d�[���QB�_,��K�F������Tm�>���X��V*G��m#&��}�_�s�{sF�Ƿ����g���~w�z�&��ޤ9��W�97�)-��O���e2;09�.`�9H�����<j2{4TRJ'�@��^���� ���������wm(��P��@����]2{�}��l;��ْ�p���~�(��!��Nn���� �S��/�l�L8I;7�Y�I�4��O���kD�+zз{6�½ ���5��t��Ra��HKi	'�Ze|�N��Jm��C^j��{�f rd�щ�-Я�q��ٙ~f�Seܰ�h ��!Ý���C��U��A��0/��P�B�:#��=�ŝ�z4������� w���$7�J�u	�@�0��k��Km_�9	��
���;,�n�56����;t���GS#��$죄�x�;� ��5�ۮ�&�ŧ���7k)*@(C��	�HM���ZD��*�X=AUr\�!�go�H�!��W�D���Ec�k9�?��S�6>��s� ���M�|�x(W�KJ���|jp�oU��S�=΋h`�1��������9��+��zaS.������������n�L� �0������*d�󭔦�C+�*=�����M���l4ua�\9�X,g����0ډ�����h>-�~������$�]���<W�H�6���Ī�J�wgہ!����C&�GM�AWT�����\���j�#�}���ة+������:��Ӽ'Q8p_o����[�s�w��N�rruR����|.�8���_�Q���j��o���=/蠓��h�����h�#��{���[�$u��NYbn�#(ޮ�$����0�S.<�#uOM{�t�k�1���2@�d�Ň���X��2S)%
��]����&+5�a��6��,�IB�{e���eOy�q�uH�j�� �q���(����K]\�Y'���yT*�CG����NM�.��7Mm�eQE�םe����A�5��;��>]��=u�k������6����<[e*ᭁ���M��d ��ds�\�q��J\;��Yk5醟le��A&8b� �ö�$�:����+�*a�h���o���2ŗ���~{#�'��Z��v/�N����E-Av���������W�^R[�������u�� RZ{ߔ|�;�z��8�9xQ����	�y��J00�5|�)<�H�rCsJV���V�r���sXPO䚢J=MY�x&�����+����o��m���1���8fM��u�9ȘTo�cU��p�t�~Z��R9�Wv�ŗ+���>|��y`^$4dG1.��r�Ml8�Ү��:���%q*y�|�������o3�Mݓ�6�pc���%�3��ږ:yG�{��lD50�8�Ao��M�좻�`�pZ�Yf���,��9:�ƣZ/(3�Tz�R�8�2��6��Z�|?��f���4���{��{M��� {�	'�L�0��.�T�-vMk��*N������b`َ��nnW� �C�e2�C�����[
߻z�&ݯ(�����4�v17PE�y�Qz� ���p�T�y���= �	�Q��#��w\��"̤F����~gC	2��N-�^���d�v`�Ӄԟ��z�u�V(~����x�������@ho&���Õb���*��6�(�&��c�݅,��aO�7��_<�	���͵�n��vRP�xv7�F�$&H��q��b?�;�dsȪQ�q�/��T	<�عIrNߛk��u�C��W��I��6%��G32c��5�ˇC�qA�G^�恾�A�)&N�v��M��D�B��o��+�,j2!xDV"�l^�,�	�����c����%=��r��NW��uW��fGW7�DʍԛmK�z̸oc�w\o7��ۏjȬ���P`r����:�d�^���� �၁����-;�7�w��Ip23�WZJ�Z�d �@�Z	�83�mIu0h�td�6�ǀ���X�-�l�L\g��@�I��n�����*�b��`��Kj;`;�s��V���nj?|H)-�'��
fPߛcB�R!���	Wv�\�ig� {��d�b���ס��ņ�5�e��&i��]��X̹�FK�G���.�X�.�Ya���MU��*�x���4J��'��Rl�FG���q�8�2�v#�&�� �
��#��{��%D� �̋v s#��1St�Gv��� �-N��t'.Z���{���Z���Y�0�3��v�V�K�%�$�ȗ�E�&���)K�Ȟ��R��.�IN�&�GF�X6 -���*x�q�#��4���9�\���8=u��C�b�YsN��e��n��Z�|�>"[���H*�ҁ��`�����rd!o��fɛ��]��ΰn�9�,Jͬ��kP;�΂�~�m`��56�q���(��U"�eD�ٲf�lZ���!�
��f��������8�v�@��6�U�bL�F�p*��؍�2�i�0�������z`�7%I[⪮ڒ(��]���6m��)���ăx�q}fNW�gӚI�s�bV���[4��� &��|<Q��ja4�+j�Ep]��.�;��zC'�	��/�Ocs�w-�\���tk�v(\$_ܢ��l��[���ݞ%U���lB��Д"{��p(�C��6g�'����R�Kل3�$�ki����ԩ��*(ߺ�J
r���>��˞��`��|�:r��j�˵�N񾆻��ϒ]y�}�yv���0)݃\eP���(*�W�t�4^LӞ���6wWL���ߔE����ݑ=_�{�s���@pg��2��*XUC6���2��1[7�JWED2�뛀m������RU�9��2������D����yL���S��0��nB�$�"vVw|}a�ى���8�aF�q������c^O��H`X�w{)v��{��U�j٫ÃY8��|��;7T[m�]a��׺l��^��`���,���FU���w7��d���M�j[�D�C/w��jjc~&���H·���4eU�K =l�a
�9K�*uv�TS\H]d�}��$�%��A�������PX����|�G���ARFi�믿1��ܕ-
_��G6�B�/��;<�z��&�n�W͋ǍBgz���5G�˅x�Ό�I��f���l��, �K]�D�4��%k�Iޮp:c�}Gs86\?���Y.��>9�g�� Q������A��T�Oy}Z �AqU� �˛�2,�+�6���|Px��z���a�=zH��oӁo;q7�z���nE&>�=��!��6}����	@�;���{k�"4��H���;o\7�Z�c�ӉV y�"�T)��PN��'G��xJi��y�0êe*�{嶎�4wݻ��d 1u�ϓL����fx$�Ьqg����y�:�2�0�xx߳I�tb�1��N�0q��M�U=�{o�-�������Ҿ���l����.d~5?��=%����ӧ���|�M����`GfLM��xS/<f�N����,c5 m��w/�>O�|�P)'	-�RÓ�A?S��=�?���T=y[�^�6�H:K��������@��C�O���g��ncf��"ٓ_�剬wM�u�Y�.)�@����p��=�F01<����"��g�w����m"�&F�<�T�yV�����q�`�����)=��F��e�����4eҍV�=�
O��'��Toj0yw��P3Dp�R�̒���ؠ��8V�	|ѹc�|:�0��XDzqݬM ��Y4}��;�қ�������A3�W�����Ca.�߿�5��#����`������k�9��cI�*$t�j��-k��*�M~��u0ދ'(1����Tŵ������>�_R��+�3A_4�8F5Z��[]��Q�r�8^��:%%�_:�c7��s�̀pK�i^A�9O�S�N0�:n��A���`���8�w�^��w����4�04�y��z��;�7��������C,��, R;��O<�����8~I�7��=�0H`��C�R���i$FH,�Y2n$�AэS�~Cvf��Ւ��&|qxu�DWk�v�H��u�B�X�D�����"��t����R�}��XX"�>Dx�yܪ�gسt�(Rk೓  TևtC,Y ��Kb���	��=O�9���С������x��fu���s�w������ij�7��CND�Z�sl��_#�Q��ȕ�͆.�6���J_E�q��p��V�e?�p�����������@��d9�i8�d���������v��GB!_���y�^�F'�����.�J��t�-�&��H�z0��n��%c����u6NH�D��f|xIz�=w�2�\�8;NFJ���O�A�y�#�Fs��&`�l��e�טj�ƻ��\ڗ?y0]_Se��P<.���2fi~.;��/������eJ�E���4>q��y�Lm��ׄn�P�ڻ2x�T���F�9�k��e3L��6��Y�V�n�k)�4��|�hSX�a`v��'��fv��^�ZQ�P�r� /VKj9j�@��
xa�Cc�~}b_��B�5lC�{�}�M'��l�q'ecK��<�4D`}L��I�Ђ<!�8�%{`�lѳҊu�,p9��G/��m�����T[�2T:�6���݆(���A�BҼS4�	��G%1��ާ�ot���K%,w�IO:]3��ĩ,'��~�k��)� ��Y�[[ ��dG�����1��]@�G6���+��Bc�r�sLY�t0v,��!��l�Ԣl��{ ��6�.�ec�VD��z�O�"�6���e�Q�v����u]��8m���FE��Ѯ���b���7��%6��?���f�VO�U�`ΐ��&K���U�{�������^<�͋���ub�Z�����*��ZvoV��tYFw�אS���"�����j.i��;R|_�y����f�H�3����{ʛ~ϗ@��5}���At5��{P܍\�(���m��jɟ��U�j�?�纃<~d0���40߶����#a�x�%'�ꤔ�i<�ͩ�MSa�kLY��@ځ�׮EY�z��Z�Bb�]�0�,���b�\�(m�w�D.��T���r-V��m�0����MP�%��dbn�Y5Fi=�U<��_:�4
9)��N���lP!�tox :��F\���ǭfל�@�(9���J�{�Pk"klpXw�݄�>AHW9��ő&P�mW'^�Y���2��E ��އ�g�A�a����~��'��u�b��n����������d�5 ͳ�V�u9Ŗ
M��`Piq�i�m����� ��cy���n�yѐExa{�Ėƞ�"=��o2���>��~���{�<y#P�A]�oL�c��6ܼ�,,��r�l����D�:sDF5*&H�&/4b����
�����QS[W�{y<�������.�������
�.�P��½AF
#86�^�Y�����"q���tw��^����ڢ޴�r�@s�՜�:�[�=�J���,)��v[�����Sq�~�m�^Wm�q�!Hڌ�У&��>�<�G���X�t4W��Op����
{��)�y���JR�~ۛ)_48�.��r�\����>r����~���F�����.�����[I��y�lJ�5�~n�ƺ�>�ҽdF�,=���S�Y�k�O�Ij�5\	���_��RS�/Z@_��6x~'�$�z�q�]j)hG�P qf��eZ1׈�]�v�7��g��z��91�d`�����Y_���ḩ?i4nf��n
`�tJBv1���x]u7���%�	۫�Z��%R�.���Ϝ�gad�},���`�Nb�z(cߧ�%��$M,����#�nKR���wZ�������sٴ$Y9	�%��t�c[�um6����o�=�M��n�����`b��J�o�g��Y��7Q�[ı.f���Fl7�5�`C������x�u�]Z�!��}���n��Pu�xK�=�W�L	٘+�^��>��z���F���׍�%��ɍ�v�t.'9�..��z}.KQ�ݒ��,���0�8��O���mm��u,���u4�m��]Y)t(>?��=��YY6���{���{ߙe��Nr�+��a��N��o��c����a ����B7Л�a���jRJh�0*��6z!�s�����@�]�Ɍs`Q}7�w�.(�r�PO�o.�7�Ln�鲲1��5��1[�AR۷�5��Y�����I��FJP{�o��d4����8n%��i*��i8�M��d�x�}���g[,�a�E?ц��?~:�
7vUU�"W�k�ƺع�`��K�A��#ػ,��m�V�#���U���x�X�֔k����K4^;�6�ei��0�Lq��4Ռ�np��������`�����鋽ݭK��?�2�n��*����FS���MN�t��J)Y�sj?)�;8����.A���:�l�((b?0��E�7e��.�{Ů�+�)�#K��^Z3�:�o��&D��Z� �����1�wf��9��� ]c����M��E1��j�o��~�0R��?��΢"$�ZxdV�vG���	��T,8q���� � �R֪1�2_�ų�8j89�js�>ﹸ��\�c)�ŁB�%�2܀h�j3L��$Rl蝍"p�(#H�۶	*`w<4Ew_���ٝ��pm�[�y�r�-5Ե����I�A��"��IM$���.��m_�13�a����=�W�>΢�E����Ȥbn���x�l��a����X�#(tZ�&��⮮ ��"o5���Y�~�ᴵ�otf�\7�V��{��XC��8X���q�c�|������'x�F��9��4	��m����^�9��"�yO\%�r�ޘ����%f�5�"���>�1[�1�$���^P�֜x�qτ�Tq��:������&�ld$`d���SR4�^!�8�J��5�������,-��y�-��Ɖ���\�C��F~�LQ��C6�����T�8����X�We���OK{\dd����b5�[n;"���Ơ,���Sg��V�{�w<�D�Fwt�t�ŵ q�.�
r�H�{��j��&;w�������1���Y�\Yf��=���x�Z��;��߽1���`�L��q����In��q����j����������84(f���������u(�@Τ�E)�f�kT1P��^HG����|��m�}�tࠡ�*އM�B�ے�5,3epۅ���|�Vy�=Ƥ�A<:/�����)�qOZ͞�g���4�!=ծϟ�0C�9> pX�� ��]���/Z���e��w�T�g u�#���ΌY׾C]ۤ��׏C[���{f�Ūe%L3p<����ة)d�a��U�� ��~�jZf�T�_'D[�E�),��)��@s#.+�I��"�:��)�Jʖ����Oү�z��O�O�#j�a��=�`B�i�T��C��8���]�l��r2�������EP�MxF7�]3��2���P�b�p� �o�W��z��]E���Ke̙3�����P��4�����I�(�Q��n��a�ު�5���0�7⠊�e�G	u>O��G$�^��Y
�*�6�Yn���iw�k�E6K��cP��Vv�C	�0���¶��\;f��Ԡ��+�_���C#�1fS)Mkڸ��ۘ�ff���b��HT�l����ˋ3
��UwЍ&�nN4k$ޫ��)\L��JΔ����t��-�X����_�_��L�*�FC�+:)w������Ө�m������$� �hk�u�&h0_�N;1�ܟ�S�&���8s����Q��l�*�£e8 c���/��䜽G��������*�@�������N��?���ฌ��5�jb�:K�6�B$d�)�y[�Ӛl�`� ��.5�*3���z���|*{�\�1%P �Kj����Y4y�@�b~5�۲��zU���|��S��z1U�x�l�;���Y��3~�kT�����?�L�]J4�8�0��c��S6���}�ƴ�K!M�\Śp�$&��+8�q<��)��XR,�ɂ�x<�#�����Z�KS�VL��wU~��b�球��'��vg��(TR������U����{U3�ǒ<� �ע� �j�źC���-�q/O���J�K�Q��%	��x���҇���L]�w�TMD^C���Cl"���zkϞ�_-�m��EW�\���SO1�9�{�S5���)1H�/��s���H;�/�hT��Q-��4H�xWf�8��;C��<��uM�r���*��{�k�5ww��}X�"���_7����bF
�����L�A�B~��L�4ѣ>�HԹ�%6=���g,� =���&��a���EQm,U��������������o�9y��7�*��H����!`GU۱tw��04p�l�1��XG5C�X������4{d��3S���W&�#�"軙�\��I�A��:c*�����:��~�H!����{ٞ���$,9�>��><$��
�
mYӟ$�+�3ҾvT=�y�6�i`��w��g���Z����Q���u���r:8��%:�vj��j���0�:�~#��a|�0�?�89��
�{f9l�ؚ�6�<F�u3�:�L:LjQ\.lB���SVd���Q��\&���40K-�6\��������8�1l<�_��
>�8��G�\�;��	Vx��s���A����T���)�E�&��D�Cq�=&���4��5_��Dl.�LW�c�Wӷ�u����Oi`4��'�ZS�ƶ
̙Z�)�.�J�vL�8E��uSe�	1���R�˒~;7)�{��٥q�{��eP��2'q&���� �\�!�B�?;f6��^�]�0D��{�%�rH��bsS�c��f��v��F�xʳ��x,�EM�Mx˷�n�I
��p�8�4a�o�%�+�VPM��~��U������s\Y�C�זj2�3ՋzUfm8�}byZ�%u���XY��(P{{l�o�ynW+�|so��ڱ�pI��nb�	��D��u^8=,��~)��?`pN���^]�꜑�0�J�.��w��4$�M��ʌ���l
m}�T��A�%��8wދ��\�=����s�HLʣ)e]��|*�z����/]l^�W��w|P^1KHN�̲S<S���5�D&+���}E&�U8H��.Nfϡ���^<:��/Һ :�R�}��s�4&Cv��8ɞ5�����FJ���&><>�WC�s��B0����bP��g����|֩�$���-` 7̐eq<q�fu(���b6ҩ�>�۷���K�/ov
R���į�̑Fg>L���h\�.H#q��,8�T~<�P�D�1�w��B��^?�N��G)�����!��՘%��~3�!���Q��t��,�ƪnn�Q����lf���[s<дQ����4]}��@��{���Swl�4�]�hSh8\R�������/����5�Oݡ<�k�2K�.�H������:u�����qF�n.1��j7Z{�T���k�(��Ln�3��:����h(šmp;����]L����D�'�e��\�ʬ�2m�V,ٵ�5�3_�v4��/Pq��<>�vG�N�{8	.�T��3EE��M�����I��Uf���R+8���O��|]�57Rq9"ƅ����M��ᕒMw���f�M�5�N�^��_d�k<'���e�AC�Hʇ�L�V&lƀrBm��������o��x?�I���(�_4��(���Ǹy��L�N�9Vo�����~�&�îN�k�N&~��}`q��{t����|>��D	C,`�:��;�3%��-b �p.tۙ��y[xx"P�>~���͝]��p��,��"�lU\�muG����RI]zc�^��;o�N�oɡ���X�,����`G��jJ8|� ����9��`wOAў�&��M*����"վ�1Q����(׃�8W[��	y� ���4p���u5[����m<�,�����ǚ��<Q�;Jz$A:����^��3QO�U!�[|&���?�{
���X�3J�d �U@����U��/^�E��F%�I�m�t+6x����<�bO��S-�s �:������.���y�\�F݋@���Wݤ8�F�����^"��=ǉ5�V���`11�61[>�	����4�v���莯�L�YdW��s��@�`l����IZFD���O?�F��!��Qc>/��-��d�|/Cn�4�Y��~�����ު�%����ܹk��\��qAꘗk�wy�����g���&���҈�p�]�l&=�u~��ww��Xxϟ_��ʒL��G0���4o^	��4a�1\��c/Z�R���@�I�m����2�ڏc�p�l$z�����*�<��zS�c��Z�ۥ��*c��x�6+�VA�������]$Ɉ@�je��?�������a�#��`s�Hc4T�b�`P�vK��h��p����b0��A�cŲ�<�C�g ��tw�*�E'Vk5Y脥\`��N�H{�S$?�����P�G#�����u�Mw��#㉅v�/r���x}>��)�$/;Ħ}
a��nJ��41�ߋ�5�:;��\��6!/���k擟��]v����$^7�K�k`Gp�^K�����ī#�w�|��z�f�<��4��Q� ����t�h��K������뱝�mv-����O�[����J\֦j�qe�W4��=*Ni|����M4?�L\t� �F@�S7EM+��]�=1-"?+�>p( ��V)�h`��|d"��-��t��p�������/�^nV����R�<�r���3�I���cv����3T�f�f�jj��7��/9�K	5�ㄱ��i�~cd�t9?�5:��=S�� ���ˍ����=�b��"���3��$���)�l/:�)KM�w��6�*��hś�W�E������q�����̊�a��GPK1\K��j������+���@�%���}��ŮP��*l�,SG��_o�rT��xFO&�e�k>M1�������$#���x� ��irK�i��:%ǉ��(P��"�E%,�=�ׯ"�~���du�w��<ܝ����b}�^�=�$���SU���yQ��w�¡�����Yt^k��@ng�O�n�K����b���/�������)V�F�h�L�wqm>?��L�A{�e�����:4��P_v�/a���f�����b����?|�X~����M�>~�ݻ��������ԍ��I��0+T����fyX3̞�U
�T���3���� �羞�0Y֪��9��ɐe�fծ!�	�6�|���6��ж��u*N6�cIK��hhk9�8��ם��Ǌm,�m�R1�AnM3��A�C�K�D��&���?8c͇��]M=⒬�����@	�`�z�����j��n�k��]V"���f�.7N�����t�(گ���[�H�.fu�\n�}�&�������}w�~3���W`�_�H��\7�Y�y�����7�6���pKqx@�V �}�"�	"v�)Ze���?�x��=.�X;�Y��f�r��b4/�����U��:�[u�Blq]YNL����{PHƪN�tO �}��G����^T,ݰ������{+����C`ԁ�{P���_5�>e��f|�;�Ί��)u��Ty�����ٷ5��@zd�0WQjdT�����H;������������im�~����M�.YC�����u� H��<-t��#,��{�UN�!��ou�o�N��h���i�b���>Ӂ0��>��-Hd�X���!4�σCy��Yk�r����#�Z!��ּ�4�S�&�c�{�;@���е������T�gK��JtTbx���ɒ*�e�����!�%��鳚���,v�;���𹑑6��w���j@�Y�j��*��V��d���d�۹��EЯ׎����%��7ގU�\,_�)xG�4T�A�>nH`:��J3h�Ϙe��\�I�_n)p�S���Ţzg��N����͘�x`մ�EC���q!g�����h����A��c|d.�kӠ��*�̚f��)-�ۙ4�ٓ#����st!�e�O��0� j"�KņS��7����E�Π����7e�j;�כ�0�#F���&b�!���:�p8+����O�M��B+��[�+{M��L�Q%�u6���7a}��53�,\ra�2yS!w��w�d��b���n�Q�_��u��3�롯���A+�Ը��=��6�L�z��H�7���-L\��~��OA�rύΩ2c̃��\���-t~��[�?/�����o�u&�	���[l�t�〴ݲ>ST/C�D��rvܰM�D��K��)~���ߧީ!��ڬ�_�Y��?�?�ROC;�������\�a�M�\���_���ߊr�.�Gi��-F�8U�;՛���E�8&K�Y�)T�i�{�4Yƾ���Y3髀j�B`�s��j����bsX����#��\���΢�+�'?�^�s�DVWH�Y�׷W��:Z Aw���������:�Nm��44S�-� A��ry.z�@��;�����AX� �|<G�*m+�/I���Olq�o�5��G�H�$[�tvsD��_^r�r���+��@AZ�����#X<P(�Q��i'�)�����kN��{v��(s!\.�6��(�ͱE&�������ǉ���ʦ�y�4L���G5�o+"j\��CC�V;���5|��������{}�+i��l��I�ޒ-�k ̡e�~/x�%`�G*�������p��u)ֲkBM�/���Z9��!��:ߥ����YK�R�������S�'��`�E(�pl~uƸ菛���H�!�C�t�}W��V,6�	3��C ���}�(�n�ΕH���S�ʓ�;ǒ�sFQ�_�W�Y��Sd��B��'2�����Y�Ƞ_xn�8�K�4섿RG��3�5_�y�1�����T)����ܫ0�-��Q`�L�]�{4�.���{� $0�@���>x���-:�8Hx �
�]ⵝ�����j��cp��{�F���:!(,1Yrk2�i/�~<B:�&�?��Lenǒי݉�Q��+�:>��Ǻ<S�
%-9��<��Fut��Ŋ�K�+)Kl���GY��\NҫJ��'�Z�����6:��ߢ{�2v�s�b��L��B��3��W6�S�����T�z��B��%1��]���oB�B��h ��U��YuH-�_��A,?�uͪ����#��`m�:%XǨ�e�?�k�av	Z�q�n�Y�-N��um���{g�O]�GbD�AH�:c��L-e���%���FP�A��`Zt����N �X-|"n�yDc*R�wC�$���q�r���t��i��R��*6���cMч>?e�N�Ys�z�jW�MS;�^�!.g5�c�ח� 4	cG���M�1��wlڟ�����\��	����Q�?����5n0��#���^���������x�Re�|�y�y�r��1��L�^7/l�km֔�YX~m
���kԶi
��pP��&�*J�-�[�[�a��(S�*V\�k�Ӧb �
�>Ȃ�#CD��z�{�R�e��t4�ǲT�Xf6+gޓ���F�2��&�w�ѿ�\M�'T?�Wa>k��P��8כ�� "2ʸ��!���[y\�L��5�����.�� �X����/�� @��<q>}��;��y����jθ�5,��Z�������'/)g��U:�U���WF ��51@���z��$���{O7}	�v���KQ��}ի�M���'���_v��&.��6"�;2����K�z�jHO�N7'\h2n{�\x]N��TZ4�ƒ�6����6�`�gF�f�ϱx�i�#�^@����w�蘃���������#�{��mQ�4�>k>_0 ���L'�h��
���V,��	���D��F_����/�����?�Y~����`�=��?�9���v��>=��S��'��15������q.��m� ���g~����#3#����SN{%�c��5c�|�8�V��ٷ'6�T������c�`�?�)��*m�����r�疘K̇{|�{�s�R��p=p�����5��~�k���1��!��1��u���G's�z�*�8��N~��yM����X�ޣ���x_�sֆ�PvN%�q\;`�ͬ;˫H|-d���(����",�A�m���X�s��0����s~x�U�b�0l���jm\V]԰�^m\ԍ��o=���Wu)�=�E��)�kIa�
Z�M�":]ca�1:K��w��+�Y��]bq�@�8�:�<�izƆ0�Z�I�� :�I�E��|��<�aO�; ($�������w��(������~*���=���'6,��	�����X0�$��.V����m+vR�B$���)�'��}� ��SN�,3�g�od$��Ս�,�v�Ɠr�׭�T��w�E�~QG]%����8��%�0|&���uu*�J�溘)��˫J�؈�:M�T1׮#��VEur�v�|^�*a�%�㯏�5���]mg���zg�7�0Q�&_�=X���9�C: bMvv��P_2�zϱ�G7�+8�
 �f�m�cf��6�0�`�瑱��q�r�%k�����,�G�9���	���d�:*���4�Y�R^����@m�'�}��H_4�*��h��-rͪY��٬<�[���G�ϛK�7�פ����ڶ{op�ٵ��������E���KM<�P��p��7x�:�jw���8�E�-*]��H��9�l��cࡲpF@���I�S�_�I�ۿ�[|v4���U�7�A����l������_��n��7�|�Iq\����*5ԣ�~����������8'�u���fH��>��1ex�)��x���ه̢Ln��R�R��^>�����葝]��.�*M�n"��P�E������\^OY��A"+����|���h~%S���f��M8+�[�y�y�~�,iLݴ��%;����!�4E`	]TK���!<=N���������R�U��9|T6K�b�!59�m�
Ǭ�|Q)��e- ��^K:y*�wי�!����n��Gwj���((�r�Y��Gr���4Y%J&���%|?T����k��k�VA4��ac-1��WϲR���X5��A�3��Wm�1�Z�2����m��X.r��D���{�*,;ݸ��z\o≙I���ԓ���	��H�u�B"S�s-j@�ۺ$%���Y��ɹ,W�@I+�^��eO���-�~�:W�L��?&@~,�!��OG�_O�I�S��eׂ�$�˯���z�R8�۬Idſ��ׇ���)/R�)��u���E�bdsX��6�lU܇^gH�	�����P�A��� �&`�cs�@C�<�'�e��[�e�������>:�H�g��;�V2�i�հ7�����(�c|��msbvQv��+mQn�1U�r��R�u�=��iu-~2�E��>�����*�	x�ڕSfq�����:p�جQQT���,!kU����+=_s��0���^��L�x��.�A	j݄�>����ۮƝ��zQ��|~���u��)�>�D�K�D|Vi�>\����6X��wod���"#�Z��S����7pxM �|�7^�_UFT;����n�]�f�V7&O�V=]1(`�������M��h[Qt��񧼁 ��OkRglMRDU�RR
<�_ڑ#���q��'�<t
8�@�s	������w�>=�����G���"�������|�m�w2=z�o�MB �t�*S�G�ʇ�<��c���ߒ��@Z�G��\޽{_>��$�G��i<EP\%��MP�(�3`�.0p-�Hp�L��awq��~���-��s< k
!���%���d�wg  ��IDAT_Ш�k�i�C.R]�.��;�lz��h���Buy~V|����$�Fx]��n�k�O?�����=:�/���3\ҳ�=��Y�\�!�[��ά�P�(��KK=~(Q����߹���z"=�1���0���ܪ�3G:HW���cu�p_��K@�[�Y��&��>���e���>��E�'��vi��({�69��I�ڌ�]XzR'������W��(�  ̚�i�vDddՀ��j��bLw������ps:����Y��� ��f�2�+k��JX�)��1\�3��,�*?�2��Z�f�TÿSPe{�1��l-Q5��jZ���ؗ�h��X#m�W���r9\����0Ͼ� j�wY�ه��:����0��[+��>)aF�R�mB��5�����������4�ꥩu�B�*U��A��E��5�u���纋s��Lӕ!,�ACz�ѷQ�qS���;^#i�a�r�=i8�U��Oz��^��m^�i3���X~��O<����Z9�E(:�h�u�y[��s��AOCva�7�s����<4�`8aDϸV��@}?�S����VZ߮��d^�,GT�l���p |�w!t�X.�F�N[�S�!�Nk\cqw���z����r`l�Ez�<�qhO�~*��	���׏���}�~R<8y�cb�P�ق�Z���8�������B�J��'\es|x�[�aq�t�O�����i`�-Q��4��;"B����ҁ��o9�5��j5j}�_$�D/3�c��㐑�_O��3�x0_�	5��'z�{J/V}ZG�UF��Hv):�0/�P��5��%
M.����
k�v���ѻM�|�v�c�pbWic���ڈ<�RJ[�����k��T�Jb��s#��~5|��TW|��M��V���^�C˚a��l���l,�r\�a !����Q�=��hk��U�8D9�)�X	Pm|]��w���1D/���^
������=1Ϸo��t��mhѪ�Hp��P-ߞ�c>��:�����"�.��w�6�?]�A;�Y��<G@҇Ioj`V��c���Z������eh����B��N�ϛ�ɀ�n^��ݳm��J�ghO�B�쐾8L��Z(s@C��)}|������z���=Z��3�(�%X]CK�D�7�J��q��c����WZ�{3͵����[�8�-��l(ׂw��Wm�L���1�R#C�D�>z"]m����bRtQ�����$��m�
>"�a'�sG�.i_���޴Ϋ�s�!�]s,эb-�T6�qA��N�sF[�5j05R	�d�d����ݜ�Z�/�&�%����B��*B�X��`!�~��ۇ�Q?������V�|K����0���k>МŲ��,���O�&Bf�Ui <S�<3A�]`o}��d!��N@R���秒���l��0wiۂ���]ވ�"����NŜQ����@��Bch�V~��c�05�?��c��!��u�>�� ��Kr�3���"Qu(u��k�������"N���,�{�|����e�Ӌ�gHTUR8�/�Abm8�'?��>�������F���� RQ�F�eh�띥����-�q�����1�H Y���мL�Ơ�*=ku�x���R\A�{9��ɋ�flL�U�S�J�D�Ё��""gЪ��=��9�E'o��}
# ��һ<�XsH���P:Jr�D�W�ċ��&S��0�bոw�k�o���� e��5��|�1ͬN��	%+�1j؏�j�.�^�B���je����2����߂M#��K�}�u��X�<�-@�^\�U��<s��:���G`���u���ΐ��o�]��9	�-V��U�W�`۰�4�,5NƩ��>K!�@�z3 ���kp!�Pp�.��ʎ^��ɖ�����^℣!1[�T��8t90�9�$s�p����}L�;^#���=�z��X��E��pX����T�Z��=��gR���HZ��zp�:P��%�3d>��8~�ˌ���駔;��O+g�s[��q��Z&�c_�yh"Q��`/ң�$��$�7o�D;�}(��~Bj�mi;���)g�un5vG����i���lr�Q��JUw�-�K������T�ϓG����a]�tVc�9�aHo�9���Rn2$݂F=�������z�\S	�]�~%#���l�51m7�62]�5L��Y�o�#"��䪟V�6�<ٖH�{t��v�k=���9.	�<0Bs��0Ta��Nh�����H�9��<C��#X��cZ���ђ<�4��Sf)Z�4CY-p�Y�tu��3�Ԧ�72�R��J��cyh"Xl0��lt
!]���;"�K���a��Pa�G
�pa�O�S
�ڐ�#%x����ft�G���P�ϫ��t��8����d��Io�Y�J[�15+��6����Ɇ�;�#���D�
Fߏ��_ߔ7o�2a�k���4�ǌK�1���%؍ ����m��u[�2�&ч�o �_��h�������},o߼�C6��_hH�وZ�׉�%��9J���==���p�ҵv4�E8��KB<(w]�g�7r4��X)j�H�X�S�L,ѻjI߅��^Y�`R��.E�/瞆\s������c�j�lޯ�����lc���в�Y�Sb�ɛ�^(�[��|��L#��(���e�/p�.���ե��G���ɋ�6b%�Ĳ�����Y�����^,��AY��d^G����0�kӮyA�������i�K�d�q��\ȇ�acʠB4�bPV��rs:UHL_B��2G5ԅߤS���N�X�㶧��>E�׳3ͧk��⠰Z}��k{MUa�q�|��ey��=�(`���N%�%C�2_�w�Sx�"�[)~�ČX�
+�!�œ�g��-<TP��0l� سRk�-v��P�]�N�����w$�[�B�5�Z#�Φ��Q�Ϻw�QBwme��~L~�zA�R�MxV+6QKF�Tq�\a24���Kf��L���\Yk�li������v�MIl���G���碽Ū*�l�]�2K�W�J����&i-�O�Y[o_� P������2��~��Wrc�>�hZ��f�@��u=G��!:q��2�K*�m��V��8e�9z�9Z��}.#�{*���n���՞Xr�S�ut΢����)�I�D��%W��d�&1�J�xw�8��i9tŦ�ʘڀ������#�Va��c��`+e�@�~a��XG�9#�z����_�b�Ν3�V��������8+i���5�-��	(����Wϑf�Z�8
��&�o���^���k��I���9���	�����<D4?1�r�b�GXD��jD�4K�ɺ�,��G8)���}� �Ђ(K[�1�7 ����>�p��=��҉B/'~��ç ��)����(�}��q���Ko%ޡ���a0���A��yd�(��\EW,Z3���2lK�Z������ e(��_l��B7�eSC?q��]���(t^�w��&ץv�mK�f��s���z��2�䎒��(����224�e�K6����x�+�B�e���wFJ��j��y�l
�3��*N�/��c�����_��^�#�C���~`/��p�z:?Fbv��}n����Y%����1���^���RNY�4�W�ZHs�G�~-��ڂ�����w�k�zg��2v�c�,<�-�<���u�P+:G	aU3W�UI��9n0���C���[m��-��Id�1���F�L�,V#-I�͕&�F����ҔJf�?�-���S�y���'d�6�MY����J��)/��1q��<��"�ڦ9����2��õ�:d����)�t��/E���.�%��j� �~Qo�%��0C�*ŉ��g�O4��Q��6�{�٨����b-Xm�>1�5� L}�ف/$pQ%E��i���u!�:�1����{��C�!z_ݤ'���?(*�tű��A�	��H��OJP���3vAV��p>��ċ��LSRo�uY������g\[󐌔L"��B[w��{�@?	ۭ�p^B ���ST=�`��"�ɸN1vMx�59���H�������c��A����q�>f�11�$�*���w'��ݗ�f���	���k�n�Ҙ.���&���1�+�������V׶��������͘�O�XXy3(	�N�U�xj2�F/�Tu�2ɄL��+uc%�a��Y���BV�KϠ��������^<	u.��O�՘�JC��� އ��H��O�$��һYU6���ƶe�|\zf��J���h2꩘<����̔��W؏��z�U�بv���۵�����_)��.�pUתr���W�~�p�*�[��Mܖ�z�,Xm�iB��nf�)`�ǺR5L!�(O�!�|,�~[�ʱX]n��D��P�%��mMFAS�_�\�ɳns�H����� ��:/E�B�5��]�$7$���X��~�]a���K'�(V��q�A
���)J)MΗ�V�K��61�6��S���5�3�4T�
Y�^Eg�r��l�2WHep �8o�K<��a�pЁ�W�V
&�Ǯ��~��ג�y����ʈ���<��_gHWc�/M�a1f�k�}Ye>|�P�qs�ͅe�
"���m����)Ú9�jN����pg�%���dh�W5o�"�X��0Rߍš�z_�*.��<�VR��+���m�z<��!�fL�	�gS�}��������%z��ɝ�4PVvghop>�t1D/r4�rz�,�;Ѹ"q��%GQ��cSx��3��k�9�җ:LNJ`�o��>&<��1�wl8�e����݇��um��㰁��K(��=����]�]���Ŀ�mRoe�=Œ��2�1�u1����ܖ�} >-�O����B��2�X��	�G����f4���6��6������u:uU�:�3�w?��������ݽ�O�At�ct��Eb�@x|�]i%��t�:���h���&~�;sn-�]?F��4�5ۺ��U@�@��h��>�wR��ۮk���h 9F�1E����!�
ߏ������S�tLΨ���^P��<m7��	�LU{ DŘ�ܜV�4���H?��E#��;l�nh=G}��!���z�5Sr�������o<)wͬnu^~���o�-����l<$%�ݹ�5���K����tzg.�.�� q��Ȉ��3'�NLюRHc�'�������Ǣr�fեx
=�aȓ��0)S�Ds������C.����4���V�tzJ���ȭP���!^Jk��Q����횝�Ŝ�۪9��LE�#��=��f9�}��x��d�qm5���{yՀP�]0�7���f��4�ZIj�'�X����������0�}]oݪ���9�c�}΢"oF�qC@ᕺ�����1m�H�V_޼���ٌ!k`0n��
{�R�O���J"�'��a2֭\T�|z�QX#�n��*��O�mU��rr�
��j�:���8��t,�џY<Ğ����X����r�2憮���8���@LP1!*�ҺZ���!mK���X#������1mCb..A�������s����B�l����1�p",����ɫ_w�4�����H�x����ρޝ) ���ՙ�IτiO<����u��K,�p�b�t�ߎ�CPO��f��S�2�2��Gڐ^.ǀ'f^g�
���.Vx����2,!Q�h���Ю�f�(2��G?| ������c�4����V��w"��:�yyBw3=���]������:��q,q��Zg�G�''�PFr�9���2W^0��݌�{��kߪ<�	��sz,b���2rAU�A2��e�����X�sr�}����gS7>w�H�<Re��������`�Ix���421���n0"Ps�o|�Bmp�=m��Q�MJ=b�݇�����1�w�w�R�P��
J�j��Y~��Hh��+x�������( �/��yI�W��԰6�H�?�5��[�<���������mmC��8�ܒƆT��!���>l��{���'a���Q�Lkn[�l�I��������z�w��29cL��t��S��n�����1m�Yu��5�n���zV���k�DM�YKm�����`eǝ�L���qc��n�M���w�0sU�,G�ml���8_js/���9jȷ�eس�jj�[��P��+=OʥV���~�S�G]ʰ��7�C.��=��B�?0��k��V3P^7�����x�����4a������q���g�uP�(0�y�����Z]���U����t�\�V����(�Q�f�K 'by��l��܄��rׂR$�b耇c\�i96�)�8Q$P�}���p�ǥ���w{�ڠ�^�`��5'��,��C�3���b3đ��zꃱ}z�oxBo�W�e�o�s��7�����5�~�%9���C3�����ƻ�5j�wN��U�I�os#��5re����G�%g��O���Z]iʝ�JͶqLW!�Lvt�A�b��Q�a� ��c�8��L�b{.��[�T"b���OYI�����t��_.j���'&���]��k��6)U����po�!�hq��XO/�P�9@�����[�8פG�h��hLˇG������q�5z،��HI���NGʔ���R��h~V�E\�S&��{���{;�@�[��J%tk,N�M�,/��u)kz�N�8Ӌ��|�j8�s������](�|R��50ג�K������Nԡ���Z�^�*��)��2�=;������;���r�����B ���	"��R'���������=۸���y�,�&���iYU����L�؋�Γ�}����!>U,��<�)��Ω%
�*{��X��^�U���:�܂���F�ڙ�i[�"�+�٩��&�����:0K@a��'Lk�)>7�y�����9eb$��?���)�O�"�d���լ�9��Z�A5���0,����;p�JQ�76���,f c�0�������� k9� ��3{��úm�����%���%���{���57#��0��OO!<�D%�H�����1����.<.��Z�!=~g/X$���h����ח]w���w����!�f����\�-���bv�C�C ݡ��]a��9fcRcz�s���bdY�^^����Z��!�+������bq=*�84Do�����"K��J��2_?_�\ǁ���=�'óF��B��J��V_�꿎u�IM��W��5�IɡO��NF���ܮY^i	��#Iz��k�]�.�s'A3����5Ԉ�Q<̉�w�k��tH�b�ϣ�����Kp�������:P��1�]�N_�;���P�P��w� �AX�io��ZD���V�^�(��!l����	�6�Za��bH�|�OY_�� 08۟�jh0�ZI�5eB+�,��z��ga�
�t�&5�]2�b�5�/i�$66E������Yi1\�g��-��'�!|�:���j�γ����
�X��dc6	��Ճn=QWx�K�.6��aq�񘇉�������	ä�x�Ww]+�Sj}t�P�Gc�U1��iѝ�sP}���L��U0��r^��rD��G���j�n(�!#��8M���y�P	�B�M�y��ɨy����^��"�GI�"�� 5��`Ms����r7���R=�n��~!�?uC@#ԒX����z��4e�Z�B�]JK-��ژ����s�r�+j@5]Iυ'J����u8��L�
U��J8j��q@8%��n�Ʉet�<t]� �߶n>�W
N�����z���Ҿw����D�����t�rm��f���^�ǟП��y��!͖a�<W0;ܩDMD�K���%[�Nzx������/(pq�%��U}�m��F���8Gݲt	�w��1���$�D����(��Ĥ��"$r�W&������(�[���Y:�?�uL�����ˮ�o3ε��U��"~'Nɖͻ�}�ډ�ΦV!�Oz�U��Ɋ���B&W|�3f����:0���cؗ9��;�A{�9���	8z񥊱��UG�N-6���Fu��|/_�q�_�	A���1'W��C����ǽO���'ەz�.�'+@-тZ��DǭJeϹD�ob��~��T�@��'�C���'m�Q|�4�+�Bs�{�D��*��9�����ݻ�����D�g3�`T�*ϗ��]*��7uo�*��U�}��cG�f0t�&������e����9����,��.]�FѤ�R�]��5�i�O�걷��jC�?[wt��1�1�����d�»�Ø
��!���7*�0��'�;,���ݧY�/��2{��uG���P
��H����8��zm�ſ�"I���\L�$
׼do{]>4Fw9M�q�Z=G8=dr��,��ܰc���X��k���t<{2�Ui�͸squn�ّ���#i�h 3ҿ�nT����$��MWңv��U@G��`1��/(\�S]P���G�>8�T�%#��$BT�������&�	O���{K�9����EMťU�G�땺PW��^M�iH�=��w���}d7�	���B���k�R&C�z�`��S��� y��n��ZC�������t��z��>aER���?ʎH�ͪCa��#0xV|����u^�׆ԥ�6��)`�<۞(��{@y�(KK�#n|�]�+��(i64U�k�o��@��a�D����K-��t��׮4F�όi�	�k�=��BF�dh�厣Hףկ���Ah��_��D,��֚�9��0�_lO�o`p��r0E���t�E����6qw0Mj�p������d�&���o�F�@mA����Yױ����0�%��*�0\a��O���#��.@n�(o�>�b��x��J�_�,s��w�E��O���(kJ�����T�(H������^U@x/[
s��������a���$�3��"���%E���Q�z���BQ�!���8��P�Q?�~�.y�^쵕wŏ+��U7�+�w5��;缃!�rBc�UnΆt�����ϥ&I��lBK�}���x�s��a��3���yx��2>MkpX��!2�P�"��/<@�Ѣ::�ؓpl^F���W���J��Өu��R$aH_��"qm���K�z����)���.�Ϯ��9�lR�e��=�-qb�b!zXDao-WӶ_�����'jjȯ:�Zٔ�=��$�^^��6%��x�zb�7�<���6�<��$���0A���qی���8�. �Jf�5hCV�M�����@���*��	RO�7�k�ͽk)3ƛ������:�̓c�kRk��U]|�s��ѳC+���g��DSN75�H�BS�c��D[;l�k�5��YO���0v����R{���7�Cra$�������W+�׎y{��9�[�2�L�Ҷ�le�w���/�B�Ob����Cm�k�l��*�����_���^I�5:Td"�rn<�� ��4���t�9����x:���˗/��>�����.�S��#�]�t	��EF}J-Q~|׳��"�ƹ��Yg�a0N�gL`>| n�!"�����UF�o?q'5ҘJmU>GnE^5�6L��]��[wQ��h7�$ݚ�Ve����ǅh�M�&�mV	��L��I�r�jﲕsTҕ<$��uؒK��ޓ}t^ך��J��n������{#���x�:����k�ȑTu�*��O/".g-��Z�j�{Jqe����B@�O�qAnT��Ss]����I��J1b�@��ϥ]�MqfZJ��9�9���83�	���|I��������ʧ��vw�����y��H�ϧ�\�]�iHc,��]��q��=#%�'�(n�=P�)z�K��OC!��WM��~a.$�H\;�H�/�� P�P�{���w �B�/<|���a�n���g�q�P�������x�?�}��J]�}*-�(�h��)�xBj!})�����ﶟx@�}� ��J��i�5�Iu�s&��?N�؎�/�W_}ɍGm�O��[�Ic��ׯ^����|��W���k?�'����e�eR�ٽ)��Cm���u�����.��To�
�"��}ˬ9*!�dX�)o���W��h#��*�u�ϑ���u�)�
ׅRS9���6��=�܂��Ҥ���5�6+�;D�3|�8�I4I]W��ikT'z���*����=Ww�p1�"�h��N|��a\4����reL��Ue��1Ғ�hkH�&�8�R5�s=��wt	2�1��q�}[x_}�u�*44�]M��\�����	��a����m���ꟺu�5��}p��r�նa���C��-�=7!�N�����Q���W0�w��ײ�a'��3$u��}���<�Ż$�l|+�]e�]�s�J�xw"[c���-j�c����]�ɪ�H栖���7L�`��~m�%�hxP���R$������?��C�����c��-==�5�ȗ/��Y���_��	�����m�|�'�bl��#[P�t(�`���`����7R��q c�E�~�X�~���������ͷ�n�T�i:�p��хa�G*����J?vP��4髰�f����p�g�`�Aa�h�Ib��ZZ�����s���������*����[��Z�����X#�t)�|�� ��ƅ�~sA 0t�h��Q����Ɯ�!��z(gY����8��:�NnEa9�*�x�EC3h�p��%��hXG촓�헵�R������#m���H[�SM�T��{wz�UQ`1�*
�`vO;e��mqCe�� � `r9eE�I�fX>���x|�a��w���x
��'�0hC���=�B1��){0�t��D!/����}/��mzk���lP��z���0����ؼ�W�!�a��AV_|>\e�aX�㐋J��$"���P4�ڟ�_�
��T
۴�&C1gn����Eu[ASwA���W�%;��q�Yg�U�f�Wqp�0�	,�F=��p�].�|��a�JDI�A�e'գ'
Z��1�	hi��st���z�"��q���2��P]�z���/ʷ�~S�zyY�R8��!g; k��^��"�b�c\;�lF��J6� �^�ܡʧ'�GIk/Q=��a��%�X~�1�ΐ<.�p�D�o?F�]p��e>�������f0��8fՒ�E\�[����m�ђ�K�:�5�Gf;�jw|?}���u�ϕl^$��NU��5����{���o����gF�?��!5-��T��>}\k���'D]�>)9�l�IG��-<p(����`���؀���*�<+�f�&�s�$���"�%�{R�N�FJ�m$�/7�Em�2�<�ȅ�V�ۂ�f��R�}���nO��x��ó*z7�b�R�����&=;z�x�p��������O>D���`?ܑ�l��4(������|LӋ���-n�
�p��%ۊ`�[?�i�����kq�OO�Hor�s,/mB��۞�|�Uy�
$�G�d<�	�A����z����67����KW��'�~~������'�#�u��e��'�b���;#Q�B(*�Ǖ�f�N=�����:-����c>��~��.��rŘ��>qP�6C4X�T�ڌ>��iN��⋢���������#�051H�J/wc��F�R���)o�'5F���>e�ɂ�(C5G����n�����[���
L��ҳ���]U��r��m���3v���i2����j��1:
Ko��\��V�k�1fw۠?��k议�?39թ�s���0��_�!OfǢO^��f���=	+Y\_;��B���ә�"�G������I�V(qCC8�S���5����6��L�w(�c�L��=qx	u�L��C�x=�������y��-%���O`x�����C�F������X�\�0���$O6��leN"���L��Q�Sxg8�C0�;9!u	��j90�`C�s��5�]%��m1��!D~��{��ڋ��.��g4��5�	�Ib^�����_���mPU&f���n�b"������������s��"e�5[ ��a��`����.��g�ox��ާ�u1#Fg�7�4U��H��>S��D��,���5ƾ����oޕ��OYb���7���1_���R_���б��3�'��w���-��_��8�L@)�d��ԏ��ʓd���EG�Btao��񖒆k���98<n��0�����#����b�W��z�:4�<4���������0�CCO�xf�""`�L�~N���ձ�r[�;�F�RѠ�����,bM|�����<R���?�[&|����3܃�6�JH'�UN� ��0_��摾(?��3�?��s`Kj*G�8��Sd�JcDC`7jr�km~��a�����E��n����%��6���L��[G ���/�Bd(��<Y$#�PN����=�`�x���J~D�v�cC��Ʃ/�
?��MP�W���N	�ɚ�2�$��3�����c���������n߉q���#��?��C��+(�+wm=�U�q�g��v���[����曯�����{;l���T�6f�8��"��z�ۘ���w�����ۡ�[��`���o���-�Ex���w����c�jlH����]]���5|+A�w6����&��X��`H�G
CzwI�1������5�g��Q!�-��������ٯ��e�|�T��<�`������ �?��Ss���a����T5X%������P���j�^�8<r?z\��]C�N�xb�=~z"�	�] ��tD?3��՞j���􎸌A��>��I��8�]�$��I3?�� OQKBb�lo)��R��*�Mll^�+�6��+m-�X��TX��K�k<���Ҿ!5ϲ>�u"��X�lU�.�CK�8W�{�h���M��;���������O����Y�iW�I�QXNp������������[.ns���a�J,d�7���81<�!`b��йD�B��RxxJ [�%\33���cL���SP�;����=�܅��L/Ix~��İ����n!���=���RO+`�7I�Q��MO�x�3a� �j���T�_m�A�T�N!}&Y�B&�#�x����������eL!�|�������W�y;�9�=�m�$�o�v�)�2�s�D<<�c񓚧��J��m^8�>�dl^��*����l%8�4:����Ŀ�#����q�$�3mX��3���k�,��?(��蕱�r�V��ϫ��I*eE��F��I��%.
��:%����Ն�ɶF�U`څ.q
��c8-s�0�����G���!Q�ͣ+jS\"��=�>�a��}͸��ۯ����liS��_X��W�xCB�;X?�����CgfhCz
Bl	�ƈ}s�!~�7�E"U��l[Acל�|؅Qjq�.��tڻ�1�nCߧ0�]�J)3DH_�R1� ���&{)E���*p=dT�$���"�vOh��O���'��(N���&b��fdDeP`x��Hw��Ϸ���u�'��t�=��q�����?H(e�K�<��~��M�0������g�7Y.�y��p{;0���`P�w�L&�#���f�%\l�%a����~*����f�ߒ��7���J���ű�(�I.�뱹�Y��"R�sJ��f3�KV�� ]��������)�m�١w�ד�}6�;�B���!r��pTDL���!Ն��^x�(��ݷ�rnp����?	�`>�lp3��5- 3�ASO,������N4�ǧh�3$s	�~���yO�$.%�2�O�<3����(����qfS+\�Gy��Q�{�����X��y홧=D;pU/^2��Dqe�V5�s���}'����[v����:����ꚗm*C�Gԧ�w���Q���/�?O�s�j�^֔wC��P�ޱ�o	��
X�ǃ���Co��BZR�Kʈ����ݲ���+2-H텅=���^R+S,+W"ܳ!�6��@���8���/��ɐ�l���Ķ��&���0X����Ɗ�[^��D)x�Ґ�F�a�fD]���Fx������1Ï���矣��nbsQM��w�&���維�ٷ��[mҳ��慝�O�)�c�~C�=�.�l�8�0����e�;�Q�7
oM<�[Q*�/jA���j�����S7���:�&��"Arz��`�����<�o"���p"�]m�a�����]%[ԓ]�(zW�3q�/7C��������s���'��lb��t��1�p�w���Ɯ�E�Ѷ�t����t�жȁZ����=�2Bez��n��	��K8$�N?��N�� I�zH�Ť�SP�B#A��6jj* �?+j`��,�,T�ȑ"��<P\��H�uW�b��|�.%�ҹ�=��ӧ9����xCȇW�b����M�\��#���s#*�o=�L35o��Mڪ����P�«p%S����v�&s
�ݴ*W$���F�5�����LцbYݭ4����U���E��y�Hr�C�ñ�:d��gy
j�2h�v۾���9��C(�/)ʂE�:�{�yz��D��4�k�*�w�� *H�jt����Q�y�������JZn�Њ�����8��WW)c+��I���cS����ƌL9���N	���W5�T�!���~N^������R���U��eZ����	��E0�h'�V/�������1Ϣq����7�D�uM]\+��Ç]�B؁��g4�싵����x�9���ڄ��L�������'�Q�ծjO;&QJ)�g��5��e���\�}{�4E]QYEX�Ɓ�����������(J���58,�]���l�:F!�iU�RJ\�Tқ2�-a�z������ΠC�r�+�sm����"kae�` �B��|iJ����n�p�M�}-�S��Q��l�5��pMFNk`�L!���=s�]I%�]Ы�.p����ث�Q�I��c$~W׽�Њy�0�}����7Uo�s.J�kE�ffp4�.z�8��d��wݛ>#�0��A���Ccdq�1Ĳ�!�R��K�^��*����f`��_�R����+b`��CӘ�{�=WrO�!��k���ay�L��,�Q)��������XC	�Cc�X�����_���G����`(��bN��<��g�u��¸�;zL��M�;6�8�wi@��f���Y_t̶��,����!6�ˏ�u�]��aX�	Ǟ{|RKo[0��pI'�N���[>�e�Ȥ׭_�3��pm���{]*������1Λ!c����l��M�>�6,tԻz+.��=���+�^y��zi9�u�}���Gg�)<��ôL���,���"ؚ���K���ܘ�����[�NY�p�/SXp]A߻��:rJ�?R�@�$n3��!d���A����X�Ŋ�0\��h'�ܜ�bϸf����sY�΢�x�D"4�j�_��{k#�V����ӦRS3
Ta��]P�`�0>���n����9����7'�*���G)2�!Kq�������H�� ��u���Ƣ������ߕ��C��_���B�ɐ���Q2ȇ|.|������������x�ΙG��9����5���D��W'LM��plHa��>����f������=	���!u��������w齐�vW%ۖX����%�Yb�P�Sԋ�PF�)hi��0BC��\_���vL$a�2��pv�"��u����=�ۛbؿ����m��`�@y?yo*�>�%"�Y���v#�]����
�i��6v�z���4ϭuj"L���Vf�`��J�ĥ��=�v�}�8g��j62�S��叠��oՈ�����?��e�9g�-a��	�����V&�'�v�Ľ8|J�t����D3���x���ǣ���a�%,�)q,��y3$�~���ڕM��� *�{I��)�����IKe�����N�i��0b��}O��v����,�g��..��a��2����1�x��/�>���mM�2�������z����1$��������葂�
����Sļ���bx� ��X�3��?mzR1�xP���)p�����j�"��t*|<K���<�&��ȚF�&��6cx]lo\��$���
�witi_!���HK�Zd&�]��6�i����9Go$W�����鲂�R�(�{�.n{�Q��zy����a.B�,�kۉ#����7^�^*]XQ��dr	��1��
�?#�y�qpT�׸��;�o8HSO8���v�I����k�(�:�����J��D���6�����g��`S��B>*1���K�d,mD9�}Md$�� �x��Z*N�������y	�>����(O����\��D��ءfq�1�JWZ�i�k���B%���$?D�^���,a�Ƕ�Ϟ��.�崮)��l3C�X�.�3~U�/Y���^���nv�R2�=�%��B��k�&���z�6��H���DԻ��-�uFs�l�׭$�j�Q�OCu��t�f56i��>��u`��d����k�ؠ�5>>�>���>V�6���[z�dE!A
���:ĤIqR���`�j���q�y��1�-Aj��%��V%�ΧS:UKbI'�/�y}oQ��j��b�BPs�C�d�h��P�&��W[�j%�`����_�f�s>K�كdn8�*#6��O���(��h�G{�X�.-U[�c0'�
2{�
>$�dSqw��b�|η��oG�Հ�����m>��o�Zsl֮v���$Y�<�]3	��:P� k�����3pa����˸���Ioyf}-�Y}ډx�E�er������\b��x���6Bć����X`Y����5��Z@�%�_���C�{H��dR+�,R_8�)6������<�Xý�!/"\OlVx0x��@�z��%��,��m��#�Q�!\��E�G���AI3OTf�����,��ō5@,��o0ڡ1�2�cx�k�^>03��F�s���R.��>��P,�톘]���Y]*�*e�FI'�� ����~�	�60O�;�|=��}$Pv����Œ�u��6B��Ma������p�z(Zs�X=���L��v0~���9�,<��Z��ԥ#����9<Y]C�
YW?Tn5Ǧ[��H�ܒ�!`*s3d$���5�ԙ��@v�`���fdk]�ӕ��y���}�mDM��=�zTt؍�/1�Hp�<u"Cf�,E�WlQ?3�����a۞�����6"���I}Hb�ru�t�i�1L�\�&�7���|��^}�6b��������N\��t 9�I3��v��9�d���#v�'�M3��I�>�{��5|NW��Ӗ}���z�!��I!����J��5��?���p���d��]�����!�)-Q�e��b� a������7����k
i� ⾔9�D�(�Nﶟ�e�XJ�t��� x/���oh���ص�/c���Ӏv��	C,k�4r7���{6���c�B���������)EHv�Α�]Y��q��f��07��m
d@�نC��.��X�׫4^����`��L��է�Lq���	�l���o���?����,g�3��1�E���wsť��]�1����cO9B�#~��~������� ��ʩ��%��o#�~܅�VeY�ç��+�a]"�dxNFTv}$���������w�`Y7��^�`^&�ߪi�}��~����G�?vnߨ�U��76��1Ro2sX��Fy���␥+]/�B�L���h�)4cS�}:�uF���ym��$����P�]�Fn}�2!�&���L���R�y�0��L���c�FscuR�b��IP���J����gE��q��;��%�Dɩv�� �������|����xU<pS����j�9Ƶ��I�)�/|P����F��&ۊɈ�ϡ6!��ÛS�(f2@]&%Z����9��:����<vg����c��.��I�wƗ�)�����I�"K�cJ��w�>9����[� v�|P˔+�K��0�_�\�7�|C���1�:;N�.��[@�0W��C:?I��E���J���.X	C����]�&]{war��'6<G䱬��>;�|9g$�Xi�s0`N��R5��՚|V�N��K�;�B����[����ϵ��b#���=Ғאa}pK��#���=�e6
��ye�&�r�|��	/8���=�.���'yFE��YmL��%�R��q�{���{�+D���4�/��P+IL�Q���:i$V�`�eeR��$���=�4�ۢaF��Kb���j��Z����l��q�ws��J�<lR�s�I揽���,��5���$<��Ÿ~���̼J9��w^%�G���3^��#�ܢ$��9I��5�q�P0���xd���jD��ܮ��F��2.4� �5�4�݇��^�!:#A�g�h%��:E��[%a��a"��RJW�<�CKB�0�qX8W�l�Y�����]&O�������S;vY)DJ0�/���	Z�Z��	Q�S1�a,�p;�nFiZaǰ��� ��o`y���� ��b�u�ys�WQY�)����
��qﲶ"��ۧ��m�"�K2|ҋ�h7�O&���J�duD5cY�xxo�Sx���ж��g	��2��hKK���w��]�x���$�*y����(C�ΚcV��Iƨ<��F���@�V�.���J�+����~�"g�B#��DI�1�������Ğ0/�y�sH!|LRxv2��I9y��X(��z��\���?Gi$ƚ��,�������G��?��+iX�ٞ�q�h�gx:��K�߷\�
�V`8\��@u���0�~F��%v���(��ږ;�@�탄�ק5C���+�9Q�q�8��+�}�֐�8Vr}���m.��?�rI�v���5<�6�y�lOT3}� ��Ƈ�m���A���^�!�:�r��2�Q����3R��F:�4�'�'��Ȑ>�z�u�Q�N��Z	d��%��Ү��SY(=�&����9�l8Cl��Vg�X[�I���>ց���ݫl%�a�̒���X��^|���zZ����N�,c؁r�����#+�6�Jnm���kK���}nN���о�@;��p���sT��iO�ւ=yNn�R���x�҄^��>_��(��� ���gumo�6�!5�1�@q�N�d�C�85J��Tr��~Hc
� �G�>�ZҐR�g0���p��s��")"�_R��=�³���a\������4��t2Ieq�t���ު���_}�q�1�UE�1�����=�'��Ht8�>E).���'T`�8@���J�z;�!������,1�0��@.p��-K�WLf	�y|����t~9�Z~��M��]�����c���[��B\D�K��6�n	`��/�܅�Yĸn���0�<saA3Ú'v=�G��u
����]��*����SV�����֩�{���p��˸���?��ch�v%�	��TU�X�k���Y�=�ġb���X��Ú�Q��sHoO��L���2N:��j%��}&�����I�]|�y��'���?{4��C���&w��s��鰎�sc�(� �`u�>J����U�ҥ������F�F|I'
�P�9D�)��_�,��޾5�.�d�uR�YW�z�X��k�%�������M܈(�,ۺ2�G��>��2¬�a]�G��2��&;fV�8|��\A�q8Qj�ݻ��~(���/��'����@U�%�������n�u�)Y����>�C	���oB�D8��eM�#n[f���1ď(=�^����7�-4O����JOV8��V����%�v�d���O�����K��E�7;u^8Ň��S�y�.��O�S$ N<h~�<�����xQo#uT���$��R�x�p}�:[�
���N�.�!�S,VY]{�����Y�#ˋ'	q�;ȁ���D��qX��柆���y�C�]xhd�@�_�*���c�҉��&I��)���Y9n��?~M�[KV��A�s��{�'������zϗ��լY�e��P�%��ژ%ıd�!���uŽ��9
/��TB%�u��v����8���=������g���df�G�y
{<'�BZ�վ{�aux��\�[t��9BQs�$v�1đ�ĉ��%��,j�:���QU}�^�U8�R3�����<�a^`�c`�a�y��g�hv,��RXt�g�7oB�|=�2-F�0��GS�7�v��/����Z�O�+f2Bq�)�Cp��M��a�=�B(�/��j�ܴ�׺P�Z���������	E�j����c�ш��o�oyM���&�l^�/0 ��,=���W�����c@u��`!��"��͟���)Y0��`;$=�Ɓ�5
��i[C�%b��6f0�0D?��Oz�7��T����kU��~d(���k�&OT�S�6� � ե�c�ŶWXauCz�gI���׉93-l<�2����3�x�k�p
�ou׻<zU��uȮ�̶/�Z��0�1�X3��¿�r�R�O]�(%�Q�G�ޟ��b���$~���0T�tP�A��wGm;���w���SG.��ƹd�j+y�\Zz�v�?��?�a^�Ol�=��5��
黰D�eRykDI����M��.�H�>j�w� �z��a3�E���=Hb�0Vؤ΄2D?�i��%h�22���x�s����$x��d({||�x���]~7�3Y�I#����������t<,f\76�K.�ĵ���*���3	^��e���������R�5�`��Q��~~�p�}o ���8�0����C&=�{e͟�>�B��X�#���a.%�b�#�YǇm�u0l�ǵ� ���e�M�ۻ@a�w̃����-�As'�������'	Ct�,:�v�w������/��F��O���w��Z�!�Ѣ!���k0��!uj�Z�R�vM��z�pw{a��I�b+�����~;���P������'e��i��V�F�6�=�|��7X�R�'�qs#ąn�.�6�8�q�1��MA��E-Ä\k�O�T�7k|�Kէ��NF�KC���j;{N�Nc�!;��c�UEߪ셅1����,��,�Mc���?2��G���2<���#-W�K<ؑs�Oe���(�*)�+�	� ��'g4��E��J�5/L#���c�{���E�"s3Ǧ��']E5Q%3�}�,->��lT�Q�Ix�O�'nc�Τ�5����f(�o���#S�'F�*��JX���$)�
���^���X�6�����
��}I0[��9��=�v
���Z��2F�Q�6ju����P��-�N�oW����{�-�A�c �O�t�S��=$p��t%�$܂���?L�F��݆�4mJxaJP��v˰�I�0DNRY��M�{�:��6Ը�K� ���ǀ�`DѠQ��.��U9aI�飸���@^��HԍplB�#G�LCr�k� 4�@9j{=e+�@�b�+M�oE�X�4��T�+��ō���*Th��}��Q��2}�X+�*:�)�mDI��P�%�_�F;ӱ���}�K��P�7{�J[UK9����`��y	' ��������������3um�����Cõ����e�L��{�K%k��%^m%�q.c,
��{�%iH���4��s�]�P~~j����l�R �FV=��  �����;�2�v�w^�1�	��租~REKp34}�g�!��)��c��!0����i���=�C����U[���x��\5�@�Z>G����ڿIc֙�Q��Cȓ��K̽�9�m��D7�!�(��g6[�B��$�l��WBD����e2��_T�b����>hX�f�អ����#�q�xF"3n�{����Z`�7��<�]庁�] /�~�R�����?D�s����D�H�d)97�<�@��v�.��*���ό�p8���OC�l碄g��F�����B�YPK�y�Y������k��Q&��lBMz��!��8]�mX�|�����d��CeCIOѢ�L�"��,
믩sm��V%�l�!ʥx��On�'-ђ�5�l��0��V�ħ
�E��Z�[4�.�?�ssFN��6���t���հ7�8�į��}Z0V�J-p����>���gM���$�O曣`AY2`�
a+�\CK�Ǡ�z���Ln�0�
�?e���/qx\�,��s���-�)<§�6�;&�Jf��!�Ӑv�Aݲ�?�ޏl���S�>FI)QR��>�z���������t}���}|b)���
W�t�WB��:�0,s�w�5�6�3�.I�_���J^��y��n���$0�,�UA�O^�"����7�}���N!��"�i9�p�irI�|EO��0��d���a�GK-"3G����� ���v:�M	9G�O_�B�#�o/s҇�pq��4W"��zL��Ԯ1s&�������&3�Dy��G%5D�+��*����Z!5���(&��ó�I��Z���;�0'�fO¸�q��A��w?�[U<��pV�T�#��'�L�j��¯�
Lcz(�ɉ�� �:���$Dr��Ё��3V�sa�����%��T������@/�fy��c��ܰ5�x���r
5�'��St�<� �t^t�||b���<���X������䰆 ����1Z�I\wɝAu#JH�܌��44"Ӭ��!�����w��γ{�wN���!��=�w	��a�tHKu�8�NO���9���E�e� d����cp;�[7�&.ġ'�AU��7�A~�"�yZҘ�!�ü:zN��C�8�]���X���;$�v��8с�?�݇S��kܟ�	�7�I���P�f�����(��((0>�a�k�k�]�����1qыү(S�F��{hNUz��C��X7����qb�1��9�^K��[5������3����#�-�m�X�s}^+
��qm�mT}�Hd֎u=\x�R�Suc�
�q1VV�k"�V"��g��ז�?��9ѩ0���d����7,.Nf�T��
����h,��^I�>H{��^�٫'٪8y�g����Y�
I'�l�:�u��<�x�pY�3�Q�?k� ��6'��7F\�L�Y^({�r�v�>nV�t�3#���
��VŦ	�*��ƅ��*YfW�0q��{d�
4u���F���TK	sE������tʺh%��c,%��t����fh>���}5�����üϾ��-�rp�}�n!4�z��LkV.ל�%
G��u��za�<:c�8�%��5�������9���r<"A��l։�b����s+J[M	�t�+iT��m2�\y�}-:!�3�,K4��C�i,$d���eaO�1�	��!�Z�U�"����x?�	�g�q��1��.f���]����H3@��k�p����L�I�J�W2�gz��t�
�퍖���&�Jz��^����O.�BHm�{h�#U(`umf��t����.��,1^4SS��!��c>[2�����H�X�Ș��Ϋ��W���=��*�ӻxۭJ�<����D`a��=S�ݵ2��6Y�m��a��J��ҷ����R�Qj��ł��VVhD�A�+Iկ1��e��.�l�I2���K���x}�v�{��k^Y�m>\�#�C)��<	F�F���Bn�1c�,�N���E+�I�$�W��Uo�#f��$��w�'~D���I�:��^��E�H"��E-?���{�z�H;�mN��z��[�Dey�fP����t��1i<��x��k/�9��G /�e���n��,p�==Ȼ�o��k�j����cDe��jRY��Կ��_�p��
	1�\R<�<�W98���i��ڝ�n��̕\.�	���M��;镆�6�Ø)�tLQhu���ɦ���1�W�����[������4�!CƓ�	�����,j�a�A]zs�4��@[��E�B�����F@<m�l^hP��xd?�W�j�ҫt��}�j޵p�|j'}�0�A�Ϙ�y�0_��������=�uۃ�x�6�'��sx����ī��`����4���� tPȃR�i��YJ-�5m�_;qE��$���ڠ�^'��{X�7kt@�I��S���8�2�E�CO#�J�ٙfv�l�1���0�sxS]gOt��mm�3{��DSf���>�u�GY㲖L\�hԎ< Q��ǒڦ>��BU�a���cw ���qx<��C&�����F>"�%�����0�����>4��0�i���������h�=6�]�t&Q�(%�p4�z�w\�r�g�������H�u"��OAӺ/��}��<����`�T���`B����G���In4�F-ib�����S@H�
r$j�ЙB��1��6�^+�e��a���ц�1�W?���1�DYf�׶�=�к.�P��L$�c_d��;t2��<�����v�-����q������x΁u�"a`�K<t]�{���]����*��G74^P�[5-�d�*L�ז�;Wq1�圸�At�~U�	���BBor���m:���'��K�dH�Q�xv},�9k��Q�v���+�X���UX��6`_��H����7w�=灰DM�#�W�j�!��ջ��?
^�3�c�z�oc�����j��3æ��u����c�]�K�{S��,��ac�J^�0V�
�hbUVR7��X/N
9����Q�h�w��aw�CF�g��ֺs�-��O��iI��Y�͹g�Ɋ���t�@�-}�+���j�� �A����lX����5R�s����]&��HVK��i<�{z����!��#i������ 7�x�cj��� ���2!0SU�P��3,_hXݳ��*:���Z;?0�"Xa
�B�g�nYq��mei�P4���Aa2 �M��pE�*V���>C�0�d�슉C��u���1&�ba�j��=��tE�a�� �{.V3�Tl��L�nk%d|#��Ơ�^%��r�L�Hx"Ad愠��2���q�=�4��E�0V�n�׸"1#]��e��`o�5mp&j��m@i֜�cH�Z�yQƾ�Nڹ;CP�lԆ���t��o8+���֐�)�D���'*V�(�Duޅ#R�+��:s�>6:�}��Jvy���<�[c{L�6K�{w"���`��z�}zo��?�ۭ��5t&� �]���^R�RG�����3���N�.�>����*Ʉx�!!�>Q� �"��|���Ԭ��ظx��4�G��&z�~gL���'�%5{op�UM�N��uZ�6q>���9���`��W��]���u�R���<������rKj{���B)�(���Զ$�7�g�&���.�_O&�?X^S���9#Q�}���Zoץ����QJz�]��2�5Y`~.=>�	$Ew�D�����cH?W�cSH����r�yS�U�C��d�Gh|c�<QWr!�B�+
8�X�
���)����ީ�t�]�;������2^�����W�^r�]� �ld����R>�m��n��v��������Km-�sqCps��YK�Hm^��1�وWY����:��~8}��?,�p�vS9d1K#����e��q�^����BK�6����DG�&<��MAK|1BjT�Z��k�.Y�VnK;z�8��;���*���r>?~ʜ�x��=�NQ�r��Z�)n�)�L���Y:`��y���`�3�h���s�uu�W@�ځ+K���2�lL��v��:So\��5�t�ך5�i[y�Gzݣ�m��ӹ?��`9���F�E?��8��3���z01Ԥ�Jh[��ۆ�N��A��I咧���%0$	���ԗ�{	�����~CR.�r�U��jYZ4�pc�l�8-a���l�ݺ$�d�6��$�ӑ�l/O��	�W�;�\/_��^Ay���%,��
!Ђ1�f�|WW�&{���K$È��c�*Ԧ| ��i�*c{�bo(<&Z�����v��n�`�LCY*=jH:��U�>O�I�3�p �������k��Y��mwA�P�m���;\��CrNbC�֐�}3�QaS���5 %W��h���@�����$v�Cqa�UU\�gnťH��=��z�"������41�,��	��@6マ�t!�к��À��}B�7��|(g�TӇ�Pey����bB�^�~�_?#�-�l���s�����<�!����U	!����
I�W����2r�w#W�V��z]�
��_���~ICtg�����7�E(L��wo��l�hlk���O%��$����C�}r��_LEA�U��C�D���\b�ج��d�o������~��O� �!#���V�I�X��k��C��"�\*���?�Vx3+��Okx�%�4��9�� �PP����f���Ik[d��}~^�d֎F��]&~���A���R8���t���f��q�<x��Yyq'��T�^�k�����=��8�a O5�M����q[g7�����]_�2Cޅ�R�{��x]��m:
h�|'y��.��e��|�����C��P�1v|��%�f��^�SߥPP��&��b�쬄���v[���*��#�:�7g�4)26C�nkf������{ᰬM	ys�`ɠ#�:���v�J�Qc?��\�m�v�f���d*�Ms��7�����z�������_;$��P�l K]�f T�M{V9�)�D�}�d4hG��w��~����̶���Px����Ր�Cu`�����ET!1��Nl�n���#.x_8 �O��m~�fL��l�S��?�")y�k.(q��������5=������m���qϐ�`?��%k�UB�*
U�&����$��D<_��4eB}_Ss�Ԇ'єzZ��8�D;hh�kdPZv��nܚ���(��M��$��ɭ��8����!	'CZf�Z�4%\���=Q����p4eK��� JOOe�~7$������u�[YE��{�<nƒun�3� x6+��C��@���9��9&�n�!`H���iL(/m�tڜx�����s����Oi��v36Z��bW���޾|��Wعs�30*�
���ژ�� %���A�"=i$[��-��YF(|`�>>\��,��׫�}����}��c�t�����\�X?=sVۖ�w�B��"؍V�
|��!��S���1��N��d����ڤ�����vaC����jn�Qx�_s�kF�3;��?�2�5��Ꭵ�#�w��Șdy�~F���q�33p��L�Ȣ	.��&oF~'.;v>'N�v��4U,L�6DdG7�ӓ�'w�C`�ڗ�RЧ��䅒-kV�H�t����	����¢϶a6�2�5Hֵ���cc�Xx,w�X��C�����l�q�<7o�yP�.i4�`��rF���y���kQ����M����(�mM��(WE���/K�Q�G*Y��f�|c� 4�۾�6<����C�6��q�7��-8h�߾����Ǉ{�ԕ}v[^�|V�������QZ���G�����0��ț��'��ֆ�V���ё��*5�����/�S���Ǐh�������O۵QUڲ#�͈�#�Ð���<R55���Q���,�r���L�h�]��<��=�$��n׾���N���{�<ExCx���i�!�CLC�dֺy�=U������$I�b�̌.]��y���,�C�G�I؎�S����W�%U�P�]I-Vm���[Ѯ��>������Ë"�wI�0r��7McM����?0��V�������V�z�7\�_�4�WV��]��O�
h�2AG1�ݒ����%��H��ϖ�Rkla��/�
=X>�޾s�V��x�x�떍�bJu�,;}�:�%��Lc)�����$�E���LZ��XI����jf��'vt!]_������3a?�p���c=� .v �ɫ��B�W"��s���]�����:��8�Y��$J��YR���$������w�p��!�1Re�W6��w&/w�o�B��8?�_�ܞ���_ыe�9��`gHV��w��Q��ܨQ��P�T�gw���YTm�b�^j����	KE�.BZ���3,URt.�%7����[9�g���@��ah}�񐸭�z�����:R��k-� k�(�=q�����L����~:J�H	cS"��1��1C�����Ո6��]��\������Ⴞ2I�H��!�x�VE�����#���m���ui�j�s���g���x�`���Da`�����t�K�l����ߘ_U58���	�xZ��)]d���47�1g�d`;mߠ=M�ū|;�ָJ�k�ey���ܯ��`��KL��jt���t*��Z��"�Դ��<~�V�08x#G�?��f۠��a�������~��W�s��j1[{Y�N]a�@��M��:��Vf�a�u*�|̆m-��MRrQx��9�P��vy� ��Ð���w+<�5�,����y�.tZ����)��<��� �m�σ��%?|(�͈�e�u_�e����>1�_l�ź���u�a�
l����K��fK
�������B����ݭ:hx��>��P��a�ޖ}�)�w
��]�V�NC��0ڨ�W���~Z�zD��.��<EDW\�;�7D���!y����d�j.	��Q,`�1�B��m��F�՘&�����ϠV��ަ�>��{���=�b��0p|a�1	��y�V���ۡ8ӋUe�%D���������?K��v��/��jd���Gʯ���7�+�����C���\����wR4�Y�*0`W��Bw#e}u�����x�I�I��FU�ifЇ��/���c�0���|�&v�<���"c#|��������<�c3���2�m��:A�2��m.��+.�'��*���y�MN�B޳�MtX|b��������D���+gI�A�����VϥU�u�P����D���I�q�D�VY_N:��gx�bF�K���NzK���fr��Y����!�pϐ��a۸_~�U����JzT�8*�|�����^����>]���=����<��N!���,_m��:�xBQ��9:��$.�#ؐ�`�H�h���z�����q%�lxN�� x���ޤǆ�o���=�S�e;����,}4�� �������?�R�V��Z%�[o���n?6%.��:�)�HoRe��h%��k�B��*C*�^�=%����g)T��w`�@��ի�������.#پ7�`��]���~f[�Q_��V����Q�?1��Ɔ�CZ7���:�� �[��5�ChNeJ�B�H-]e>�Z���1�B�m���u� �q�Z���	��ZE(��>��,Թ��Y5�k@2�0nh6�������n`Ha�ݠ�3��P���o�����v��!�َ��<�1�'I#��`����>H�Jmƥ����(�%��p��υ��C�2�9��`��6ـ*"� �j,�n⾸��J����.�zI��ң-�Llv��/�������2��#���*���5������s����_��C���������
����q�L��_��(S��,�:�����=ҋ�}�/^��������?ŵ�܊���ٳ8�#2��ݻ$޳|v�^Ԙ���[���a��1e",(D��*�ּz��?co��q$FfV�t7I��fg����}����I"�7�:��473�(��TT	h�P������9>{���~��r@�Tΰ�'��]��웈�:^�7���B�����;P߰��3�!am���K���f�l������{�߃�̲ҧ��ǈ��s�+ƞ1�#
V�{���Y�a6�{GG��,}�% �(P��,��q8�߳��7z��^�w�ڻ�[]�)��(���s����E����۝��]bb�]V'E���\�6��#T�i��Is"1w������+R��H�+���a��Q�O�H����O?�(�����}_;�fF����L�Er5��]�/�F9���g�_�V�4��g��=9ApaGE\׷�����%�����d�`ɋ+��6�K#%�=�ɕ��%�uH�f,l�s1��l�;W�md[؋C�m̑Y��Z��4�_�� �?����K�2�!�|������0�2��gR�>F+�V�������D��zۈx?x�NJa��i��b$�������p��?|����횎L��'���=� ���5)~�e3�WC�Y������5�+�5X	�Ԏ�U���׮���U�9G�l@ a(�Ȏ-�٪�Q]a�c�0��Ӷ���#7��^�`�QQ�5��	���j�b>�(�"0勞lh���V�p$�K�} �X��!s�]iݎ9���ꝲ�ik+��N�����/��4�i2'-�u�摶ofC갳��2����YVd�#�pu]�ϔ�h����>�g������B2�ť_�P���$���4��6�:�`�1!*����@4GL�8�R$K��NȾ�0`�K��X#�:.�G($A0<�sdP?�
>�X����
p7E�t:����D�c�c
_���:P�����I,by�)}7L7�׬F�v�8N'yħT���}Q����t7�AQ�t��ԣ�I��J�ge��MNm��P	���
�? y�M��s��>G8��CM?	���əY��К,����߻�xL)��M�y�h�)��! D�^��.ƚj�L6�JyT��!�^#�ެ;��=b�~1ָW<L�k5f�ی�]py/gbӅ����]�Y��(�1����%�(�0�C���W/q��o�8�4��+[���#�_�@���NIOt�s*����Ÿ�ÁѨ�MCr�t����:E�S8n7����4���~e�~I{�e����W�}{��J[�wԟ���y1xm�"%��e�q&�0`��j3�]sq>9jQWL9�ލ:�X@��)��V!���>2����2aR�#}���������O����y+�X���i[�0���q���+,J��Y���ҕ5Ðv!x{��S|>��+gb1��2xćX008�a�z0v�ې�c�E#��H�����';�fѱ�!��G�I7��o�zN��2DU���,o������R�Q��Y_�"�))U�v��'�������x�?��>Z��!\fa�'�M��#x�3�=��9���$��G�Y�������F港�R�$��Hw:l:U��H��=RWŽ���jZ������H.UڰK~����!�ǔr>֨��юǽ!������sQ�U�߈lP�W_��BΘ+F#�J���-�|?��z������sxPdUY&j�N]�C�{~PKq��w1v\K��1BĴ`F�E-�Tw/s(o�ƴ�m��u��qH�M�>q���:�L!E	�ǆN�o��l�j� ��.���]$. �gYL}PP����� x �D���tL�m��u�X�z���-ۥ'C���vǘ$`F�@�4!Ģ��!Dq��/q�D�Yv�Y^9*�]�l��q���y@�R�^�8��;����`���e��c�n}$+^^N�5�$/�v�~@�i/l�ka��p
	�$E��p���B�	�.��y_��*�p(j9ž�0�vo/�UyQ�x����M<ewem�*��Rw]V��a{`gؐ����1������e��nG����;uJ�w�	�b:�R�%���Fu����1i=6�*XG{E��kz����I���N�#�z
�C��&� s&+_�$��I.�+��b�`��I�Y4/�=-��7�h�AR~&�7��7J#�h���VBA�dS���4�NV��� u��޲��:�E�YM�$Hzg ����ImR��ldY����2*���"��dΪLԽd�1O�bü@'4Z#����7�,�7������:��&�K�}y��6�����Nde���D��܉q�(�9
��>/B�Yc;�-a�c���(�����[B��B�Hn��3k�q�/��-kme͖�l����]y�V�b���[�����g����d�/�����J���ڮg�a�>��E٥��P�R�[�O0,�|�@(ĭ��0�����Qq�&E*0ե��Z�c�J&����ފ�6��//'2ҋ���]���ʨ
G3�r��}�\�xUr�M�e�9Z�.�g��T���e`H�糄V��;#&8fXLn5��CVEb�M�7�j�J�"ӘY~$5��u��,(M�����0��o��o���£��`������-J<�mªr����x8$�g e]n����K�Wj����-xbJ�,}�ྑH���P�Β��=�N̒�.�g��Y��2_㞿4����'=;�kIX /���J�	Q�4�i�]�h����|Wa`I���S�"���>\��w�����@���M9�	u�˧U�����80K��D���hNG�H�w�����q���1�["L2���$V�q
�{z�*+1iD���~E.ݗ�����X,%w���I0�O�6��%��/��B.$UT���-%�`D����$P��f������%�~�XK��g?tpf���Fq���;���/c<.���.�R���#4�!f�M�6��������0>V=�5��c�wC�	�kQ���8�[m��ۑ���t2�
q��ؕ�_S"��wd�EP��4�pquT��<�s�]!����!�W��z�71�RZC ���*��k�j��(���|���t�)i=��x3��d����5GF�1�6��%8��~���p�z� >I�kʪ�h^:8���P�6���a��P��T�Ev&2��������n�ID��ꃼT�5�6�6��rIWu����Hm��kT'%���������׶�L�nMյ_��f�a�B���n�����X`/�7{����&'��G��%�媖�+%�T,g�Ӎ����n�k���֒H��H�t���CQQ3n�2�p�I��"Ga�,<�)��1<R&S��O���a����&p���/ݮ���FZ�}�	�؛�F%/�m♗�-���Ң2@4�Ʌ�7d@�jQ�6l;$%s���Hx��0���T��^��U"�ӵZ��� ��vip��y��
O�<�亳?�f��\�X��]�Gb���E!�0�b{��׷���"���4�b'g�We��]��:���6?�oh2���X�Y�{!c!Zq���4�M扞�������՗L6/sM*g(�ђz0�8���"�j���Zp�^)��(���Y��zN����	��I�[���*; 0�טA�S}~��לc��|�{�gOr5����k�R�GҚ���ԕ��5'���Y��=7�Q�T����rRVSt���v �wE`v%��9��,[mt�̠���F���AE��@�QTT%�(OnH!�S��,kz��ĭ&yaK-a����"h����U�E�L�����^C�|�����wa�������Xy+��"C�T�a��)k��9���}�� b�����)��q�{5ɢ3���ܜI�bxgv[	:��I���;	�����o~�5ᳱ��P¼�$N�Ćղ�7�~AȞ#�Ì?���|�F)����`I�{�|O�T���ͥ�.9
8���ciY�,u/��k��5��n����-��r����0�8��#�Xr�j�:��b�5Ǝs�&����9y�~RM�,�H�c�8��ry�{y#�fq�|[~�`�Ũˌ9����_#R����/�H�sV�,��6pǵb= �2�۽���� ��;сx*n����� cK臒��G%\�,4�k&�m�ر��7���T%[~�mb������lP�+�|�� ����J�㼈��b�h��]�OC��BL�
-n\�FZV�%Ɛe�ͩC<�a�CCaHA㘩�c"s�:?>H�O��P�.V)km���۝|WM@8䞍�5�j����odn��𧠺 �YCteR�]�Э�C�S"��#{�!u8�E���]����aXq�.5�[��4�]z��/w���s���1�$��րDv4<�;�2#���°�-���܌ij9�('}Ì��-��[����S�� C\1�-5P�lM����2�Ɖ� ��p���N<�z[,����Klb$�X�t
.��l�����`������:��u�K��rz��a���t� ����S���b���];p0CN'e��Kzڟ�B&�0�DV�&1��w�#0�H8a�`�p����)�ۏM)%M���g�*�=�����*�ދU��}�[��馤V�6�F�E�W� �7�m�#JC��!�6�<�i/�%�)��a��{�5�B&br�Ւ.-�����kc}�n��)�,��*�G�S���-���dp�3�P���Ъ�<��P���{3Y����"&�r=�a;�Cf0$a�M�cM�*�-�xH�4y�ܐɩ�^�{A��4l��a'�)l�����_���>�0��Ҟ!�}����<Ix���J���3Ԯt�G��s�jQ��u�T'ϐ�u�s���W��{���hM��5��7u�WI&�'{�q����;)4�-������0\�\
Q�� =�ș]#S_ˁ/�4�C�v<��,��M������p�G��\�kNTfg�N��(��(wz	x�����:L੝�"���E��8�	��#���?
��A�ͺ?�#���}�� �@� �5��4�>��A[{<�#)�h�6"*E�0�x����?EH�z������n��-��fd�u�����dl��Uv�+Φ��Y�{���Р���E��P���Эq�� ~���f�V����-ڮ���e��$���:�\��H��g}�a������I�1wT���(��|3#�V�(9����z+mm��=@bUL��17�[~��7n``	�U��.km�S���T\��&��T�=��޹K%�j9���~����JS�z���!�Uh{S�� ��\ƝD����I�Հ�4b+3��=�IS�E	?��h�b��o|NNo�Ezv7 ]F
��!��x��G�H��Ø�yIl�=vjoq˨� h=wT�a���Ab����~���M`^X@q�}�w�|*+�T��MlN��`��s*lB�37$��`S��&z kA^����G	����˜�x�T��iQS�H����JH&/�+EE�?Zh��;߈��v��,���o�w��>�O���)�?| ��|I�����w�s�<O5I���X��I$'sW�;6;�u����e��9�a ��=j�`�XD�kE�]���W9>-NZ�+��4i&� 2fX�ޅ�k5���Az��v��t�QhM�|<��;���}�^3�gq�!����Ƴ2��b�f�ݣ)W�� ���̧̒��paޔ��R�jl�������$=�Z���ͤ�MJX)�'�����'6(K/Q"������*����f  �WB�����З`8���9�ZO�?�han` �E�!Ø|���lw�m����~g:����˛����`1����QɵP%Z��1����#ta�g��*�{���b
D�&������C���P���<`�B�k
ܠ��Y���#w }����k�S2��A#���X5?�c����a(B���O���ew���"o�����#�����(�9��hk�o�&�+w;��Hu0��c/���k M>7*���������������Cw2�NSڮ�w
�i�Ae{�H+���UѮW7qH	���vm��I��&�ZZ����#v�kV�"�w ���|�yOyj��ΗKPW��#�1�W�ʐ
#5UTz�꯭N�V��B�4Z"s�DJ~x��z��Xn�aR��@%Pv(1�](�@n����O65SM��*6�T'���rN�r��
x�-ԉb��,N���\�
�9���\P��ק/Q�!�h!�D{wW�+6ڶ���������N�N�z��E�:V�X�vM��B�-<�K�
P�`n��S7��L�'��m�Yj�Ȩ$ͨ��I��0�0
n<X��C�����(�T:�/�z&��훸w$��w�OOa`�6����!�Q8�,1z>�~Kա܀:���G�c��j{S0H,Y�����Ps� J?~�nC������}�h\�蹗;2�K�dG5��,}�_m�ʐ�i��n�C�Q>z�>� 0<(��ケ�������������fB4�ߔ������h��D��]��*E\��ą���+pB�0+�ُ�V�yRe�޶��M/\�}����A5iͣ��8[o��&��=�Ѵ��x��k���~c���b�t_}C�:;�����j��	���$�"æ�̰z~��X��`�v4.���J�:���y�;v�a�i�/V�
�`��Hè��,b+�9��\5���v�P&:DZ���S\UxG�㟢~z����&���{z��=�lc�F�=�=�D4 `���?n!��X��9ل�yM�PI�6�SD䇁B(�(L�^Z/c6KH�X#d���Q�V�t4������䦦oJz�˚!�H�1��o��TB;��a��À8h�����g�(��M1�`:���L�������S�͔��#�dF��DYl�mgk���L�oL�{�#������r<�4'�"�1�m�ktx,�9��I���4 �b�6�LH]�#�ヮc;�q}(�E���	����X^�ϗ������������ט7JlBbW�#��.Tۆ�%t�v1���X>�s?Pkk�c���	�r���w_��i=��m��������ޒ^gM0�J�S;��ǵ���Ȗ���LAkMK�\������%b	^�H(����?�J�ۼ�������������!H�Wf�k	����H��]�t+q
����V)�O8�m�^���XlP䁌¢(!ݮT'��Zx�%qXj ད�L�v=����������˗����5�*����EaA��L�y�SOq��
7_�I�q(���E����lX��Sx��C���%�����:HB��L}���캤*M���6��۸-oi������_���?��Oq��!0�sA�	O�ġB�<�����_�k���a=Z:o����D��Uh]U��7:	��px`����ت{��l3z�6�{��p�ᷳ�0���Ѳ��Qz�>,���ӟ���kzbu�_��桥�W*ck1���3ߛ�a��p��QūX��y�|Yc��#��������)
�7�J���-��{���N��D3?�I;\~p<�w؇����^�P����I-��/���RigQ�AO8ztO�����ř�������=43�Oc]���>�����&#�ũlٻImj^F�Y�ɀ�u�� wmYS�:�E�$77Jwu��L����d��V���c$�2H�b��_�*][�>ܝT�z:��F��^��pJ��7���F�R�SfI)6QrX�JEull�*&�ӧ�[��a3����&�A}mhH�ğ*�j�X�����,LL=�b��d��@b�=
�õ^B-�`�O������5��j�=΃��df<�67Gxx�kcEۍe��1��PI���|�xT]�zg�8��z ~���aH!�����a���H��	��2;��ڸy݄�X�ġDCJX��3��{Jhڞ?�C�=PU!����;te6�+� �x^����9�Ž��4�he�׿�5�Ƹ_J��Q5�D-��Du��H���ʻfS3��44�9�ۯhF1"�h����y��Or^���bMR�Io��ivg�Y�s62�)DιO��ƹ�|/˗�w�7�.R��U}L�A�?��XF��PT©��^�z�a��f����F�	���۲�Δ�%�m6��E�ȩ�!<��Q��E��ܲi��ȉ$r�/1H�=�3�Ђ9���t��v�m��[PP�%8`�����mH��{��B�k�߮o%�vH�Td5�0ٞظ�$P��D��|mH��P��@�ݻ?���������O����#�*�4��	�)D�jJ�-��7�R,�����?'���~/C�-C�҇q��|x�1���X
�b��1��?΃�*ċa$�{<��J�9�B��n�dx���[��s-a�xl�58łb�#�X���D�&�3�p��u�=��_�e$�c��G,E-Gܶ�t9x�_`D�>�p����ݔ*�!+x�A��i$$f*���9`,����Fi��(�(�Q-�%�	����B����N�!�"Nl�G��u��Z�F������k�G������-.JF@�ݏ��ZK�=�*�\��:|S��e̤%bM�0��H�U���6���R|� ����k>,���<���e��T��g�8w���e�jn�:��<�ր6����u��_U�����K���d����E�j���z�'��ߌ����s��:y`)�ܳ#ט��J�g���N.�rw¤�
�CҔp��q�ԋ8���{��Dۀ^��B�t�Z������;���-���v{�k� Y�-ŵ������q�jX�@#J���/� ��pK���rg	y�kx2T!��-u�_�x���>�t9���.]��`��fYj����IB��O��;�z)���o��@���YcxyC �]352��{���u:%7�H�!��Ir|m�Y�����7�4v#���|�A�C`˘'7p����7SSg�K��O�t/R�Bb��������� �P�kj�D��b�/��\�v���*L�y��+���6���}��UHY��y� ��\A-�,���悮)�n�LJ/58*�a�Z)��
A�ߵ�����Y�ƈ���M�6I�(��IJYBo�����|=w�pg'S���Yi�O����K�Xq�8���˼ġ6P�>�{bb� ��^�	���`�L�v��w�қ�o����R��S��~��!��cp��l+�\4֏Qq���m����h���zZX ecӘ�����I�	8��0��5W��hA�m�',�%��������������I�0N�P����k�wެ�5��!�e��UA�T�ҎMo �"=�1�j� ��N��$���HÆ3<7�
���W�d|��n�X�4;a�����$����&��)#�^o�#�F&�޳G
�8���e��b��B
���d3¨ņg�=|�MmN��J�c��������o^=��y�W����q8Q�e�{�a����-�5�w�tf�ۏ?�J�҉�8;�0&؆H4�:	�����WX�k	�����db�%�Л��C�n�L\�@d���S���|��Z���j��^0ڣ�I@g�����a��:/q4.�d]�j]�����>���|����12vK�h����,�|��+y���^S�h���'e����0wo	�u�B�[�n�fu1}�U7�S�%�v����m�0�A�]�����h&�y�ġ�I��~����m8���́41a��#i��Kdv8T|z�Mj�ς�����D������q'���`l�3�oC��]�3Q��v]�̆TViq
x��=�20��Ы���H� ��п���5����5	� ��w�ƁЊ�`Ȣ��2�a,7C�v�^��r#�ʐ>=똡646?<D�N�3t (���yV)�˹�;�(�k�i~��=�<�O�_��J��)q�g}���cs���P�)��A0ScرM���Y�\����I�7^c�n�(�D/
���M��{R�\�����)"iɲ�s�4=�Z�%�L
�ĺ
���E�t;�
i��n��S�sF�@W#�d0"�5�\K:;p0p-L�����ihP7M��S���8�x�����>���B�p�9�`�
IW�	&�9�=�$^Ӄ.�����B���Y�I��4Ȯ���b_'�k�ii�����f�������i\_�H�_|_�u��{�]q=y�$�
��F�̜�^v�v���X�Z�pE�qB�rb�P2�
�e�+�P�xy![�&����~�s�h$."[�*���f��y���?��B�m��bivYed�$~'���X�?B�0�d	 �{��L�n3�X��((!e��>��B�
/���9�uӓ;8�J<�V�k�g^ۅ���3<�)�N�dƈ�*��ł�̡��O'�Iz�k�N �e���"�þT���}�����O�В���"����AqM�M��m�}��B���h��a�	���� �6a���vzHZ^s�P)��S�`��7��!��퉯0�g��A&���cC���q �v�������d��^�6��Ř1^L,.J����懶�3�x���Y����{�μ��A�{�Aq~��6�r���L�iNN�e�J'MgteU����%?'�1��e0�-�(�Z[�{��p�%��������]W�+�V~D�L��wu���˴�iD��O�T��o�T;����Ѳ_s�-��dj��n���M�f�6keG�N�D��o7������1�Oj���.�+VQ���![� <F�F�j� Y�Y�L�/}$
�������&�h1��]���s�Q��b�IH�⾭D �j��o�ah�nބ�3�F��wؾ?l_/{������<�q���C,�;póp�$9[8{J���y�:�%hf���
�|A�Fk ��{��fab����/5"�X�x�n�\�U�&d��;j�Ѻ��ց��Y�k�HP|a�-��篟Ch�k`׷䃚k���snLd�*q,Y�vQo0"x/�0�0b�����
�M���X�o�$����0S��\H�m^����/f�5�N;�.G�l�hٌ��`���c9������z�[���h�Z*#g;L
 68���pjӉέ:u6�$�7�M�2Y��QUێ�6>U�S{NC�ίA�ݏ�-��Hܪh;���C%�Os�p����]�Y>L!;��g]g�җ;h`W^ҊE�η;���p�u�������J�
{)�k���Cd��L��(�c���k���Ϻdb��nj[{��^��Y�N�aa|��>2�l-��N����u�+��z��Q_�x-�欮��E��ɨ({�*�ݥ��HG%Ix`\s�Gk�b�{�=��s!Ro�ޤ�R?8�&Qc�o\tOq(�f[��I23ܟ��^�>�{�U���,t��\S�R[|�;�+�j����p��3o~���&0f^�����#�9z��U�$�Bu3(^��:�t�S�a�@��{�S����zM;��dX�YG+�Q���)\��s	#��˩��0h��C�8=�RC�+�U�Qq8�������	#�P�|odn�j�5)1�`���Xv��)<����xS�ҔE 0潔�Kw��������\��믌$/ّ��H@'�IG��E��K}\OW=R�ש��/�JjĖ5�O�*�d	E'ɛb������$�	����o=Rf���ҹ��N�T�G��JE�Fsf8�!����3ae�Gʒ�蕔��U"�0h3�S��h�-7�U�!N��W����}-����p(#���%�A�m�GƆgi��m3>��(�̉�B/?{ܐ�\,D\�w���a,������/�q�SrSN�H�c���(qoT�	\p�̥�';aֵٞ)b���+������)�ŚI�B�Mp;��,�[���82��*���F�f��p�pHQ�BUubџ?}�>D4�%��3�dx9�!u�H��}u��ݮ���k�g��-�7;$�T�����8*4�ݐ��=$��=���R�u �h6D��B���ꖬ��m�݈Ra���8̖�	�wT�r����GB5h�ѓ[�'��5�#a�c����b��M�JO�G�_��vۚ�*g����o$�MO7=��i_,#�ݢ�*8��<��M8K�>Q�А�2�� A�5c�l7��&2���J�V��I8�OG�k�.�[j�Z2U���j�>�v
q��kM���I5�1�ᥭ)v���8h����D�Ԕo,W!��/���1+E��׀G�+zq,�����Q}�v�����|�U��uc�$Ai���L2�� o�C�򮾯��B����[y�EgU҈�h~�����OM��$�^a:���k{n4��9��z/�v��M�:dw�|Vg�}�:Z�ؤ6�+��:��v��-��=��5��M��ϙ\��5�y����c���Ϝ��V���T�n'&2ݓ��2�t���}�bzH��>!�eC<V��^�ưԱ׆$��Uf\W���ι�Y1�a^q�BWQyz�[V-���L( b`Ik�F�	x��vE��y�=8�D\�X?1���2OR��ʒW��Ki�@[ϒ�]�vơ�9�I�����e[xS�\{�=�2Jͯ�J��[���msO�����y��>��>*���MM�!>>����j�x��(�8�K�,�2����J���>P�xk]�7�u C�l�(���֪��x 9�k�D���(�f'�|���L��*^&��2����q䱭Jp��pC�ә�X8��7fNy\�XݔĳQ�gu���^a�9�{�Ck�^��f��<Kc�<I���6�r'mWc9���Zۤ8�]db�������&|��!�R����M�k߉�ʓ����74F�DI!N��ajV�d;+X��GC��{�S?n���
Y��X8C�&qZZ��K����`t�_&;G%a�I^$�㹧G:�Tq_Ŀ����=������cHF:R��׾���)�Ö���q�)�o�A*Mq�l{��Z,zF
$I���*i����S$����JϾ�c�����;�a�#�{�3�C&5���א@t�eb�,��Co���R��E{is`�j���e�~M��>2S_��|���Y�]��un	 u��)1�7%�m�N�O����*�lF( 	8
ps{q ���Tg���1x�I�a�@6������B<��;�|p�ZE4fƿ��.J\��S��T<%~~K��4�X$
wbiw����S�Nɫ��ha@㹰/Tv��hn��N/Wz�{�z?�<x6#p~���w$������d6۫��2�뚑D�Yxa��ڧ`�R�r�uS[�P�U&���ˬE'�U���]u�p�wl�֢3��90��tr1色�pMDuؙ:0�K$p�&vC�x|6�<0�s?#S �IH�d��z!6�$x3�ö&$�0p��q$�:`���?�����Zד�5Ԡ=���M�Bl1.��yf���(��a���7[}������w�V�����r��ն�O���]4Fڐb�̓��o��à�����%���I.�������<����{�kb�s�����<��l�i���e�1x�G��a�LcZ]e��"���o�]��:�^T2F,��EaYf�4�>��H�w]#3���o��..��M��� [�̵���p8�� G,ȵ����P�p�Mg��<DSYz��__^;.=�/&����R�zOxYK}J�x�^4��o+�B�k����J|�2�c�"brgm~O%uWXE��[w� Bv��H��5��n)`�y�D[������"���3Y���оq!4ELO!�x����<|{�_{�f��늉�U*-T�#ݪX*`m��A���o�AP�����ǲ-t�gG��%�9�kt�Sݰ�Q�ipA����Ε����X�{B2��j�5��*���{�6���,,���G���4��'��c�ӗ�o�ڎeP� ���C�;ڬ�������a�v%�GT�	�ar�h=�i�{m�''�*!w�oA<&��<�.=wG���C8�~ʱ[h
	�7�1�w6�J���g��kN&[�R��f�~�j˷�}[3���N�Q{|�v ߑYb�z�>� ��Za��4PL&����7�yδM�,�!��N�IwcNT*N���Ɩܰ��Tc���<��&�{_+�G�#D�W�v1�5���Z���/�S1��f�z��x�˚�=���
Q;�w�J���L���k4�QQ
�@�}�o��d ��������	(�*�]��e���ȯ����Z�*a�Z�v��8�ם	��� ��	;��,���uE�39��	�c7��ҊxO�h"��t��*K�q'��q�>�{��E�2����mvr:꺪ɍ0⥲h`�.���pXGL���V����#M�k�N,^���6h�&���l�֢k�5:��k ���;& �Ŕ�x�J���]�kz��!��&v.����t#<�;�ͷ		X���y�9������g��t��F��NX��]-u^��ҙLZ����iQv�&
�$��a͞m1��|�P��'��=~��Z�ۄ�=���u��AV^\ԻfV��k�c��/Sn:׊����c�+<�RuM�yQ�t����ڠ�=���m��4�����X������-$����q(��L,��g����=�R{4r��Pc��wj�G���/��1Q�3��&%|`��*_���Yd��:��N�a�'���b�D��J
Rr�U*�U������y��EF�V�WY�-�e��ΐ.����lb<�B��F��q����6���]8:}2�[��5���k��^M����W�tM�G]g�>aL�>��zLq��5��O'���%qX���D��{|���
����/����v6^������5�19���K,2ƾT��Д�����*5ئ���
A#`�'HQ�_է4֥��{�]����!����?�h����q��=^�א򄭓��k�I�v@õo���%|_�!N�x≁G)�+��{e[ {�5\�ă�R�?�$B�;�u��]��z���������=����T�X}�����̺����>F� fe{�u��#�������f{^L�p,�[�P	�h6&���x�J��{��N��h-�J�5?��^�Պ�!,��'$d�ZvyPZ9��Ƀ͵p�]8��,w�1���I��O���`��yP��q=6�L%�"qٻE���x�'���>��M8�ݍ)54/:���:p��Pv]��6�yPX��n#v]5�;�e���Ν�p����x�u��;k���FĆ�E*�*ʞc_��hbWrAGv
�(�Y+/�Y����ԡ�Ȧ�LX,[��{��"Wt�8�c����p�H�C� X��,������_�����p#D;e� ��f|VN�z�y�A�������i�M,]�^O��7��1n����͝��R����Hj]~,"R=�5k#L�4D5|�wxj�A1��:#ۉ��s'#$]�>x�!R�Vq���d#j��bC�W/i�<��_�t3����_����qa���;y�ʊ��5g1:�x��^^g>E���o�hӌ<G-i]׻��r�K�V��k��=���J�]��]z`�3�L��^�1O	Dy���Ax�`���:%��"��݌�ݦTkzMY��8+u��
싸q.���oӔ�37�q�n���	:WdD	�l���/Un����F������C}|PD<�d"*�*K��hM#y�P3bՕ��(!��Z(��X;�v�e3s<�Q�]
W-���`�/Z�M�u��Y�C��\��M�)s��3�� Q�cѯǍ
V/w����X�7�R���v���4Ѻ��u�����N����o{�2J�$p��eć��bB������Z8&�>����<��R��^����LU8]���,��J��k�C�:yэh�L�]��٢���k��G��BlF�m,��zR��ކ����V�>F%M�x�p�\SݑW�	Wy.�{D%˲�w�����x��=�c��:ݱ �L��UZ���V��o��8 ��/��gQ�,j;rI�� pq[�"�}��d���s�qm�]$���[&@��UOϭ(��:Fu�z�]��w]BH6r��X�p4�A%�s����1�mcFf�	��å5z�W����G�}�@D��������0�K%���>���ޡ�p#:���pPұ֡����n<���c�0P�)�%��xs"�s�C ���LNE{i1jܘ�纬�3��'	�D��f)ECb/7���)�ɪ������������6�ڊv�x����Ա�O�s@��!}y��Q�à^N稚�tr�juF+v�G�i���s9�3t����|����=�-OV/�rvQ�D�4�R���z�
M�+
�Nǣ4<��I���U�\�9��n)>�9hY�&��N�x%���Y�
�ǂ�6*�~(V�!��eS���ZRd��8�.�ܐ��wi�,'�eץ��^jIa��l�{�־�z���$�}fuǬ�2~�V��i���RNnQ��%3�֑���>*�X��].�	�8�X.<:m��|�ڣ�'@�����㲨���YO�.bWV{��v�{ݼ�]1����Sx�oh�u]���lFW��sB"/�&|N=�(�܌�K��C>�a�)�6V���2�+���*i[J�ب1�S�4�� ��A�Epz�9���W��䱚Wno�k��ʗlJ؜x;���.�B��'R���Xv�/����L<��'���1�MCZ�xLK n�*#�B:�ol'����z�D���y�����l�qr�PY4%���
/.]t=1VNK��P^5ܫ»���ny�j_��M�o���
��bO��s�Cz�Wm��ٍ��������Q�kUon%��O�n}�䅈D��`�{��H=�b�됯�Ē���6�C�0���X�~O��d���s��a&5��fzPc�R�+Ԓ�RK*ãɹZ� n-�I���^�}�QLk�Q�a���c��c�k��U�@F���H��5��Ns�#����H
m�'v�u�ڲW	+^�T�^���ȯKdC7d8kc֮
��C�.>d����oE���f���'�;cr<C`�Y&���*<H�7v<� �T���V��4��a�`D���tR�$Ɗ}JW-�ݲ�W�d1�I2�U��|�=�Dv�x��m_�!_��;ϴsh���דM�]3�tK`��N0�4/�	���!��#N�4h�K�/lA��=hĂB�����������RccaVK
��C���d,���b�l�[���g���	K��i7�̸��FE����QmS(g������A���97P�2*jTu��)c��H��H|>^��M)��DL�H���u&��uU;�[⢫�yW�������u��a���r�.*���?��U	_1�z���eY���cq�������O5��ʳݩH-kf��e-�W�z��������,��J�pZ�*^�$^x���]'N�`ϰ^�o�����יִW���x\�����3E�U�A9���������(a��wQTIUb(��{�um����hC,O��������&f���w�%�<Z��/ۊ�|l}2�՝~}�V}��
F��/@OJ*�>�IM.��=v�E5d�����O��\�ᑋ�����4�u�Q2*��a�גX�iN/�]$�G�b����eᬀ��|?�ȼy2Q�%Nil��
M$- w��SY��rR��m�� �sd�a@v��V�����{�YӮb�� I�s%�nTqBu�z\��6��w%�vm6�&jfU�C�%B�m�a���5ծ����llx�7�[F� ��-�?���X�X1�Us�^O�`��\-ڲ�ڶ�e���.N
���ľO��Mw��U�Ȣ�-T�w��o2�J�p�rl��N�:���;d޲��v{J��^�䯖��v��E�\L2�9(^�z�)4f�[G���S���:]!b�\w9��{��.��?g�1x�Kh�^�Ě"�mL,��s��#�X�{���E�#{j�&L���8�4�P0>ꮤ\��6f�q���Z��lp1pYM8W�0�ˠh�&����%婵���w�����i�;/�%Cu��|%���wq�_g���r�"�db(�ǩ�剕�!Y9�)��>H�ԩL�T<�H�왘Xw�p�kS�V=&f)��5���&yb؀�2���C����{�?��I�*K��9�Lu+��5��R���I�&���<�R=��*��Eet��4�0wY\eZ�̅�ǽ�}GZQ�d��1S�g��V�xA������a������9��)�:�L�)�s2g�J�(��^��<����4�Ri�cޗ�f�E�h��:7�z��-*�̵۩rN�n���W��R<��X���1�Ӎ�!D�1�HbfDf8��~'Ϟ�e'����]���N�PP�g>=})?��S@](|	�-���-pO1��-_6㈯62lB��y�QU�����U>��J��HyVcj�t�@eN��	N(��-���1%�����R!�bj׼��z	f��Z���z�mZG���U8��j,�C����z���[��l~W���3����5���"�޸��*<RO�9��r�2IE9���|�<�úg�-gp�Re�lH����:��u�Q.�����$�	�#}s�E�M/�y��fQj�p�5���{fZ���@wI�Q���cV�"��=1���/�ѳZKT���&�H������:�Hx\�����{�n	�A/�ӎ5����v;|�1�HAW��ޔ�R����`Α�|��x��G�;��d�����2D^��u�z�j�=D~e��" x���%�����k�N�a����(��|�kQk%W�6����$�̛�7b1��K�E�:������,>�,��ƾ��~(���b6bP��厞��"ܥ�\2�/���:#Y�.��⸖���qL˭mK_-fRiHb'�G��z�)�e�nkYwe�3=�&����֚��gz69s�`$3�!q�HD��^d�'�f3̣�������&#On�@p��{�f�XE�,�kk3���`eҦ��;��}��p��1�>�o�`-2�פ_i��&kWT�,���;g�&�tà
����
��WKV
!�����cTN��/O�<^�)��������!D�Yy�x�S�c�ba��M+ӣ�S
3�M� �5'��ʫBpư����>���'�9e���{��[�=y�5�1(1�z��]�~X�O�"!�j��6�����u��f[(p�CD��F ��u���V{��H���P��p��|G�1��	=��S4Un��?"R��<�獱��;&|�����բ�QXk��{eK8��(ʜjR覆o�g����I:�WF�r�c_
;&����N>{��7tÃ�9kW?v]��5��k���AM������k~�x�Y�лo<'������͓�Mr3=���3�h��0*+,*P�%���D�T�f�(=���l}�d��SE����V
O�7����!��^C���OT'���y��}����S�L$<Z'l���{QYtZ��6����7a���N�������P}�6���]v�]�,�"�|C^��{�X�_gO�jD��ט�ǽ�/+�w�^��#��yR+�t������PM��� �e����t��a�Gv�k���u���N=��!0Jnr�!�Ƙ��̗m,��s��0�ͪ'\@�J��������)Y�!��J�b�0^ļ���L�i��RĂ���Um�FE��<�kI�a?���!a Fe�����y��w{V�BIOKvC�UC�C�8�ҹ6~�~�!���J�anΈ��&lF�© �أ��k��ߔw�.���E�~MZC��O����6?m����ln3&¯����6i(B:O�DTU�u��j��Zj��N7�4(��oY�k�4�z,KU#ϧ�݄�.ٌ�d]�dc�,�!�p���ܼ�o~W!�^�>wG��|���� wN,5"֋�s�a�V����.K.�ҁk"���Fqz�f�K[6�w�D����+U��4��}V��[3�Ъa���K(�������k��=�p�S�l�a�uJ�플�e[c��{��ʟ����F���^�u5m��c1f,�}�.����RT��#1����<�t,���K.pX��rhN�y�/݋�
�W]�!/�VO�EG�h�R��B��p'ެ�*�&Ml��'�]��`7�$���O��6�N���x��H���,�P�cq%��65Th ��V�֧H���Ed��䆯v��4�����7�bm�4���������1m=S���#�����yu՘ti\pC��g�,X�e��du(�r�>��j��H:B����C5���m��9�W7]���е�ӛ��2jS��r�u��F�EQ�p�!r�T�c����J�N��
sU�hW,��&0�8u�O#1Mt(��c��� s�@w��'�pN9y�Y��!x�8�nW�-����	��΋��a�J 8�/��}�����9U���8iA�4ٻ�G$��v"��k\�}W�Fd���ø�jZ�q�2
�X8���C|�b��J��,�i;���B�Qx��Û�����b�5Z�`�,W�.�!/�n�x���y�0�h�8M)���j��lc�Wj���P���q5s�K��-ڍ�k^K��'v��N�b]b�E����,k�*��h�* ���:�F��TL�����>�
����K�o�W��4�t��H����j(CW��S��J,uPwԙ��W��K��׏zf����ߵ��?ڛ<lCj:AhQ�)��ȯܫ6-�g�?p�CD8���A�.''��J��E�����~f�R��6᷺�kaC8��pmWU�����W�˩�OMF��.!m��C�Q�˪�IFuJ8�%}���Ȱ���y��B���M#�0�ُg����B��rn��}��x+)^P������Ҙ,/h��L���A����A��a�E��n�:�1h�2��V��uM���x��Am-�ā����� �2�J1���TFɲL�u\.0�E%����{�b́d"���k
�Rq\�22�7&�F����6�)�����d 7���Yz��ż阌�A�P�e\E\��k'"�o�j��
tb���M�C1
:Y��YT��	$mG�jH��^@C���)Ա���a��U��*��cF���]Ib-G�n)		�g��Кmd�p)�����ְ�W-_��_�[���-i�-{��%�k���=��1��⃢�qx���&=��n�� ����n���E��y���f�نT���ر�g�C�Gڋ�%�8-ѕRl�uYű���y��)k�@�b��N�v~k��f�=)6`0>���:��瀿PCp�Ka3���>�(=%��3��f�Ӆ����5̵�q�ILS���h�Ø�@�1���>�_�����X`��4�_�Iq�>�
����U��e�x��8�f]k��V��:��-5��e;�m[W�o��}����5��k�I'п��Z�y��01���rUy�"���%%oy0'.W��V�(��[ɚ�5���F��$&z����g���N-�6e�g���$f�N�揓v�9m�
tW��P�ڌ�5��/�{v"O|v[�(��~���Ȅ�@��Q�Z=�Ю5$�����3V8���i�n�>�o�����cӷ	�jn��GZ�@����v�Hca	����=r�����Y%��aEx�
�%�$l���cO��r0&���=�@�o�`dFu���'��d���%��j�96��k?�4���z:��V��O����:��Px-a$�&��l�f4nC��ޥ6[�*&Z��أ�%����)E8�B�CK����ZT-b��\�����،�.@�CׄR^G�Ҫ�M��]$,��l���L�y�h`�����Wa���4Yf�-���&M�5�H�H����T���X�sɫ�ѡ{c��}���=�{i�rkuŭbp-�,�/��PT%���A�ҳ3�)(i*, Z�D��/����WW�i8[����*-ks :�s/�I�2��pT�Jv,��uU��W�������)D ��wa*ٙ�ὶF�WM^~�&3_߼G�gB{ߴ'�$6����7�S��F(�bRE������<�I�GX�� b*/�-TH�`IO����µ��|����|�og�VNJ�"�_�밢�Z�y2����qo����d�{�oV�M�'{�^��]�	O~����jVK^މ>,�$�0<p�|����!N�c������Zk���	��ϊ�v�c��`��Rhܝ�ˑ�YM�Y���H�Q���(�ۉ�*���ZLt՚��_Q̔8sSFo�Q�����j���IJR��
S�Xq���c�(��rwh�=�L�s&9ZCw��W�۲�`�:ו��u��ap�0�>�Ӊ����6'���4Y���)$�6��F��r��[�ŞpzÅ�Z���ƿ��$[(��9VyUf��	2�5��Ŀݣɏ�4὆�%cVn5����z�I�E��q�ZX���HKNX�������O/ϕv�p׋� ���]X굗D\�xG�+mHټ���K@o�Bod{�L`=J��I�V,�R��A����N.���^�x�2s�Ϊ���7cr�|XуXR����~�������B�k���uS�k���$�D3�,�ѳ���DX�_>��:d�߽}������n���g�)=?�z�@f����$���cj�6��!]��'ʚ}F���W���g��:��:l�5��Đ��j%[T_��0����_��&F�A�k�������n��p_&�#|��R[�_����Eq����(H|X����F��1}*{��M�	#7O-L��A<�5��*�}�����\���=>4����߯w���I����I�A��u���[�)YZ�]�m۞ؐ&�D�C���/�m/ڞ��c��?}�֤���ʐ֬�-zK٩�E��^���2��h���ɛ.V	�����$��ca� p��zz��W}��d�J��;6�E4$���=���(�K<ɓ�*�`��A�v���7i��ITx�#-@l`���W� �څ�e �]0ۓ.sS�RSU���]ӫ�CN��4W���,�|O��*OМ�v�2�.�����s��
��oa��1a��&<�ɧ��+^g�Rk7�޷>ܳ}F��^��J"��{j vE�G]�m�5��:�p�H�!�Y�t`�2���ϱ!(�<�QÚN��|��Q��Yһ�BQ.ZH
�b(h�JJk���"g��]I���3¢��tĭ������azc�k��#�ӣ���E�����ޢ�`�I_v%-j)�2�Z��۩�K8W4ص�i��u��Yts�c���_-�	�i��_vk��WƳ4xWJ�@��Q]j��J�PV��T�?���±�rg�M��tx%ʞ�(�67�{�g�A��>��,J�_�����L��~��&��<~�m|���D'��J��9�cj9_%���%�>&e��Z�W�'�-ԛ ��ϗ:ָW�~w��N�K��kT���W!h<��١ .�;�Y�b���O�ɳ)��v�alġ��lQ�)H��1yj�.�$U ���B*��B���b�쨹_�o&�H��MY�� z&����4 P��A�>n9�ɬ�xɇ��b�Q_���%��ji7�A��Aǵ8#��h�]$��R�/
��@:ņ�t����'*������O�c%��]�?q+%a��#��,����کo�r�F�ڙp�i�=�t�@=rb
���ӧd~�3#O��(�|TH���O�FC�C��������R�����ب�k"{�R���kRv{=�ad�P���5�MN5���mwG����ҙ8�buF.i}5�6���^e��W���F�I���W �2�^��{w���P?�֯	�����y3�Q�=��DX��G���ߔ~�!�"]�.�[P�6�O�2�Y�����>����� �UZ�;Ȑ�HSV�B���A�y9�*3���1�>�]�n4�U��Exd-�;K�[K���Hӱ&�����2f�lƲ�Å�UjBJx!{����AӁ���8s	�Un��nA/�	�c�WV��6��]W�|R2:({X����v��Z0C0�Qʌ�vi[�&JO�@�� �#�i�1�Wg�����*�q��:���;[�&�>���#"ϫ��?*�(&�&q8L�6o�rԡ�KU,c�&ޯ��P�B%�U��Huߵ�m�u�Dy2���&��J'Ls(.[���*87�}�Fg�Vޔ��.�V��Z���eؖ�t*�Y�5k�R��;g�>��߱�u瓱�Qz���qI5��H}�Ixd�|��WjR2�[[�2LiN%v�>C�e��劒!��`�]�+�����YU>��|&Y�5���+U��M����a�k�o� �#�͌j�a�������nI.�q@��t,��'N}f�Oi
'G&�#���m#��_�ەr7G({\#�����>W�Rm�.���_���̿�՚#�U���A�5��&��;s�GpTw ��~��.��%s�a�<��Sb*l��Q��[{h���G�w4up�?�ˌ{�������> N����c���Tq������L(�`�}����k��1��Yk��~޻���vdL��zN�ߝ��`<{�]T��Y`��c�����}FC��!9��3�;/���0���]��X��O�iD
\��P4��н��ߗ��`f�f���~�TC졖�RF���Ң�&-.��!bN.�C'��d�mB��
wJuA��9�,������X�;E$^b��f�
Nv7���z�]gע����N@����ow��x#�����$V��T�/��u��ș[�WKW)�X���G�B\�a���YJH��lP-'F��]l�����_����x�2�����}\��vVoX�zK�x��
��kv��0�W��ɧ��:B'̾�=��	Zp�"���D��=�j�m�t]f��S~MV��y��ૌ+>J��T�p!��C�v�]x�"�TY���(|�Gʱ��P+X��.�I�$vk�[f�W~6���1^�É��5qVg�]\	��H��\v��K��b�L]�A�O<q�X�6���pw4��d�W�L]��d�4E�%�ׯ�ၗu�3�{k(�p׵F)�h��|��<<I��\�^��{��o�x�L:�#��R/��nc�'1�eN�cO�X46���e-�!���J-��0?�#����!�[���=��J
X�)�+@Y��X�g}�<^Y�W�_���s��i�=��P8�v�� T�Tn/p'tR�II��a�l�)1�(=,P��� ��Z�!��D����7��L&��o?��'|���}uH�A��rr��T��Ξ3�!�����eb/2�s
yX~m��1�u���`�OYpb����$���=��T�W�*t������^�`�r1�W�pMzT���1�Ga���yʄ����'Z[THlWL7����5�Z���=Fٮ�9չV�ti�)L�r.Ge�5KlT�����h_k��^�"�(7��б9�����u/�2���3���L�H���ʊ�X�"�I��N�α�Ux������h�c�u?ġ\J��u��2����hc~���>���Qګ.m��:>��_'�Vҧ�������rQ@�!���^�4��]�@Hp����j){�֡�g��cm��bm2*���������Y}�H���y�ʂi3��}3pMY� J°W�N���;�Ђ�;�@:�q��7e�[��5��6+���k9���vV�F`�+z�WT�yLT�Q��`9����le
^ʚ׽�g��ݡ�dW��Iz����El�(�KO��J���lf��Q����ccٴ�)�bp�,��+g��,�J������b^�\*��ZoaJ<�uO�C�n�hWҳ��/湫(���+�r�5���h`�VN�sOOĒ�^߮���-��/���<�a�0�Az~*������;b��;@M�lFN���\�SVRU#�1�����q�غ�U��zZ����H*�R�vv�QT�I���hWvE����ʳȠv��w�B�gu�8W�0�/�ad�6����׀Ȩ�&�����%�v�u��`ɚz����L�~8
LN]v�u5ު�C����7��t�����:�g[��U�����r�����~����z����WU8��q�XǕ�A�G%�����r�$�Eq�MV���ր����r20x.�+�e�"�(���.��n|f��n������6�P�Eg{O��3� ���qW���-�V�R�x�N�B�j�j�t(MJ[�
a^�;�F�uX�!h@7ʆ9�����"�b��� k.&:D�|��һ�r�y��Z1�"��a}l\%�\Aey2�w��-ϐ0�1�NQ���խ�ſ[���3�Ɲ�ɝ4AyȄ"��k�e��ϯQZ��\�`b�@����jed�]��k*�ʬ��ޙ�[x��wmw��2K�����4-�$���u��	����*#{�UȈ��jL��~ތכ�S'm�(M�����.�/[�������"E}f�}�y��U��5����oa��ر����7���x'��)�s��V��2�w)�R1P%?=/������#���G��s���;�Z�Sw�z��#�]������ꂉ�\�r�a9�>�k����ˀ�69heB���u��}�.I:g�@}��Noyn����%�̤���]I����T�-,����΅���@��̃�ix�xN�<; Ng$�JI�0f���DBeύ��֒F��	zi}aȖ�Q���>.����Iw���ғ�����XފJ����!��Ɵ��T+*��SV ��g'�M�Ë�ܪ�Uz��]Զ8��%������`h0��y�l��y���G��a�o��S�~a�`jԪ1톒n4�7F��K�͎���ǌ]_��<w��c�S$��zd��h�)A:��;�{���W������*c��rۀ�u���ǜ��������8�=�JeH�O�;Ц�\��
]���h�`��9�a�M�����n`��0���V�i�5��4�4������P�<���V$���&�w�v�2��u{�[����(�"��������҉\7���MhR�W*��XC��v�r(&|w�bp�W
[y�TI5��Sߥq�ڃ�B�-��k��.E�9��Q��64؈c��w։ff��ϝT�FR�8M��5��P�;��A^(�.czc�`ovS�X�Z�$qm�U����MWI�����|�!�� o�vf��T����|!�c^خ�6��C<�=K@)/�a����Vb���l�L���smS����U��k���a��`�H:�X�W�Z��+�w�q�g���;+���T�ٱwה�D�*-ؐ���hZW�{�r�e��өn��;U�R�x����7���|��!�EP��ۜ��4Gq}_�X�]g�� <���,�X�M���/�^��:�O*�މU�z���O����3.�1�u���1�꣒U�U�K���ժ���b�4�.��Na�t�!u� ��s���Z}����=����$?�W��"����Lы���DI6���GTl����/p�_�n-�}�T�I9dg�Y�u�!*���ֱ��$�H�M	���6�-��>fe�Y�r�GJC
lu��{_�NMۘ�FI�P/Ah�K�z+�/�{ZtJ�#*C�^�q���I�H�!y讓�XzP>��p\��Y��0lw������EU����ݗ0��z�g����{L��ue9�׶��>p\��_��ܳ�;wI^�Y��Qҝ0s�!<�E�NF���:�7F�	����WľP4Ќ��J��6肊�"�6PWm�}^��~� �p��3����)!*�NVmYx�o7C�����|��L?��S���ۛ��n�����	����9��g?'n#���`���A�{R�G%�;o�W0�_������z��<��x��5�Ӱs[��lh���2�Є��1�d���(�t8�|���4j�^�ڵ�h�\m��������Wu~cP)���0ŧ/U��Τ���N�8d����x]/5qBos*G)��|���f޾y����R{���?$>\�g���V��}�ކW�\�<�
�'���p��r�ȐJ$�
��0/�O1�0j�-N������~���a3d��fj-PrP��}����N!�Zq> Qb�ڗ���Q���岴�Ɲ7�s^�P�to��iv7��D�!������j׀U�1��sh�&EK\����xL\2*�8bp�#�h+�o���W���Պ}��U��Ry�v@-����x�1[-פW�8�0�n?NFE�'޾�uτ�SR������GBzO�_y/�E��%���c�哆1�I�4��?���ۯi��9���7T��t�z��I�i�ik��͵F�N4��<E�Y��vuOmM2f	+��7��WiFV*�Ҵ�v���n'�Vo`��᳼�Evy	ٚ�lOq%*v4U��Pib ��Q�]�B�5�Nt,hj@r�Gk���9��x���u��5!��D�1^>��iJ	-���u�lI�N�x�yI��K|�b���(������0S;g�"9�z描��ݷ�E���qd��D����^e���/5�p�P)bnҤ}��J���UICL]QW1���g�e�Ϟ�AX?�:�3kG�bm���~	��0�1�`N\K�зrX�	��t_I�!���m�Z�qa���A����gy�c(vUϓI-�=YSC���"n�\���y��9$��B���r�VC������r�����DR����o�h��K-�#a�`�H�w�-k��Ŷװ�0�Ad�U�F�5���_�Sݐ��7���I�I5r�Mo�}I�!����o�H��r�.i$6��wF%�B���� !d�W��J�XP�F�P�����x������C�����Bk��x_>��P>~�(���~����`�<���w��o�-�����trN�y'��YO���!T���*i���fm~���9*N&�V����ph=�K�e~�¾������]D�0�x�W�c.�m��������O������5��>~�@C0I� Lč���+��o����p�DT'>|?��q�I:F�U�0ø*������S������l3)pGa��ˇ�C�Ł���p���Z�!�A�A�������"o�^Q�-�2�~�n��T�O
����ݽ���j��|Q�5���I�I�G;�ų[�pZ]&�H�׆�Ѫ�!8��u�'S��r6�5�kCK��r�0�6l��X�&�/�H���`����������������oY&������{e ��oZ�_7�~��(%=�4����U�����Jj8$���gu_fZ���{N�Y�Qڀs9��5�qwҭ�?io�帑,n�Y�v��˻s���?�ͼso�%�T[.\@��[D0�����lfe� ��p777/�je��e���UOo`5�Y�,��Ř���y�(5��a�nb&�;7'KL�w����n�~��݈ޣJ�!�I�bJ�_�zI�F냒�ݵEg��5зw/������<FC0�x�d�e���׮⼏��6�&�_���T*��?E�80=��yO"��0ϼ�q�wS��{��MNn8��>`m��Չ�� X���Y����1O		�������<y	87�;trU�0��z�]U���\,�l,蜐��g���C���;�֕7�.�����ʅ򼷷�^^���v�f��%IL� �t���J�V��@
]��� &V�E�K��4DS�V�~��q^���>�CFo��x��e`�;��S.K���]��(,Թݵ�
�D�ƶ��ҕ�WlE�ڎ~��V��Ԧ��XH����wK���x��ϓ����ؙ�DλG$0l$�]7����
��fc��j��I�gJ&���#>��]�1��R�`�vY�x�#�������W���^z!�|��ۤ�o^+	�{��E�EY�DOlOa��$���#k����y-hKq�(�\<ZzzOG��^B����onI#�cѵ�eT�]Ȱ\G�bO1��"|��O��2��H1|?I9
�ߑw+�&�����X��z��=e�o��l�(-p�g�wi.=�$�'�B�&i�n
�޸���c��\�1C~�Q�I/QN��w3��O�Tg)�"�a�7$C��A��<���cn��B����&�^/N'�%��L"��:�� J`�--ўa�Ǡ�B�z^����B�s�D�k��m��Ebv����r��1��|a.���8E�-Q?Ye��ps�.P̬�Q�n���Ι��B���{�ŶF��xJ�>/)�-�i� �l#���9Y�ϫ��kv�nW?��Klԕ�ƞ�)�|��C�#Z%S�1�ֱ��|���s��;�;:1P�u-:�?��}���b�.1��r(�&{��}���X�����]���%��������J�Q�&��>|�A�7�n�_�|�L"�U�^��7<�.�X&h�_M�=Cg�?�{)��׺�9x���M���	��ŋ[rH��@z��PD�Xũ�f���������F�'eT� ����`nj� �-=T(*9��y	}?||�>��{��&^ב�ZGS6\��F�U�GM}^&�)z'9�c�;m����a,p�`|qm���J��qz<_,���y��m�S�p���b�l�wN^K�������uЮ�`�R�Dv��+VD��@CH���������SRiK,�:��=�:	f��a
����QYk9"Sx�؜aH�Q����=U-��pJ���Q��!'��{R\e:fC���S���~�]�%�a��p�D�� 1Ίs�����^�d�+���9i
T��E��	<i�x�T���Y�^�-�']m����5:ӐV;��M�l�]�`Xw�܉�-��� ��x�[��!2�S�G*x@��-�gL����#V���SH���ǔ�iڎ}�1�d��ݨ���M����/���M�>e@!j��#���o<Gx����+B��8��n,Jߞh,��?��=�����~/�*���}QB��h@��c�G
e"\���=>V��rC/�~lw�v����,�	^��~�Ţ	!>�s\������o����n۱D �c���M���w&�p�?���'lD!����-�|E)�]�U��*�2�9�<�����#�ae�}�H��	:"�����bQb��@d@�Ї԰n�>|L���W���74·	�s�U��zcvȶ�F�����1Ģ�{����miC�4���A�ݹ#k�tR~T8�~LA����(X04UwЊ]�v=�܎c>�~�N�M�%\��=6�}�[��;&os��/+�e��9�i%B�&g�M۲�7<�� �>ĺ�g�w�r�X��-�'l�7���f F�w�;�99�k��.*�9�:?�y��0?C%���<կ?��SJ%{{���n�x�2��T;�ɑ��"�w��)ė����8���U(� �]*e�s:��Z��C�"����(	�{�����BNx�x��������D�u?�����;>0";�T�םq���ijڂ��+ZZd$zi���?�g����W���d��cū�嚰)�v����.�GD��O?-����IK����!e�7���m﹡2`N+�l7˫��+�*���>2{b���1�_�1%�S�G�X�⏏bJ�C'�-���cA>>�>1����ȧT�A�[��
�7���נp1�E�\�����{�J�jYV�ʉ�����2�Wq��n����pe��8i�xzZg���_�{;;ic�k�5�B� fCk�O��$];Q��	{�L�G�q�%�����wW'	}4A�D5_"�\��3a'���1��,-��l�y���E;3�*��D��l�y|�q�V��B�)'��J��-�X�\v0���o���6[�s?�~s��J��.�֢��~4��B��T73�S(�7*C�wm�1أ*0� �W�ccq1|_����_��z����aL `wL�8�8�F�=m�A��&g, ��Y[s����d�g��q�bl'�1f|-D~OC�ب�tՂb#3�D/
�Ft�Sb1�}v��1)�^��x�{�͖s`Rky#�f�&y�H�L��Ѝ2�0\�7�2��x¦���^�:r}���%�X�G��~Z·��i�F��"�!�EE���hl:8>5����M�Yo>+q2�ksFXk�� �����y�]�xo�?y3�|M/C����Y�;�1�w*�#x��B5s��7��u�y/��:X!B
�˙a�6� ��5D���{�C���ыж!�=��xraE�(i2�p�po�4MIf+Y-�.�"��T�"��!�u�"RD��xy���:[_+��F����e,��/�Ϥ*��_�;��Z{c�uf�Ύ��w���`Rt��~uU��^+Nv��`�_��l2o/��Ljxv`(wg��2E�,_#��f�ey�K�i<rM��7��_:p@y�eAX����;��y섛�����L*OOr~�r��mf{��J�um�3�aHʈg	G�݋.�� 煨�bD?S6����cj̫�"䑞X��ǻw�;�K8�٬s)��$/��KдC��F�&�� �o<Gb-=/<؋�<�kLṹ.z����y	M��y�.x���=���4�i2��k���8����n).S�԰�F�X&�f��5a<��☙x��mDfYZ2��cz)�R�+�[ݓ� xa�xi�J�z��2xrH6��WQ��S�LNFS�
�B��gr-c���2��U��GZ�\���#��NRTV�.eCz}M)'�T������	�����T��si�.H�,kВ*�l��nV�_��7��������=��h��8�?<�B��Dty_x��n,gv�s]�o��1�&'�����GQ�Ty˓��pܘ���7�2K�b#K�)佨C���B_�ÌZ����X0"�u!ϋ�7d.�0��Ы�~�P�q���<��z��sm7��Ԙ�t�=4=�K�7N�F���*�ι�f�,b׵�E�e���$2*�_��7����EL!�헋�UE�E�^yLMQ�r�Vx_�>Ĝ)�ӻ̲�'�w���r��L���dZ�9��A�r�<n�ϕc� ���.��!�����E��?��k=Mj��j�*R���M�w�^�g����ѹ�1�xN+4O9��b�Xm�}Ӛ&��F��_Z�#	馀hi�4�L��|��1^u0��|s�6m�i�N�R02l:�U^W�t����S`�K�����쉖��i���K;�Ͳ�;�������{M&��w��.��09�AF8��M"N�����!]#�O�OM�XG+%s|�P�#ͦU��E��SЖ��!isI'��u��P�"�'P;㚝�%����i]����*_.�A��""�4n�5E�������=j�#��Q�Ѭd
զI��U^�|�.X/� ƄP�z��H��
!*iR�J�c*�p$�e�ƺx6Zt+��]c��n��Z&���a�?�����_���{����{z��5y�H����d�Ԋ�c���<-�� ���a����
s7ߟ1�Ѵڨd(�.�Kѩ���;����iP��GF>�Qr�z���<����������$���-��)�,R	ׂ��t�!A�k�9wI8��KqJ�~�\�܈Q�	M����/A).wI�z�[�SV͊�t�x�!&ݏ�X;�<I��.��g�ꂻ�� �S�.�a
WX�z�;�Yq�}³�8IJR�"5�$��F�{�Q��E(��}�/l��m$����5MW����gc����B�-���1��a����v�^�D���� C�
$%乖֨nP�kL�nY8���ь�s�lK1L���F�x��` �%�p�4P����}��t�<)ک��[A�gM�$���N6�5gj1��!킃��&=!��4�Ԣ,u�g�h��0�'N*2
F�$!��0<,=]�yw����FS�1P��uC4M��@X�����I�Y	���:K�����7DR
�������_�i����p8�-���B��$�1]2N4R��Y������?��H����].�w�Ȭ2އ�p� ���>�cj��9�3$����� ��p�����&ϑڸy�0O��r+碞�� E$�Y1��̶��R!�He�EoL�18��\ٷ�Á{ Y繶nn-�<��@c��X�Ѐ7��\Z��^��Q5$ش�1�m�3�uQ��t���K�F���Bt�ק�V:����P�:2������]����6��o0�/=��p�@%%a���nc�3xͤ;���	/�\J$<���=��Q�͡1�F��e֏"Ja�h,�p�2;��q�����ͳoS�Aۅ�!�ζ"�z)C�0��`����D����I}��1Z��Z�6�͍s���4aD�!�A1�Hq��m��D!p�Cx�����E�ۻ܏�c���ӕ-�8@�z|�s0�i*���ď<�˘�4Y�h�n��JeAEB	�o���x�2����i�x�;����Hu]��t�^<ʮ#i$B0A�}
�(�t�c��'])�F�*C]|GT��﮷�t'+�S�S�Im����;�����F����*��+��S�%�D�/�Br�O}Mycè�[[�S���  ��IDATPYe��h��(;1L>����� j Mlw�ˢ�c�
8?P��i�P��>VGU�U��1T��WٺK6��IY|9l�i�b�k#aZ�;��R���Ą1�<R�'9��LĆ����
����S5��l�$�s���C�ɆT�+)����R��\e!�����`pQ�O��U���z��J�[B�.>�Lm>�%Qg���h�E��7r�����6T�����{�8��Q*R}�<do��.��&U+�QB�H�4�������+s�rc��n����+��C���Ix��1�mh�<!h�/�7�Os;g��CC�-w���i�����Cђ���@"������s8./�H"�l�e�A�ܯ��8L� vL~�7Lz_KA,WG�a�yN6�l �5"��JMܤ.����g��ңmb���عbsC#���r�y5���)a�pV�a�jf��9�?)�L�@���K��Q���*�)'�\����<4NY&/�h";�ceg&�R, Ǌ-r�_p�\UUY<�<В���񼦚��\]y���Q@��t��UrA�RdQ�7è�NX�#���\~n(���~��=��Տ>=3�_!����_3�ƭ8.��*�,��5��h�4,7�B%���e�:��ء��1ӂ�KS��j�I�T%̬~�0�c�cp^ �Ls���[0h�2����F<D�RS7��N���2�n�^�e �Cy��2Kn�����e��FoM��y�<E,����\�&V_���$��>H��l0ɽ��Y"M��%�x&���!��2�����h�����C!����j�2E-{���)A�Wu ��y{sԝ�Bd5�&h=8vo�d�%�a�T%d�ם8/A�K���Cήt�uRr�)�*�����̕]pIY�f��eq�)Z��#h>��4bZ��
��C�����Q��%������cN�D�h�OA�p�P"7*Ҕup�	y���f0�_�����yj����aqx0W�~*Q�γ��s0c�Ic�� �E`�e���ju(^�`-�]�/ �#3dR.]m�ҏ͑H��[��ײ�_V.=���{@��D�3rM��4Iy�4	�^�=�s!b�h�	��!�X��vp	f��c޻���r)����:��>F��Ꮼ��*��ց��.o
���X��OcU3�(/d�b�뙮i���l�H�mB�t�F�'���Q��l��>�0��ȕ�-��J�c��X�zS$�0�0p����:)[�!#	zh�f��,C����TBAD�aB^P!�c��j���BCm�%�6�V�9�t�]�O�t�u��G:���:xR�����KR�Bų�u)���|�U����������S�iˌ��j"q%�PT��[{�1��pO�㮚j�҅��^e���H����"�@�
a�ŧ���6!w��4#a�D�Ou��,�s|�b�s�����]y�}@l�g&�wxٗ(�H3ƁT�h�q	��y����D�C��Y1(��lt}���x1&P}�z�!uCL'�0?��i�y��Ќx�)R�e�g���{4M����C{�S�*>A��	�H�x
��|�OX���/�Z�o�ʕ@�020�o,��KN&�Γ��N�v����YgC_�@0�����L���sL4z�{�L���w�sD����e�m�<�<>A��Y&"����B���Jэ�^"5=�>iLa��H�� j� CD̩����kc*P'��|���d=fa6�^?���1��	���af	�"J�`Ԕ�$��~�w�oB�c�н_�S<E��0�i�^,�BS��2yPG߭���|�N���x�00>���E�בOc#�d���&�Z'��k�͉�)6�>BV��8���x�S=���
%���7��|�??���it�����=�(�;&h�I��X�#˹4��ײ8�c�^�����)��󹌻���	eVMEx����d�x��[֭�t��]$�����׃ǣjXE�%ʙ�F�+Ӿx8�W~S�Oבy=z�oz����3��69;��A;]��^X/Z�n���@�'�j�M٧�ꬌg���̬i̝�R�\�D�Վ��x\�i'G�F���\V�����	Yw��7����5�����8�q����Lc�p'K_c��+��[NkVbWF=;�c����&&#��6�Mn�V���r4k�`ln��{���>��2�i����֑H�a�4���[m��R|f���(�����> �3H���G1�i,1�������K��^A�qoY�~����L����N�����)B7�{w�|A9DWRs	��ep���7�T�L��箊���56�ɂȎ���"9�8o(�xV?(���:�6��q���r8P�����Lرtr��,|�A��������R����e]
W�̈+,5���{{mug�����&Z��R���qiOm2�LF���&�Md�\L�w�����zw;{���K�38�)ڀX���w{����pw
{�a�c|.�z��^�Q�8Z��([��Ӹ��i�d6�F?�������8�ӕ!�������m�x��%+����U;ߵ��m��3E�e:-7'��I�\�C��"�]��4������_�_��b��u�0���ls�=o�A"��8�2!`��OU��>?��+{�\ΜH����B`g=4���2�P�R��Ezё���x��s�XtQ�G�q`��JT� ����a�~��0,��I��"�B��,)�O�/�%��U�2zq�0��p�3Ce{��̩u��y��p+�����ł�y"C
/_�u�lH�4��(�u)�G��U}���[.2(����y�P�8��>)ǿ--6�����0G$��ݍhW�Qv��L��d�`8Pi+��j�"�#̇��cA�����~3�w�$CNY;u����9����p�b�Tk�-<NC#��ǵ����
�w�tn&�%C_E�ϩ`��s^J97��.��8.�+�dEG��$�2K`��M��C߅�9�s�J���9�a�ٕ���SXy�_rb�3������<R�dʡG��P�QKa�KX^���b�V�̸�B�C��R��Gw���u��U�����	c2�uj�jX>�x�w5���I/�!�7�YO��`���׭<'R(�������CVW��T����CJ��PEb<6|?�x�@c�a���dC����V��^Z���.�7��L�d��Z��g!H�5���nh�`��3<��������{XD�w72�n�B�c�� �t��3tP�R%���>��ݝ���x�!�b0���E�H��d�ժ2�߈OyD/���孳�l����ȱY�J$3<.�#=lR�[��<�)�����U�N�,���65E�[�1�!*�MTx�0�R�zAhO;M�zMS���Mꜙ�Z���A���E��9a%��"0��0*�e�+�OB4*�<��������i� �Q��ې�aV���٨;
�\x���4�ٌ'�/��{�W3)j��\��s4�d��9o�H8f ��n�4��Ɛ���E6��RTd�z`�ƵJ��f�pF��0R1:��o.*S���ւ�4����rU�˽\꧳v� H^�e~��p���K��]��UY�%9��#�<�c���a���̽���*`����g�_����Q��91g�1�\��5�$�^�]��?ޥ�>.���2���q�-�4��<��A�Lx�sN���u�9D� vn�;��̃�B-;ڠ�F�#��\RM>#,<#�{�5�?�MC�ȋb�eW�`Q���㑑E����4l)Zu#I!&�Q����q�g§x�G%�\���bPV���1Z��>��I��UpsN�\Y�
8��g,^UI�W���ߩ����&�A��`b�U�J���>8Ņ�g��ھ�c��QZ�iZӠ*���0��̥�Q��sc���c�.���=�!��[.ǝ��yV���`��R��U���y��<g��{�F���}�h�n\M�*���q��_�����WZ����<�v�yҫu��-�Q`1Ñ��դ�S��P` $�fS��
����:�)���a��hC�:&�0��.,�o���Z!��0�0�W�މ���U.G�Am"���>zѻ?�To�?���%������5������bpc
"�)����*���O�6�f4%D`���oC?3�R���Ӂ	�!J-ɑ$��z�&��$���>�M���v��bi���%�י�ۜÐZ|��G'-K�ɋPR\^wauƞ�ߐ�{x����_����)�u%#�s����Py��a9�{W	nq�iT9�Ӽ�}��chx�Q�s{��8�J��� y�G�NP�'c$xԗ�<�Z������K?�]�E�����D�AY�s��X|�B����K��_⾫
̎�+��ؤ]԰�뷦Ja�\(����*�#^z�J�Z�.L�̛�%����N���Wخ��X�^�(���X�,��I��.����*��i������ў< _��]�K��	����,��%g3�����C���}��c�bOq�=� Q�=�߇p�<x"�'؆We����b�1e���v	�_�o�v��+�e�n�r�epD�j��ۢ����!O�,�?JC���.��X����+/�\���X�������>!�a5˿��	,�3���J����gE���IՎ����XC\ML^�]l,cL�K�6ɭ$�q�}��bs����h.JD���OJ�IG��J����P����4.#t���S����P�s�MGx�e��D&l.��c3>h����YO۔;4�i�(��oZ�)�ٳ����q\�B�4�Q�����Bvo�]v�9!��%�ߚ�,�,8��;���m$^�����U����1oǱ4�:�ο��(�E�-���t�5�Xz����`����$[]e��Y�c�{l�.Ӫ��4]j���Q����O�؎0� �`�VT+���t�(rF����M�����.�uhoRrex��+{�2��6R���Q�kL!a�ɜI�jBx�m�&C#�&N^�����97A�QT]t�mצ)��Vb�x[��r��ᖎ�:ވm���I����ي�<��V��x�������
�R�!��?�	���{�yb��q]sg%�A�H�*���/o�^)p�U���h̭� Ɓ�<ga�j�r�Ha�mw*Br�A�����#�7uE�L�_�+4�E�t-ˇes���-��"ه��k���n��,��D>qL>}����ӠO+�}V�
)>-�s>�����te4�mw�+x�z&��!���x~�j�Om�S诺�\��}�TIVV�r�Q��Dx/d
u�50��<u���FW�F��� sa
݁N��S�5ݪ�kz#��鄖�:�`]'�JQ�H����B;�\����0M=y���4?�4��>�{��I�MS��S���9������ƛ��s���I�%S(�H�]���.(N���y�P���8N:����ν�q"������jǻ�&pdH-���q�����W�>Ϲ��jF�����z��tYwc�^위1����%:`n���:g�6udh~���RA��S���{��-E$��q���5������C���O;���&}����}o{���s^��h�*hx��r�~�9W"ΏS6��U%�S���u�僙>�P��$Oq�po�\l�+�6�ʀ?�?����1�pG�+E8��-e �r��k�_��K���.�/��Nm�QE,n���J�޳0��z/b��%��M��T8k��������z%O�x��X���ɵ����-\�.=�pJF�Px3��S�Rj�ioiHk�w1~W��I��ǣa��lW�,*�v���*ڥ�N��M��Ѵ��wb��#��1�wu�9vWu�(���o�i������Ƴ��<�aL���đ��&��� �k�ŋ}�o��ֳ�d��ܲ��-C�c��`�L�c,tL,�ﮌ`�C��ϱs��M�@�&�q�x���� 퉕%��`Տƥ���\S�N�R�*�m�~���s$B�M���t�s�����-.<�U�t�Nkn�� ����6�+E��&�W�bN���1��s`K�g<�D+Q��	^5�!��E�K�@�xȘ3�迅�ۋ͛�)qxJ�H�C]��@�(]'wh�v�N����H��P�?e�-��Qrj�7y��zOǌ�q�-�#�s�,���S����<��m���C�����=���2�0��N��I����r{�Ґ�'e឵�Ѷ�ڷl)CXp���Zy��C���(
�C?BUfk�sa^J���6���+�ި�&���$���7��4�]��C�omʌ�&�_ӳH��(�((�d�d��9�%�RN`{|�6�ŘV1ͯ'�j�EO쑆�i�������)�5�!�4W�����G	�L�,<Ҩ�c��0f�4Z8I�=�"w�L�r�>�D�H����JS��L�m!TYGIh H���92��tc�T8ڊ�k�T'E�w~
����xۍ&�.M�͑�-B��-��>5A�A��]FѲ����LVcf)cg&E+k{ɉ#����a��-A9�v��GnX¬.U�Wi/�_�s�#�~Y����D�8�fv��<n��\�dkJI
쮄u��Q�O);m�V[�wӯ�N�C�Q��DT�����"�e> B���XL����k��VM�$,�y���?��ۉ�9���Բ�]p>*)�X�c�ZP����;U��8A34��jf���h��Sf���<�F2��D�L�f���$3�Ҏ�� �2�`�^�S�E�zHQ���!���zu%�E��E
c������c���a���R�v9Mynφ�lc����+����.0���ޣ^O�!�Ě�,n��]�w��"�!`C ��6Ё[� �N��Cd�Ι����H��@_��^B�b ���XJ��'.�I��{�}�*�p���qno��ciQ��YVO�;X 0�02�(cܚ(�LA�bM��vx��!�ҩ�N�+�ğ�wJQ�\�
�F��p�ƃ����ƈ�u�i*��<ct��""�8!�va]{y�YuW�>M�FXS07'?��!�W��w�D�OA���:,�x�	>g��0sq'ݙ2�ax����H&�ޭ+*�*�FB.N:q�jC��}s!���J���Q,�?ERF��"�����x��z 06��U"��9r	1gm4ovQX�}���ǜ"��=�K�S���Ӛ\�m���_��rTR�)�
�1w�����>�{qݻ�8s�#Ā�Ԃ'r,��S��ں��(A��C�W3��x.$#IĎBA����UEh��
��k���l�G��Gې�߬�5��1[��6�.��]��.�]��-#Z���"��А�dH1p��C�%=?T�DX��hCQ��M�ݴ�0Ȅd��W��E�3�à�$(���;���w̾��3�y�g/Q]t��]������2˸������e78�]܍+���������V�g鉎F`6ؙ�R��O�����
���a2*��f�9:��t����j%��+}W�����l�Jxh}Ty��	�˘��)��-�h�G�C�����)��Հ�_&='$-og�G��	R�tZ$A��1ۘ5�ԇ`��$7���Աm�eU��S��1k���.�N!�܍y��%�;��c(��Qv9�F�l������^ZES�!{��(ヾHF�I��El�۶�p�3lP������lG�S��W*��<����%���L9���=J�����؟�'��#�Y;��r>.+55j@⊘k���	}�6�Բ�G.4J�5!�9u���U��X��}�~.8�1H��1���7��j��Q&����f�������b(�ĂG�`��q	��A���$ٷ���T�<��z�y���D�>t�:5F�A��Zp�.���7�~�ԛ	�Z�����ڻ68�dkN
�y.+��&ZY��-������&T���m\W<���RL�6x}���Y}#f���K�wT��7���snr�!ƞO��-,�n+��������s]����fڎu]	I��]L噊�q>�+��w���&�O�9� {)�Der�*n9�\y��'�eG���#�A����Vx}�ы����H���ܠo���͐G?i��gvy�MO��Hs��/C�����*��Sb󒶩� ĭC"�d�K������͌�	7���b+�/�;���b�_T��`pAm�駟����Ɉ����[k��1]6��@7��_�.Ag4WYc;��V���YI�ψ� s&�A��=������6��f�U� Rrɕ�Im"������k�����cri�@���c/�	�I�[۵Z����ҩ���v��`��v"���1�H�\i(5�B��Zє_��H�p`2�c�%y�Mϛ��x'��(t�j�kgWr��]�ͺoU7ѠEuap�՜�ؐ�ĢE�:��N5�E��sS�4qLMS����uZعWV�G3��6�Km��Ԅz|5��89y��Eg��,�.3\J\����>f�i<\���
";3�R�'�����1O���M�I]��d�8�56w�F�DjVD;�&YR�j՜J�����]�����c�x��G�#�@��jm[�0��5-V,���aC�d�\��	g��ɛ����E����Κ�N������]E�_5�ϭ蜾�h���/<�"Ag]AS�ܒ��i;����񯺎5y���n����q� ��C���.x�ێ�Aл�������d��ذ'�D�55�/ш��=��ۈk ��������Ń�ڵ-�xƸ�q�F�q�Š�)p?	�����H���D�U�d����7V�a%���X��~��#�߯Cp��J�����3A�����a������k!(a.e҄6�����U���ݠ#>��4
�a���x�nn\����|�}��e�Z՜r"m�7<0Y���>���a��2-J���]=Y�@�@�t�r�l\������Tĵ�%1Ŧ�W�K��=���n�E=�sn�33kL�����C_3U���f��s$��l�8�!^2�ĸ�a[�E�5k؞�&w� m�1�]n�"�2��Yb>�ʯA����!�\ѩ���]Ń"�i�N��N���x�Ϟ�v�G��+��kƔT��x` �����Aw���lXQ�ʒON�[���җ,F�&2C���τ�,	g"Ivg�t}���>�� ���vI��dx~��I)e}�r~�
�N5�h���<���R-�k���FX]�*{�����/�B��xٓG/��0E�ᄽ-�7�bFQ�[a�ؐ�������!w_mKF�<H"��7@�ݶ��Q2����������	����ڥ�%Qg$�.ޣ����\��������� ̩qױ+��^���><`c���~P���xF8d������1zw�o�&�Q�1)x�NܳKE%qe-�92���W9�"w"f�K�$��M�'^c����p��v$��Xc<f�k���6�H�vc(�[ fb��.Z9CC0{r?�g�k]k�+�j��N����L�gf	=�i%��0��.�9a�-�c��~�1[���o�C�6"�E	$$Z����ÑaC�n��z�l��T��\IԹIW٭��]�^@c�O&��x˲˔�̟𨰁��[���6yq�D[ʘKJ��c�X-I���a�-~5�OQ�}���8Gd//�>�(]\�!���h$�})�zr�^�>�FuCW���"�Ι�秫R֡8t���<)��H����5�	��/�Ƣ�PJI�3����Yb3'#DV=��J���Dω	��<���#`���x�!�3n�ίg��iL�x?�`�E%��	�q<�E.w�+�c�s��3�0�L:�e�~#�~^�!gx
������H_Ef�FS��&��V��`��jYG�F+� y���S'{���K�����1n�}1�p��T8���(q-�f��]{%���F��K$�앚cZ�%23V� jP9�n�##��Umflw�ƙ��N�`�'��g�V?Ex���髏9ciM����:g�bfE��26�%������f������5��Emrn�>X�N��6�5�W�켟�����Rp����}��榺����B�zƃ�	��VDo�K�[���n��Kf�+~���W�����X����c�x���y����1�6D9m�N�8��g���&O�K�g��&���}`���NA��=c��������H@A�xp���C]�>�C;����8WX��fM���B��w��n�*��� ��oB�%�=�u������X.+� H�f��Pk�!���~/���b���!O�9��	:a嚣}�U�6�@��C����2JB���<wBQ]��y��w[�:I�p����lQ��F��KKn�v$=)���ׂq�8��$G{�Ӝ�T�-ojF���������&��6t�+�S$�Y�����(��Xx��K��jK�?������9xN�G�*��q*��BR���&���5�����H�}Q�PL���ڐ������n�V��S_0'�R1������l	&S�d�Px��`�Quò!����U�h	��Dٻ')���ل7�C������^����Ի��g$fOS�"�>�hbh։�9�D�¹K��;�j��F3g�YN���]^�2������uv�����d���)�9�ǁ^cD%A�P�K�%5Xӵ���YGey|�D�#�p����m���H��a�=^�sj��T���̖"ژ;y�h�����:0�&��C�ҜY�*Rj��S�>o�K�������۪��gET�����X#�Z��V��U�_M�������\9B�H�1h^M�rv��&*�v����+���>�k�u$}�/����ӥ��l��S������� ��[q]`�Aߪ˽sR�+��rKDX^��}n\+K��i��~)ü��Y�IB0�!��:qh����-Cߝ;"��g�	�=ɶ�H��5Ì}����N��V���9��0�]���n�j#����$]�X���\D�E��<�x.?���+�6��A0�7��OgC'aܾ�*@���x�7o�r� *��,mă�XM�JR-X�Dr,��Pܙ��Sag�0��e�V9�M� O���iO��dvAln+D$L8�S�n���7�~�Gc{�Cqs��8�1����H|hvƽ�8�C�ŷ������H�f�3�h������~FU+���׼Y�sl��O�{�H�Z��<�ې���p�E�xP.a�*;T���j�f�-|����p\SzJ��#�t��Bg ��k��8��J�[%��}��-Q���6�.wP�XQ�7���bH���1��M��%�"톈j��~M�p\]��4���L���hx<�`wr4���*�>�/���}֯%}w��ژ����@��y��l2%*B�|�eeꨋ��2E�O�|�u���9�}����&y���$m�%"��+P�re��̞&B]ݤ&9	bH��%�W���I�,	��U"�U޸d�j���M#TQ\ͷ��b&����v&)g��Ʀn��<��s(��`�3��Ha
�!k���)��U�5a��ish��,T���nB�x^󜮼Br������(=T)��0pq	�T��>ۖ���R<���7��O��*2��H �wVfB'(;T�jRM��XƗI<Ѷ�`a��)������;ww7���S�=��8�J's��:pe��HV�P����KV�z���J �kC�(�!�4孉r'���F��v�2�&0w�+\�s�)UWT����!$����N���M��^_D���K�r�g��!h��z��)�zI�����]����[�o���㻹a�A6n�.��H��{��1��������"��U5�<8q�{���1�Z�#4܊������w+$n�]!�w�C��V�!(t-ܻ�+\��)b�2,��y�İ^�� �EQVG���6㐙>��U�L�`4I�C	�mӔ>rw�B�LPŐ�,�ۖ�hO��"ߓ�/f��}`����y����yr�>�36������Ԇm���G�?�o�"��¯��Ǽ��C��vT�VA�W�>C\m+%|���h�7C�%�`�=��FmP|�y,d�CZ5]u�]�C���%��V�06�HN�{����͖������z��WB�(:�ΰs��T�����!�]�ެg{8ກ�tY{�1��x���~��ni0ב�f���O'��Ԙ�[W�6�%
��ę�h�<����%��5��E��-a/�`r�7'�,�}E�J)(]�\��D�e{�T"�(�T�jDdng���Md�o�K��ό�@\�sV�n0��ۚXz{	'�����5�4l�37�:B���^)�Yk�/�����I)y�hu���̮����jr�I��B��d1#�$t�t��q�;Q�d��|u�x��P*�/�C�L�mԕsw%���%,1xOؠW�pN�Ñ�ܱ��kNr�;��7�R��S/�Cl0/�^�k��[u#M�N1V�r��1�"fS#��0�?l���Tb�fo��Ʉ�%`����7V��:C5��Mz,�m�]W�S�#D���}{�?=E�M��I�+�7��]�v�9!�ǜ�8��a, +��f�jbc���P���4O����q�)7S`ԋ�r����b��2uY�p�&�t�M̑d��~�aĿ�!]��]tW8`�X�R
�������0�>��h�4 �Nv����<n�=����mx���KT�T��m�zl�\���W�M������Y���q�;EC�/f���x<0G\>�Vα�9���Q��$e�.ӛ����l��f�-C��ک������9l� 3X#�T%�W��z-fu�2���������4�6 ��P��I���������8��8�>v��>ǍxZ<�6��P�aHD|������յS�$(���å��R8��	����E����R�a��zHw'a��A͸<�@��͆�Aoj,�)L:�ډ�P�	���#�����o7�Øܓ����fW��7�M�,X.�l�\�Ŧ}w�93	9�P�Hno@���)&.�G�)p�.2���w�T�j];b�nZ&��2�諒��]�ʫ����-�0�l�r��.����t���@���K������5؟�չO���H2"<��|�jJ��i�$�x��;qbI]XsS-$���훷�j@��
CJ���c��mN��������Q�-����j�����Ԥ�%��Nz�f$����_��-�S�7b':sk�H��#5��v�Ϙ�b�L��zM�_nC�"�#C^!H�x�!0فg�Z)j�"�ms����yNn�Ҷ
�aH��g�q����̌��!3��� U�deE��_�u_㡳�|��/���!\З�K����l�r'`$����^<!l!%�G��
��/�!/6y�&�G�ʈ�NIv�o�h�9L�6�+��i6�H�r�u���B#�	�j঺��ۻZ�N�������Z�QgsK���E�4�:�xOH �,(ã��%����ڶ���6�x���88y˄��v�LB{�Wl��8���ڸ�Ɏ�\@Q\���%��:o�C%�p�ʺ#tfk��Õ�;��pC5Z�����D��;���6,�j���?�tSDT�m�>"�p���v�/2�(?V��h{�CUrd/��c$T���n�4����v�>Z���Ŏ�Z[���li�1�E�0@�C��0�b�,�b�Đw�r;7��(ڿ�������A�2t3Ny�?�K�]@s�>8�a�nK�*ZS��)g͕�*��5Dk���z�Q��d]�	p��*��1:����ʭ���8���=7��u������J�#��ԔJ��c��iﺴk��dNaf
���!���<D�0��=�7���;���V�Wig��2U��9H�[�r�+�RC]��_sQ�0n�%�r)d�����k�ׁcm�˅�W�h�����n��b��?�����)�=S~����m�/!w����K/o�to����T��K�
�.��|F��������}�.�+1+��M�To#���J,(��]"���ϼwmNr�59�B�ɭ��jD(0����e,�jV0�����+;v�c�YBN1eڊ��P�W��\�"TBC��������@�Æ�^�yI�0z*�����͎E�{��àc>L���ެKrs�̉��3��1��RlL��Օ=M{�b�
���2�R�K�V���!�D�%A��p8�y��T�����K�z�\#���n/�T��g�ț�߷U.��rn_�Sj.Y}�y�*�^�MW�9Z>t�����~��lSR��PW��0\O�Su���{�1dC�e�|iy;=- �0.�Z;Ĵ� ��u��r
N|�S6���esά {�;N�m6��@�>�d6�颤U^�1*,��lc��<�*�QdZ]RGjɬn�۝zr�Ӑ���\#��Ř��x���U�,���e-ry��L?]�Ncľ5˸���lu'g������zu��`���z��҈�_��62�T���2޷�/���������8E�\S��s_&S�Q��gx�cb�������!<�B��|����g%�#Gt��\ "�$~$�����|3��%�&��я<ɿ��s�I��,�#�!uG�1".i���]�w{��	�s����z���n2}�1�.��)Fw]�������K�ٍ2���M�,�!E1Fx���͜rI�;ǣ^�`���p[�2�`U�wj�8_R;?x0��XG�S��Wt+p�ϼW�d2�������霍mz��lG�lb1��=�~��U����}@���Mh�9'������Be��#��;ע&A➛���
�%$�p�L/��V��'�����x+n���Ԏ��SZiW��s�Xvu5QFX�q~�
�{�X���P`�W�7��v	�N��m4�p�/��9���x=Rzp1�ct��VJ��e�����ĕ�*a��<�����y���W	7���4�QE��6��N˸��.s|e0T5��nk����=���P��9G��[>�nJ-�Z�9���ޔ�8�t� L����y���ٚ�:�
/W���%��h1��@��1���T��I���^�z��k��[OL2��`_��=�3ÀJ�f��%��
����=��n�n�#Y���XK�K9��+��x�/��
�5�I@�mЋ��rDF�!�c�K�� :���ec�e1GO��:ڲz��Y9��+UkS��p����YU��"�UG��ҝ���::j�'��[M���4rs�%1����Ѹ��<_������3�$�zcn�����e�t�v�N�c�����}�u�M̹��g�Đ[���%lq�{�j�p\J3�h�ǰl���!3�c?������q@����m���Iҍ�!��L���U�,��m��D�������e2=�9�X�h� ���A���F�7���ݤW���:����@��y� h!�;��Z�F�u�dL�,�x���wm<�ɖ_��+�t��*�/�1ƔKy�X����}�w�M����O���۸�{�ܓ4��+�!U��zA�nu5����+�fl1b�Ô>}�ϡW�`k�@.��	��"qq?�-�������?���I�����=���ś<��#�H�lE7О`�h<}�~��46����zا�4
3��0I���7o���}������xhK�Ԏsǁ�����a|���F����������e��::W���B��K�Q�]�y���x�b��uj�6�n���u�ڂgN�D}໊Xq���=+������+m��,~�hP\��p�y��
�sl�EeQ�e½�;#��s	ӝHz�;G�n�Ve�W�J� f�fD�y�W�ȉ�d�z�J����[�|X������m}�o
p�)J��a�0)��9{/������m��n�]|�g�0��'�jҕ��V��ZR}�8�9��4��&��dVWO$������{�����;,��͊���c��h�a������&�k�L��vd"M�2�!ii4�(" ft�����;�L��k�h	!�
�Yh}f�,Y;c��
��3o���6�Qw��y��MX�Ȩ#�D:σ�t�E�^�x
�������9��O˩)�����Bgv�2�,����znsd)|���!+�K0f1>���!��ǟ�O��-���i�s����ç�p<-��,�ܔv�l�6��|��m����Ć��z�����o��r�S԰ҊpEd�œE<%�%�߿��OB`4�T::��z�VT�����K	p�� :T
̐D���I��t<��v�s�T\E�s��"�8V�I;�1i�>J�G:�=H�_�C)�&W�1a�P:8ݝ�/���E��7�0��\���S����]8���l9�E6�஻���q��Y?�kW�Y><L?EWhgeI]80^i�P8�-���)X �#ue����G:��u��u�L$Q�4��g�"הJ�8\�}�oA���9bR�B�*�T����}����v(&ҧ�md�&e�������<��wT�?g�-���i,����~ym�s��u��D��=����j�/����bDOT臤�n1�/_�`����B�?��K-��H��mt���ky	Lh�VzJ�
^���O�u�C���%d=�I"̫U�(��T� u'=�a�+��ό ^����+&A�m�X.�&y�����%�~w/�J�|nX��͔���l,�N�<\���}����2�(���u���P�m�J��p��(�Uŏ�~Z6�?ӧ������x!	�~>�I��C�0�0�^�y�~���?���`����������/���+F��w�|�FБ�&�	|��o�r�)?3鈱��G
���	M�9����	�w�r�j܏�Ζ9���~0��A�h,�f0��{%l�k�ޤ�v͹��i�"�9-�U:�Q��TրP⩋�Et>P[�
�{��Ex��i�ᢡ����\�l�Io�o��@ö�ŋX*L���336[��"��*�Ԩ�0QA��$�S^���$��.k��XX&�~A����k��~�;��o>��X�,��ɕm?���~E��ؓB9�e�<@X�x�ъC8�6cdH������V�Cb��g�ڹ�|2QFMё�	O�G�[���=�6����D��~ܬp��@|��Q���|�	ju����냐�LJ���K7�;�����f;y��g�q���0[8G�\Q�V�޾���U�7RJu�@�X�?+05����g�c83tSc�đ ��ɠ)�#���7�1CV���XN1����WA�W�!�r�"��	���7��X��	����Z��_����_����Y�.��6�1f˛����%0L/pm*�6^5����.F��׸`�Y#������74h�3G.�z��Ⰶ�+���P%�po(2-ĵ	�#��݄�ng�:(���ؚ�B�t���pQ��{�� ���I���o�NT�#n6��e.����3Mp����IT�I�a�s^+9ǒ܏J�����t��F4��Pj?{�%2�}��k��=
��Ե��V[y���hq6P�,���*5��y��1@$FT�'�[��jڐ��fK��^^�ƀ9�J�hC����\�<�a��}�����r�G�g�>D���g��i���2�{������d�����|�(�ؕ�N�(X�R��ǳ{�br�0�O^�T�*:��R���7�z�ԕD�h8�R�K�jwV�U��Z.�:���A�P�[4h�y�]I�9JW��e� &�=Q��cU�H�i�b�/�X._���^�,�����o��.}��w4b�Nܫ����￥�������8f��fk���������՝t�2J�W���*�]E�w�;`Pً,�7�s�{�����׋ф�y"?:�:O1�$�2j�j�'*B׼m�_s���qB5�ؤ�2+�9��6ox�7J:͜�Y��,��Ê�������Ms�(������in�ۼ�Ԙ/��/�|1��!�S��{S��`�h^.�|��[s�E�%��ls�^���=�P�����aH��u��4�~���!,��H��i/���M�+�ΉOy�~]������1��`���vhkB�1�#�i�1�	ə�)0��*W�ecó �/߁���k������)H1Р �A>P��z��XT�q�����d�Ɓ��\��-f]״[�ߴ%�Q��8���� ��7K��-ѓ�b��n���!x�nG�Rי�E��p*���x�G���w` ��ɤnJ0.��Kg��Hs��l��jX���au9�o��7G� �X-F��6(D	�?��<�g���_	�������^�����O	���[15L��:�31fC��jh'�d�)T�@�#�̞ߨ�c�j �6�D�_����s	����@��M�{+�{�#�d���+�fe��]���˜���]��Zs}���<�9��������n��=+!:DiÍ~�2Ow�d^c�g����y��HM��X8p���}�^�i��0�)��.'p�y�G�ϳ~�ިy'�/��־�H�U�)��N�Ōa����
Ƭr�c�ջ�PF��-��V�C�`C!t�6w�Ӡ$E�c�l2N��Jd�=�8�n{���&��D�m�i"�ާ��^;�%$[Srm��C�:�<��?�w��C*dE���h<Wa����n/V���G�o0�K�Z�ω�ϡ���Q�)1�<5�,��s�H�.���j;�ˢG8E���ZQ ;��@B<I�j50Y�ٔ���QPTc��ǜ�x?��4���ᔩtSH2�4y��!æ�ӏ?��o���8o@X�����@O�UA�h�E�c5�����-���jEDG��D��q��[<�r#bBF��(1�x���_hȥ�����9��b]E;�L��f�LC�j���?�9���ܯe��q�����A{E��"��W�ywںUۿ��m������=�Й���%��Ys��a��:ڑ�h�3��A1���ʓ4�2��/�����L	}Ơ�cP~N�nU���A���ĩz�x�]��J�ꎜ>��&�S��2�0{��C�H|t���� >c<EU6MrC0�ש�p5/�~o��؊��^D���w�ty 2w��ar>�i�,*�Zww|l(�L�s��a1�x��t�B&��I���d�>5e���;���l'��D�����e��MT�zEX7<g,Vp���Ar��V#�hEb5�6�0l*�4Q�|X��6l<��rb�C3�>,Mxw�=h'��~5rj�4=�(��#�2]Ox�?��st�L�F���Q���>���kF
������M������e<1_F�U��h]�1hEl���镼Ub:v��w�r������x̠�=U�Z�$�Tb���+�������NZ�AA�w�1ccAD"1Ϊ����0��_Rƞ!�)���|F�����{�'���D�Z��$��	K�'Ut�OWx��H`_��T�х�<�bD��m*R�*��q����)�o|�&���|��>����hyvaH]Q!���!Mj߻5|[�9n�T��  �v�]h�Ӝ��"4ڸ�{�	�{8 ߐ�ƚ^{s�-I�������0��k!��E{�d�G	�T�=�|��ux�=��x�B$z9����/���\�&w�?O��>����!�Cq�U@�V0eO����\�<�.g7��U!ԘG��
�`:DM8&�&o�wR�xY�jHW���K]�\�q�5��7�]�܆"3(X6�%��8�i c�l��v��׺׸V<r"2��8d��g�}�2�y�6}����}g��0L�_d����{�ws�������y�d�}��)�����Qe7D�K�V-Ԁ��DT&F#���o�����G�޽��>%ť���Ue߫Wo��m⸂�J��1�Y���æa�
y��@�*�C��nal���u`�q�9�L�N�*��O���&�
L��H��
�:����$�Wc�.P��7_x�^+�1,�)1�⸺i.t6:)YP|L�Y,-�k�(/g����v�7!�ڀe�6���R�����-B]��<K�g:gж�@��3i��N���6↍<R-��H'y��)��q�D��a�&(�kVBϳUh�rN{'}XL\5��ۧ}��1�v��=!D�
���?|\<�O�V�`(|�Lh�}x`7NH�a3px��pߝ)g�ex�:ҡ���9���Iʤ8.��H'4*d�.^S��������X���O�,��"%8nr^���0gN���U���S9.h-�ˈq�kK{%ЦHxΐJR��G�뒾����J!
�kÆ���q:[U��3�ىs������sot�ϟ�`��J��e�6o�8��U_{z���s����I��p$v�����ת���H ^hϬ�(K�7�4��+p���cF��M�Q��F��@�[޽^�9�*!��r��j����_獎%���i��a!�GCW5�I��y"��UC�*W��T��M9R!{`񜛱4 ��Yzh�����9U3Xd�
L���HSع�wϟ)º��c�u����R����Ӌ��R����X�m��\r&�]$�����h�4��U
ÊQ�*à���}N
�抩��-=�M�W�QGޯ�
+\q��ߗ���Ű������V��S��٪_g>���x<e>��J]�e��)q�Pk�����ד	!y�
��Á�		���;��� �#<h^Έ+thtp��ܣɚ�� �Km����~�*	�a�~�fy��,��RʃJF�,�՘��^+����p� ϡu���	��D�����ԃ��|����n��5�{ 0�*E�d�T�-��+V.�����t�/��̐~���<�:T���0���LnaX<\�\��D"���=�3x��k��H�k-$*��14q�3�s����͡�:��X���ղQmyk�j���p� 6�M��4���{��HD�ϔ$j�,k!dv��~�1ob��9c�8wќ��?e�Z#5;>��R�W�+�!a�d#��(�cR��vJ��kH�p���$�ֶ��7hO�L�YS.r,C�^@=냃{�{��gā\���Y���\�R䀹�md��zC�*Φw�3�R��p�$�a����r��T[��#����P���}�Zv�4�U�}�}�ʐ�x��"�F�E5C�D�w�MMk�������|�>Y�<�.!_hal���QыtZ��� `����C�h�h-N} e�����Ta�k0ygO��?/c�*��/"4��Q�"�c�)ƃ����^=zRr��^sI��f�1�!�r��s��T�P�e�C�%�Mt�-e�H�`LXu�d�}�~Hj�	�Q�f@A�r���4�#BoF$��� �똏�By,s�&6{lr���?}�!}|���ɱ�mw] �x���V�/��hvK�&s>�X�$`䍧��R�L9�Q"G9H�/ב�d�<燊��t��[�Ug
X���׻*@{��T�h<�q����X��B�չ�*�d���'GƵ!��Sd,����\g��3٘6
)Mՙ��h�dI��}���$���Y55᧔����r%�$�$�N��$,�H�X�͜�}�6)�[¢�/�M�v
!;�=ڻ�F����lı����D(#HC:�#qq�'JoT��F4�YLSeH�\Dzn�x��@o��v�2��٨�$%%k`̇h�P�3���;��O�5��F�ڧ?P��tgZ����L.��Q�=T��n'�Mn^.�EY΁qN�W��?0��&	pjQ��Ǖ�]L
�l��cx_$��9��5�����͹	�=Rx��,��T� _��c�ґ~�1g�?}��͎b�Q�&d���3�8.�����R�o�~C�:0B#5i�u<-ǖG�t���%.h��F�$lfxR�g^�M5��6���n]^�:��lE`�xЈ�8����e�=ۮ�����l$OM�������	hm�q]���)����>�?F0P�
-j/O{�ִ��4=TQ�;)sqL���S�m_پ��h�ƪIW;�W����w¼&�_ь�9�p殄5���B�R�a޵���2�Xp��|c�Τ��Т����hʓ�������v�����@X�(��g�v/u�u��n�';�dd�Q�V��h�"��c�F���*�qTP��m�"E
|�Z��g���'��mt>�՜ͯ���)ZN����t��8&�]"�p,L�t��;BR�����}�޲jG�4�V��iʊ,ƠD^����Us�PN^Pm!{�Ә��%5.ᥱ\���3u5;�J�O��B����	Z��q<ED#e�5�2B���u�#7l��D��l��������2�q�ߜ"Id��ןKu)s7E��e�織x���+p��]]!���Ű����'}�h���a�M%�=��S�/�Y��Ҕ���M&W3V҉�3{�M)jP��AFxtr�>�au�@�f`��K�Ũ�_�7_��&�\�����dIm�+u����Y�_�������x�o�ض9A2��%)�&u <CG4��nEޗ���P���3S6��E�z��`,�������EB���ˇz,���t7[a����9 �dq�ݻ?*���� �,}E݁]rU�b�p_@O��MD=���ˤ���l񻻹ͤ{֛cG�B�96�c4�c��[*�x"�ӂzfQ�)��%�I�����K���V���4��wO2`�qbROك�!Z�J�:ȺCl�Ǝ����R�tΟoA�j��S6kCT;b�(tn������Im�72���[Sr�R�M���bq��v�GJЍ�C��3�4�I7A@?e);��VK�X�8^�!�qkW٘�>E�!�Oz: }�O�(qNY��h��n����a
(`H�=OQ����
����J����"<�ip�����RT�5$��"����el xnO�h�UaiS^<���D�%�m�f��܍�i��$�X��b�����y!�dJ��uŒ4��ޕ��˧�i�̘r~�z��h��4�2a��i=�bb���%vqV��0�O�!A�;��?/5y""��E�rQ�SV��y��(�iG��X�d�������\�rmOO��}�A��J��F����=�-�ت^(�q	C�9}:]h����Z���b��Z\Ӭ�ވ�K��u�Y�]���SS�(�[�?{}6�
�ֹ=2��1<3d��:c����Ĭ�J�����U߿�ԭ��=!'u!P햛�SH�ɻR?��X۫��.͙�P��!]�Zg�3�I�;���aՓo�:x���TȞ(������Y߻�B�i�"C�ce�4�4�c`�dy,� �p�$�`Y��>xYC��b⓰�%W��[����c�춱R���^�q�Ȝ%B#U�UD�����5���#,������ �?���9���r�-�QѨ�n�vyn�*���<�s�����^�:��ht�I�3�ڔ%�q�u�L�͍Z�Q����5@����<���fj�0��b�w}eC����X�Da�<�ݪ���-$D�9��5�z��lmC�JU:��&o���3MA��8S'"Q�w�t�`���a���ĉ~�E;zz�G�󪖖��&x'X��ʹܵ�l�֑pi#��%�`X�7�w�{Qկ7�z�=�"�#x�kqt	���<.A7��ا�k�A�Q��m��:%���7?�qs�1�T����<M`��d$��,3�c&%n���0oTQY}K�c��ğdHy��/��ʨ}uT���<Nt/}���!��K(�b9P��U���C�Z���AlH|b񁆆369�s��o޾Y����#�-<I��eLnwڠ]Y'q��3�PfIY�p�P����Hś��Rجq��c��� �#�6hv�1��U�m\I���Κ^�pu�Ӝ�>,����X�3�{�!�/TΆC��zf�M4E4<DGi��@&���W)_��3e��<�>I;��u��T�l�Ӟ�7D|'�uL��[�QK`喛�|\��钡&z�mg����*su�������C}󟔈�p�J��{k�D�Z�up�t2x�R�ìE�$�K2W�]BJxiY85�C�n'��Oו72�4�:�BY�^��i�-�5�� ?^�?��?s�#Y��S��9���ܭT4����]O��d��ޓeOjL��Л�(���ٛvG�$Ib�G 򨫻w摻��������73�]]����pw�\f����Yb6�	 w35UQQ�b��F� JVȔ�j[��*�Rj7v��[<��=��x;s��'~9YP������f�Bֆ��B�8Nfq�ee-\ے-���BkiE:�JD4�p��P
��̵m�%'�tД<��ZZu]JM�!� ��X>W��U��ͫ�*w���*�#+_|�܃V1]��\$�#ۗR�)t5D��le�,�=a���l=z �T��|�p_���F�Cm����]��$%�T;i2ֆ7fZm�}IVB5Xo�rl�ڔG�N�l��!���~���ӣ`=����g�p�p������s`ct�O՜r��2�u��η��c���se�����*���k�)��GBײO�jg��a�.w�v��s�-�Yꆦ�ͱ-�4<��lޜL.᯶2` �`�;�����cv�N�W%$+�Wl��Ģ��kB���ܪ}��T��AEguSI�$
*��ԩڻ$g�ͩ�T3����ИHXf9��!q�+�M0r�^^*�<^I�R�(�Pn2ۍ#|o���$	�	^�!e��0�P��f�; ��b�� N�x�w�q�U�Jj?S�/o�'�*8�Pw��m�Xa����$����$����i�M-"��pM^_�\����gW��|��8�.kÄ�!�}n�����T��^ȭv)]�g�acj�:WCa��:s��C8�!^��?~���}zW��L�T9J� ���y�6�Mn�b�]�ԖvZ�]/	
�<a�//��f�2�3��x0��a�@KNj����x���R�ʠ���7ۖ@IL�� ���߮y�q5���}�(;� _��dZ��.�֤p���_V���k��a����4���R-���e�����`�B�P�9%h5/R������t'`�()�u�ϕD��b�z͂*; ����
��أ���*�w�C�$���"Bt���gss�I�����>7%�A�F׿�Hqf�]���կVw��Q�L]�$+�63�[ن�hTu]���C� t�F� r/��z�y/��:2Ql�w^�g7���.�7HF�*���f�6���Bޘ5��Ha���kWtM���J�
N9Z�J���C�h�Z���K\-�Ji� �2�~�L&Ͱ�f����m���a5#�ԬF]�c՝=O��zY#�'O�2#�k�R�VA4���*�lq ��5;	��X�{�bU�o}������q<�� |����ӱ��R�h�R(x�������"�˻�qO?|��ғ�ܿs�� *3,&c��osBc�L�iC��)��Wր�3����A�aZ(R��E��u��j��9�tew�c}=<�<�t?����]
�.�7V@�H��˄e��v�=�n��Q�	��Rs����_C}���䲰W,��ڼq6g}��\&� e�Ud3�����jF/̀H��l�٩�k8&��J���s�]P����d �2>
F���ke���-�$68�U�ЦؤZ9��������9��,k���.*�����kp��<q(�l"�dTqmSb���Y�\��AY���̓`�����&�{.���-�ͪg�|����ԎF��\A/A4�^>'U�X�f���-�]�י}�����x�FZv���մ�(�5�{��+Gi�R51�qʹ9��9���� �
�����P����yM �]�c�������o�e���5ʲ�&W-�����$cػ��JL��Z�j�6��>�QT�)U�M!,\��p�2����_�ıyD���϶�#���	ߊ/ueO�W ]��Tȥo�誠GA \��7����vo�5�����Um	\�NemJ� ���_�=���|��-k	�b�����]�<W���&誹��?3s9����H�N9�mW���.c�C�楖�����F(����'ˌs�jQ�RD�r����C�k��Vg>��+�/�+��*>�uo�oiC?�϶�+�v��R)TyT������A��@�\���.��YVO�(3�N(��T�����J�=��@T�+���dY͈R��Vz��1t�1[���F����KyM��q=��V��W�T��v�Q5�K;�]%d��P����a�Mf�W� �<$�rYls�;�2���p�^G�>�N��o�fk���<]*EI��R'�8����E��P1Y�(ax�(�xY�ocC��#�wU�svCs���j���T]1�F��eׇ��;tt����(Mu�rn���s�'؉��*�&�������I�`�L?�3�
��1+M����w*��E���$D�Q��lú�4�K� �H�Qq�^�.~��2/�ґ#���ə�����X�[M�:7��n� Y6i�vn�	�efr�윳�Y�x&a�K��t���8$��PZ"C{�6>���}��]��D�yb�z#�	#Nnh_���������q*�ɲ �B�7z�	E����K���2�*��F3�
#AL_� 81k9�K�v[+���?7�N&�����a����Lt{���F�yWޫ��# FK@^�\���@:֡�L��N9$L��A�M�@��?e��`���ؑ<앵�����6\U��b�=lK��>\(i��n��)GF�'�OQ�R�Ҫk��Zs�_^5�|y�Ը�a0e�\�}.�w���A����/�#��ݽ����u�M8&��=�@j:��XY8��/�.��컈�OT��Ņ��W�����g+:����P���š��̓�V4P�Ĵ��:5���o'����U�;X�H��ݻn�O��5��| X�4M�`6�G��
`h���¢V�:m�L͞`u� !=
J�����e��N�m��=�7���eM�\*l��d2V�v������b��f&����q�jfL�<�Y%�����֧� Wfj����|;�õ���J�����?���j�{Rr�Y>��ù�0F ڊ^�,e�wQn�W8D�;75<>��_�x��vM)%$`e����Lg���|��#�k�=(�\�B�l\M��q�	W����ў��K�y�u�o��v�VX!YQ���:��ܦZ�����d��D��#�����iZ�}�Ɵ�ftv���-q��ȡ���o�[�c�YU��g�u��3~:I�>f�i��������$x�Y+�]�kD���_K��뮊J6_ת�a�K��2�J������+^�JN��xjKPJ5����oƃ)�q�)f�}���V�����?f�-��+C�@+��!�e3p�7�M{3��R*��њ�^�i��*�^1�t�͒yk��<1AOB7�)3wT�Ѱ�N]P�{�mr�e�Hq�^R�������O���X�ݓ4��l�4ͳʙ���`>�Ue6KE-X�"k{��H��W
�h�f2k`�AY2�C�����׻�ֻ+�:�T�D��z907���V��~o�~~wh#v\Ȫ�'7c�:�H,���ȱ]��TBm��@}:ߠH�x�un��Ɋ��6YSi荄�$��xr����܍�X��\"����3�G�ܥ�|7>gLUi��x�v�Б����ŪW������p~?o3,%0Ԛ,��gM�<ص@6�[ �C� �7��1`~�~G�Jg�	X�\��N���Vԙ�Ǒ�Zګ
��"�:�!�62��6�����T �����YdQr!W�s�	����E�S���;������z-���+����{��J��w�S��ѕݪ���[%JJ�5�n-����g���k��]J�)����ͬosm�EzHM7����$VGm_�-�$�T��n/<P�\��XXE(��������/n�C�c{�w]�B��HU�o/f���ظ�q�cF*��h�*lyl8�%��lN"�����D�����Pr�sY�/����%��󽙋��v��R���9�tU�`r�i�ќ�<! K}xp��o�^:��������S���0`L̼R�3��,�Y���L06�d[MԱQ�f[�s��c5|����g�l�o&�
s���a1gWΚ{��	�i���hK���_ه~�JJ��L���R�����L�ԭ�To�9\�R�(��c�����8̳:������S+��Zt�0�H�!���� k���u��=��֨k�N��L30�`$'?����2�� ������d�-[�~	�ے���)�?&��Z���+1q��haݯ叁4L�}7����$����\C�r��ΐ���ܵ�3R�ͺ�O?��&���g�E����ހt�[��V��m����i���_�k�������s 똡6��a|�SMĿ��^|RNv�81V�����QF�G�z̾�Vݩg�l�73�K�W���X�X3,���TO��ṫ;���Ӵ0���V@v��6�p��59����)��0�q�QB5j��zeԢ`u%)�y��:��k� NKd��3�t+�/|wN��=j�����$w�'� z X��7zr�<x��l����bLB ����8?h1A6�����٢�S����r����lH&�g���|h�0�v��w�4?���wC�K//Y�F+&X�փw�����kz��hG��

���Xu���{g�ſ��/u�L���&AY�0���Ǌwʉv@_W��ACu_��I�O���Ҳ�L�-p�����>3}D[v�9n�Gj<'�p\���(C}1�d�]۹0����+��TD��������e�Pl���fJ"bL���r�h��0;���;a��IfcO�Ƣ�xz؞����:���.�Ɏ��������l�g�c_��x�?�]�|�Wc���I��ga\)';7�NG���y�PuEx [���yq�{��gk�t��F���ݼ��I�:��I�k�����#�_d���qJ2,:ȿ}��~f�:�I����Ar7gq1{F���|4��#�\�{��S���
����矊\p�3��.��*Y�<�Xg�7��v�#i��WY��<	�r�n,YC(�A4��\3�Ҳ�uP���Edh0	\׫���#�b���I9�]o��,��X3�Q�*p>]+_l�+��w�]ۃ�oa�'9Pt�x]��VoZj%��s>���d%��믲��DҏЎ2��s"6��I$�V|t5a�M�T�=�Qn�2�g�ð��R�}/ݽX��*V��P�y���蝶c�2 �޵nT��m�;���Q���f���&\1��K�"a2u�6��ѳT'Y��R��=��!G�����K|+?N�?;��<��z)����K�5�2d8�J�))H�9+c���E4}�����I ��S׫�x��=���)b���������|�O���Aԡ�_H�8U�l/�4��x���0�0�e���P�����1���ʵ��?���U�,�7�$��g��9�P6xwV�ɱ[fw�$ie��
s������+�-2��M��t��Ρ��]Wn�2냃e�=�-m�vXK#V��R��ɲp�o����*��uW�0����(��L�e��S��?�<����`�E��Q�K�D��^Nl�j�4��4ʰ����%�~k����m��e�oqS/L��������{��*zQ�7�6V��\���J��g�'<>D}�����MW��k���g�Zj�v|nj�FMj1�p5o{���g�Y?�}��fb���}�B�J`�N�X��f�����Ev��� 뉿֎��lIܬ���J^.�uss��*F���řc����减Xf {�9�ۍ�������Aj��Z��9����;��~�!^"��gbKT:�SwRp�a	���q
#{��_\dRx?�_���,3�NA����Dǆ5�/����u������H���|��Y0�,�O���&���<��F��))��9�!=�A�=���]����R0��� �u������\�A0�����v͓��î5ڢ7������Z�.�K������=�~Cx���t���J���F;ԃ~�8]׆󆸞\$��wX���x��d�� D1��`��XPM��3��Z��v8���#1��(.Su��iWG|�Q��ҩRC�h�I��-�IW��/�\��ޥL��XGG���
�?�W{v:�K��O��x-�G�V��o����^.�l�����u��\'&Z�[m�L6ܧ*��S�c��]�Jl�M�9�V�hwU���ٰ�i�������7t�4���lj��{���&CU�^dYuLKK�~w��_*Ƒ�����٥L�'��M�v6��D
k�"<y(�kq�t�����������D�;O}
+P)]����� t����ba�Bs��,����U`�0��3�/��s04���=�_7#�X�"��ڼ�-}��a��M�w`��L/�_~�I>�)<O�g~����!�}&�T2w��=�F!��f�X�
��?m��x';�x�Q�����"��(��8�4�|l	ޞ��R�K�1(���<��t��D\t��޵ݷB��k��Jq��\�����}��;�RQ��Ww��k�8�<�&����o�X/go�V�
�^7'�OG��3Cm
���_�p�Fu?�e�&�$$�D#�C�4���&8j��a?��[-�� �v�t�����'3��@���l6(+e96���I����x&��>,�XqX�+��VV���e����i�y']Zu!d���p��Z�S�>�Q
�"�<��X�g���3�:k���ɻ��.���b�g��6�3��Q�t��]0�]@hI �E�p-���r�����MiV�I�9i�U�h1�zD���"���GM.�&O�3�dw���b����ww4�� ܳ�����V�u"|�����I� �f5��2#=q��\��=�>5�\FƇ�p�� �37Ȳ]���M���������x�����v�#�e�ˤL�}y�20F8�	��u��^�bΠD�ٲ�&bA���%6^�e���\e�]�鯩������<��T�җ�_�
bFur�%�����~���"uU�#��X��Vĭ�ays�hVۂ��t�d�|0���_��.w����E�w��'% �N*�:q�_�AO-��T��F���;�	��A�uUsK�ߍ��/l���x�p�ӟ����_~����վV���]�3�k%��L�m{���H�{~B.6�ý@S���SN_��@q�Mq0UU�����T��ˤ�=tn�6u^�6�'ׄp�Em�w�wб�:j[j��-:ޗ��zmk\t��*���|E.��3�c��w�i���v@��x�gnV:��ӽbP�p/6@�B��R��X���<�]~��9�������ֹ��Uy��X(Ͽl����3�6e���*���SƄ�b��t�o���w�/�e)1�j��(�ДO�*FMe�9�с��Yc�(`�=
�6�-(R��F��;��"���|�A�@�,Rg�O�i�uz7UɿX���F_����w��3ʭ)�Cm�-������_^>WFƃ���6�tlX�u>i"8sC��:���8������ٛ-�4w��ݪY	�\�����|��L��ޙ�W��~�87��_-�+�#o���<�/yz!����i���[�)]8�� ���]�T|�W[����WHY�졁���
&:���X�0j��Py�Z {�(����:H6`u���c4:#��w�I$d�x_"x�����T�o��s%�DqZ8{�a}w�}�-LX��\i�f�z#�w��H_gus�b�j�A�Y�����O!Ϸ?1mmA�M0ݳvj�5���s2��a�HuM��W>�&��k�@zs �[�[�E�ND��>K�����e��`���q�y�\Ɲ\��{h�O��W���x��~f`̜-�#����e�{�,qv��ij.=3�Ʃ����������Z<X:z����`˲���y������L0Fu�ZH��52w����L��?Y�X�Ќ��1��l�������5�/�tI�M'����L�B��qo��l���VN8�x <h��� �u��w�-��������n���PB���JHp����x����T�8H�:�zr�=������
��34b�V�	j�3��Liny])-�,����^���] �}���c���p��z�~C�ה��[Q���ָ�n���5�����R��` ����o�<�~!�����pSn��:|4��H-�K�j��u�**pE?o�)�y��Z�O[M�{�����	��9\T���0�:C��>N%c�I�/}�����oƠ�7�/��kEa����ochp�?ӮQ�G���.������Ͷ�#���ke��E],��b��f�'���l�4�>q�ܧF���Ha-�Sr���X;�6�f�L�q�O�N�/����pN�s�q$��_=Ut:);�=���l$m�c-Ii�(���C���-�<�{=Uy��0���Miz2ܑ�Zf�9�I(-;>��Ł!^o��"n��oNR)?�/����4VjH�Պ"c�׫n���4�����8��6���ٱpclt��__� �~ ��AWQ�&36N/�*���t���i+�>y��8y�'L�ݕ�md1e�>�2�GZy�cP&w%��؄^�ρ�F
|�q0>�Ú�R�8����N���U��Ҩ���F G�������ߥ�o��K�u�k)�'3��c�9��* ֆ�Q	of�a�0�h����ꤘ�+�k��}(P��4ݍ�P_���5Ga����gW#�[6�;������|�nf�,x��\2��$����Di��#�v���l�m��zk��"n6@����\ꌬ������H�yW`��~})�W������7��H!����b��"�XS\u�W�ǥ�'��y=�cz2ٸ�k��c����S]e8�����<3�-+����r��mdc�������:x$5�1<|@�ꤘ�X�S�ĵ�?2�S�}s���s:K->8Ny�c�
糲����uց�Nx�pҜ�W:d~�@Chb�dUS|�n�չ�ar9��k��݄��n�ʯ���N�),Ȕ 6��?~-�x��՘*4�n�K���3����d���	19�6��ަ����.����J���u�1{�������A%|�?��2PT_�}fV&��VL���[8LSQ"�ܮ�to",+���#�;�Wa�i�������{��8��G�w��U����+���Ӥ
�	{��%�F��x������.��D�
�냃���?G2�*k�1�����-@�z�WJ��Jw?�#��{�4*�n�fQ}����`�&�V�s�ҵ2�%����Q3��S㦮X���ț��/w5�"���L�����e���1ݲ=FY=:����Q��A;���%��Z��͖���G��_�dͣT��T�c��� ��;��Kw��~-ͧ��x��4��XF]ѡ|�J0�������Bc���V;ͫ1�⒝��E_��oZ�|}�=�sIԜG�C��vB�¿�J#�}w���K;\�Ԉ�O��y�ZU|h�O]u����ܙ�����N��|��߷����ݫ�<�\o4>;HDd߈B���;z�_O�2^�7��d����Vc���^1�I,�{m0N�����(�˟�K�l�R�0�AFH�{W����YhAY����M�HO��p��Z,����:|���%���IR�^g��:`���`{d{��u(����o� '��"qe��KU��%��Kl�����|y5Q~�"C�A�P�,2��L��~f����!�E�XW
��E��=JIw���6L�����_��mSfށ��K=�Sv0��[٨o�X�����#�v�Ics���ˋ�1�U��uWG�h��9��/Δ�~�:��b��n�
�r�3,�3�ȏ�Z�c�q)b|�&�v8=����MC���@������r=��.l
�E@�BK#�'��`R;�I�(K�XX�m��)�4��ɨ4�H�^t���r���y,QM�(J	��
\���,�� �^����3�x_�__�o)��,��Q������z�	M
d���ū���N���]�!?��N��������Q�"���'��u��*AG��
��!fO�dn�'��	��*�n��&�C@ȔP*���扜��V��A��w!����$"A�(��  �N�6�]W�@ F�(�.R�l��:�;���^����D��U�4�W��'r���ך����8���\M������6�����t-�J���b���:���[O"���+���^�����A���Hk׾��oS�҉~0�Q���|:qZA���N&K^�Cx�%����'OiL$��F0��d�Bn�,���/�9m�)��e���)K�i��/n��<,���J���O�}s�>J�H�N�#p�}�d�&�GjBn�8��z�)K'�e�Ց�V������?_oM̫��ص=���`Q��O[&���r�{m��x�~֚NZq��ػ<�kT��%~zd�q�.��912��()������=�TO��K��a����x�QNϮ*������տ�q:2�����6[��V	��E�MR*`�l���M���b.�γ�F��u2m�0
���k��OKl�A�F�R�����������~%M68��
-<��C��ÊǬ�Ш]ڡ�ks�A��N^���q��Jە͠��-%���n���ވG�VI��D�Z�� %xO���T�$vȲ���믿�#�4��d	1�Ɂ��Ң����(����:��i;pN�:�]�7�1.o�B��B�׾v�}�݇�Q���_��i\��6 ����6��`����H,�M2Ǉ�g�����#�2��"�uo/� �}��4a�:�l�PԠ`!�*K�}�n��1Έ � 穉PZVs
���p�5���4�U�8�z��'@޸{A���s��f>\%p}����K^���0'}le�|�����(��G�>����+�1��u�|�)G���6�bU-�
�p��O|I��n��)�e =���yRQ�d۰�ZWY	����Hu����韬.?�R�5���Rim����N� S���D#�U��P�ƥ�e�8_~�u_\!����� �H�d�@���3q�����
�����u>���l;
V�e/�@�ʵC����S���@
~�G�����|WqteM�~7b)�q\�/��2����U�����K���P�8���������p�X�n��
1I��3�=�A+k='c!�����5b��̿�"�Tl~-�4���Q&�t;�[�,���{j��v���@���ߕ?�d!�v����}.�2�k��2�.5�q�J��]#[�� ��i>�A���i!�_a��)הJ�b��l�7Մ��o)���R�|n�Tb��,@��.j����3#]��'e���jZ��z���}��md��u�a�T�����J��b���lG-�BF6�,�c�]$E	��-E�����q���c�:*g�8�S"K:X��s�o1D�@���#2Rtg nTDw�Y���><�] �|r!~j��P������w�:���B��������A��i9����33=9��q6׬�SC����@z^�u�/���-P?�Cű��.�V}WF�Ȯ<�%��A����@�������r2�k��t�c��De%���y���X���x�
N�w`�}u�������o�Q����?����O8�̀�PC�F�>�uw��2������=j��G��w&�ͧ���x�N$Q�ik?L.籞��;�bڔ�ܖX�ⅰR:J��-�׹��x�7�j�59�M6�i�oDQ�&��d�yC{�v�s�#`�-S7�qe�:�p"�W��D���s%R��_�j��E���p�����e
g��x�-
�/a�~�;������`qE������Q0���̒
�����.R��K)��k@��,r���9L��~b�s��I����P�����R�����K��2ƶ�3�p�8�g���L;S:t��$ʿ���xq��V�|��3-�cvS �Q����"��������ȉ��Ã��ޱ�����Me������{^���h�b�}�x�o����!܌�_�9apj>0��B�j�oޤx�7W4�w���L�
w7%�(Ac�܋��*˹��m�QX���
:>�t�ޟ�Q�[q��P%��=��g��5P���%��V/�^ko�,_��v�.y��7VL���<���IMd�m���&�k�C!�we_��m1S�k�'���g�z��^i���OU�����i�QL��&���Z���pG���>z�R�� 1?O^��P~�
��gdU���X�|~e��p6�'bB�IP��2)�?��h"��8%�k	i�(����<Iu�]��DAɉ��V{B�}f�S&���S�
�,z4�r �2�d��r��|׆�ٴ�r��_����BJ̕핛�ݳ������ ��A80����X"ne���^�޲�=��dD�~�ޔ:�Ƙ&��_ܡŃ��4RӤ����7b��Ͽ�S����ؒHɩAH�jy�)[މ�/x}|����ߘ�r��_������sB��y�N��M(6��D��ɴ��ަm�"�3����`��3���kq���}�=#@��δP�͖�����ֱd鮄o��� ޛF��>����r5�q�_P	�wMR�K���`~��'s�����1R~�A8d)�k���ؠ��u7��Y��t�	��66�'�
��ʰ�o��r�`K�h���v������y�����Qal��^*�jZV4$��S�լ����nݗ�|����]�P���~��{u�+\�u�-��3�t�	r�D6�����nv2^��_��P��`ꁛ�x�M�I��R�T�Jp�vS�6��!#��^0s_.hi�!���D��M+[@�G� �|��cU��U
6N:�̎M�_��(�CS�8���b�̏[`}��7P��,z}}��ݗ/�L/�T
��zy�a�,��R�	Jb��-(;-�QlZ(#Ǯ/7�s9���5�g�};L҅����?�@�L��`@$.V*��H���=�T����ȿ���/��_8�y:K�`5W�����:̈́��h�\��b��ץ�+-<N��zJ����9|PpvY��rsE��;�gB'�����'pY�u1�:C�-�ܾH_�`x�sr����@%1W��Ls�\�3�A����յ��\jU�@�C�9M( ]^��~�$�u�vW�������c���Z�����uTyL��Ca��ą8qh�{�����N�鋟]�B�8z��9'9g�K�͵/+�η�e�6bv���	��ث�Q�M�Q���,�ר{�q�6��z1�����'=2'N_u�Q�gw���C:{�] 7��2�[}��=���%ݩ��w'����@#A
J�������eL ��m�OO� =���Y�T�z/���[��e��i"wm�ApUiL�>��R<��q�l�a�<��M��n8em���;����q�����#�-E�R��~�r|�|��������3t��G�+�o_�0�'v�E��@3چH�Ye篼�T�v٧Z#x"�g�������Ϭ�d7����+�~v���8<�9��
5���8j���N���J�pf��i��?�	��\[/�t�')Y��M\�O�a3w�eأm�T��&��n�@C��yTwL.F� �V���j����k��T�ȫڶp���͇���$���=+�.t5B0۵��w~Q�΀K\F#�)��!䫛U��?�U�sk$��P���Ĳ�A�lo}�Ӯf�����7���;��v��R)%L}�E\�œ7���2��@U���NX��(*��PkuUL	��m� 8�h�La߱&��qZ�z��^��n�!��N��C����n�Zn���=�����U#����Lժ��U��4\��v�t��ה��q� ��2�
xVp����Fc�=f��P�zS�.�l��g��e�қM:��"���R�l4>kD&R�����C��2l�S���5��GvWTb�w:�^��]�7
����nK�˳����e�:I)>!k�2uЈ�>���`a�����M��0�P��6-ٵAz����_�cv��mt:v�M�Z<}���65�46��,���F67���_ .|kSX�_%��nx����,���dū�B��	\i�;n
QϤ~وK�)4'40�R�K)	���_�M�𑯅��Dq�j��R����tʚIG;�y0�}�u�O�+�@3�}w��~e���)ֽ���~�����w����Z��\�y�0�����N��9l��%�
(��Փ%X
)Ur��g�޼�uN㙔!N�� �hv�$���8�b"�������*�s��`lm��b��`���q�l�pT�A0~���ȆR�}^~⟾\�T�Q���4�@��&e�������D��Y���\7�u^�͗�A����+�HP��EY�n7<����En;K��efh�eQ�nf��l?3�xsH���K�*�3��+�6Ov����]Y�,�ss�~{/h�����l����d���s��<���-P v@Ɯ������ �kf&n ͞]D�/�a������'X!9�Ek��-^K(gG�Ƌy1�ܽ� �@6�)�z!.\��6�c]k�t���*�H�u��R��,�V���`���G�t��c��-Y��撁��+#&{.�x���d��\�Xv/Ǘ�w�2:��|:�+���Zi:�#[��(��[��k0c���v}6�([I_�s��i}��/&�"�=�|��dl��yї�-,�&S��e�T���Ԥ1���m U�X�B+�F�����x�����Y���"��a$f�N7��J��E�)�e�I���H�I������4Ը:oA0Z�P���3/]��K���~'���@�LP ���
�	��H�m�NlW<[?W�P���m�����,-#�٨��`b�{e"{�M��=��)�˫4���!*�B�}��2�q�nvrӽv���*�CT̏��)#e�	��C6m�,a��&�L��u��(lr�ؐp�3�"���f<�x�ceW71�|�{�b��?�t*�k�X(n�:�"�?8 R�u�����<�����/�Zۍ@��^���y���ێ�!�xTAk���µ�����MwN��sH�iPV}�=�a���ܰہU��*`�J�F�}Wa����M�rF�ᓢDJ�SL��N��o�x��p�e9� `���c�1�l�������R�7��@���w���{�\^b�������F%1�:؍�y�I!�ry���N&�&��1rP-��fX�@����@d��tR��3��p?0kC<�f�&3J�D��X�}�]�-덇�x8q�b�"�I
HT"_��C� ?��z�<�_��Y���q�#�}^��	�}}7�6�՛����昺�ť���@��3���Y�����zD\��m�H;������5��<
��z��>֬c��&Sp��B�ƙ�����ͫ�нR:���ᰄY��5�m��0���ck3T8�n~�����{R�ah�AM��-���C!}x��
�(K���{�RjC���X�!����^���zt���GCU<���A�@��X�Gi7sV+I\%౽� �5��kyD2my���G��Wke�,9��Z������vϣ��|�˰[��f�
Gޯ�7ӓn��b����}�H��]��� ��I�H������܀���_�|�aA�p�D�q�Mz���&\n̓��B���eX|S���V�z�t7�f�I�5Màϧ�t�b��M���C��/��CU!�wȒ֚����vR������W/�����@��-��H���:ƫ&r2_o�7�q>�R���b³T�|�#��֎di�����R�{��U�R�p����d��tb�����y}\M���c�&��󼡰Q}jU�k���xr��l����3����^�D�8�S�0/�Ц�`��e�n�b��~��rQa�����P!�o� ���bX�0����!FnG�>�D��z��ǒ�0Qfy�ŷ�������O.WS�p0�ƚ��6B�%}�g�a����t�PTOH�[�ڸI�ƥFq�����̓!f��`���񺧳�2�*�>���j��|�t��ܬ}������e�u���3��SK�#Ҩk̥���E�7ͦl��+�Ԕ�� �͕�8�}��:mq��#�����⩳�F�y������SE�=��[�̦�����@ ��1�/��D�����Ӷ��9�S�u�Au�|2��i�X���$�1�M����&�K�~�woN��c�������o�/u��(<M�K��q<Y+���r	.~vz�*d\ۮ.g:�#D`�@s�4S	*���T^K�]+��%
����V���/�ŝ�⍮�Z�8v����C��s�I""a�K^�>X���_������\�T&��I��V>��Xz� Yq�Sޥ�,�S68�>&X���N�#'w�ϕ2U��3���� s1G�f�u����j�p�հ�����}�&u`/�^�_NVC�P:�Bx�����h��1L ��]C�e�oゖH� �x�3� l��V�I||�>�z�[*��nh�A�AVN���ҴhT6��8��*x���+��a�r6�vL���h�i���7��n�#1�>}�?F������T;W�3����O��KM����Aʕ�)\g6:q�C�^�B^k�d���lj�'Ns��E��AJ�d��9v6[,;�$>�R""�;M�Lu��dů�<O\K�zAc!�DF�E�M>�Ub�����I���WMA���LgX�o
��LG7qn�C��e6d�e/��W�N.����U������
�g�߳�:x�N+M�|�k_9�����5�l>�|���[���SS/�2a�g]�X����ϞL<t��f��?�1�C��C�"�Q[jCZ�<"4k�W�[5|��Q!�~�T���*��4�����p:���:�">�w�޶m�
����U^0��u���z%������̭F��g�㞢TD�t��H�7�FP��hhTά��`V�����$>5Ϧ�I�ppj��4��z�Ϧ\�!��͕G��hyOk�;����0s�>���X��Mi�cD}�#l�_y�lj�sx���j+'o���D�(h�m��k�<&������p뢶��2��~V�y��F��9ܖ�?|t��f�*���bA"������[M��)�:9�,���;X=`v�n�˥��a$, <������⫛)�7��ȃi�ś{���*��Sv�XiS"߯U�*���]�q��Iq���r�s��J&�_��Va�A}�olNN�s�������;1_���L̙�>��_�����~E��x����9�C��o���%�Wg~b��MƱ���)#�iv�����첓(��K�bVs47V��^�q	���.Kq��>|���[�X�4Q`F��M��tXw����q���jE��2�s�p�J)Q�=���%6��-+��������'��]���?����%� ����y0�������o�+�G�2q��?X�4:	3�+�Gуo��KZ!�^���Y4�:L{&6k�cխv�I)��>n�oBg�Vw��m ��+ѹ��ͬ������FE�A�o2���Cqd/Q�>��H��*P%~�����O_�m	3�� n�>UA���� Xvvr�?�F?Y�Iֱ"ccS��t2ɷi�1�"FD�8�l�v)˩QfX�Zo�J����ѯ�����vs�H�����&��|��5l�?wIPO��8ؠO��x~d8_=�q��#��F���B���x���\���]�w�쀠�b�qf��O+�<!3����8
)Lt�7�0ZXe�<Hj�ԷH�3�����6���L�c�>d�y�>��I�r��\���AM��`��j)�c��0��bq���Im&�h��~������#����}���{LVlSsb�� ��\�m���5����<��R��`�- "�'q�U�K���$:D�c���p\��J�K'��_��_�P�ۿ�+?�vx�6SS�B�I�+���ĺ���~�u���d�2>��;�-NL��1/�_�?��:wc9�&������7wy���_�e�� "b�T�hn�l�q8b1>Äu(��2���}�?0�b�����d�asKmG|���T�� Y�tg~��ؗ��4Â��!
;ڱ�t.w�kc,��F	�$��Ju��uI�Z�,5�j�t� �F����W׻*U�k�;_�S��tu�5xD~N���L�`ۇoŋ���]*��RT��I�f�Y:�P��/[ �Z<��8�:k~ܘ2F�]��u���ɫ�v_�;P����R��ܽ��'s�_�἖p>{�KӇ|�>����'�׋�6��]}������7�"�F�5�22�qG`ӓ����.�4\u=�A��ڎ���@$e���++�4X�bSÆ�˟�ˠr}fy��uR�"?�􋼙�p�͖�3lCh�J�/�ٚ�f2�+��OR��_h�n� �oO߫����hG�'���fó�q�c��Ï?2���˿����X���ȥ%1����owilA=�G���/���֪k?Ն����I�Ib�h��O��߼��v�����H]���yc�n�Ӎ[ �->�.|��^�z��=�Z{:��3)��(+�����D|�(��+D����'�c��_-t2�j�� ~R�y+Ǯۆ ߭�@s���~	�mB`�){�xc
�ݜ�GԺg�$E�fJ*�\�$�E�D�(=�<�\�W
�`���9u�w[�����x/�W\"��Û\�*X]�.U����PR�hf�0(m�w�i��ͫ�X�����m����������J�NO!t�,|+[��)��9�����=����^�u�kt�NƱ���>Y\�	��&EUO*�P��S��l��
�A�C>�5�L��� ���\͓T�ū�j8�w�1��n8`A۟#Ix��o��2SBsi�T���>C/d��Ǟ��p�H[���Spq�}�]�>Ø��7[f� B���{���*\!c�]�Pf����5E�e��׻&�"L�)�+5	�j?�� ��O<Jbڸ����3b�:��U�`��ާ]�V��)Ş�W��j��=�KR7[Ì���%K���5�?u])m��}�޴�ޘ�0`�bܩ�'�v��"<K��RJ��Sj��^f��àE��)?��;	7�n�We'wz�?9k�ƣ��Ǒڥl�1���E�F�&:Y�2.�Ƞ<�;���3tw)n�����9�_�1k�/+G��|��;���:	LO���#�[�O����J�I��ڶ�m��8F��Z��YpUl�N2^�M����c�M�y�wlNj��F�y�-���d��13,��O��	GdBPw?nY%2�m3�c�`�ejU_�����~|B%���<�~bP����`���9�j�ƹvg����Ayג�a�[uv�ԥ��Y��3\5cN��`�o��]�!r�v��)_1�;M�]5�ò_���l��b����8�z3����b���&�M4�Dy+���-����Llbw^{�x����S���v�!������\�-Pa/�w`�H����\zޱ�/`t������t��ζ��${���n=<=�_��33n�@��~�~w���!�ö7�z�l���,η4�Xt�OAU3�c���D��O|�W�����P��d�]Wꁮq�H�BUV<v�4���Z�<9��H1-a4�y�O�N�R���9r|p�"�~>J�^_��t��;��q���R~����]y,��㲝�0�Cq�����v�x�l�Rfa����g���_[�Cj��Wj7�;\��Tʫ��N�X.nH�9�7Սn�`��Ձ��&3,x8�(������/�y8�KU��c͖��.�"R�,��m��(��X�=Q �/T��+�8����m�˭gPE�,���;~_�������>��{�9�b�B:Yٗ��������Gn�����O΢���L�`��P�rJ����
<����L��̩�x���ޏ���M��ܤ
z�G�ͅu���;O�
8sⵝi���+���
��>Ax[t=��H/����0���t�;�HlP����̴pH_�{�2�sM@�蠐͖��^U����=&�\��~��O�iYp0#���N�S�:�;�n��"�k��gLUa��� 
ϳ-"�=l���?�"�ʠu�zy���H�q�u <<�y}���7mkH
^{����80�QԵ��1n}�C��A�&�v{fО���b�}i@��N�{�~Hy.X���y��������w��&�� uv����|��C�8
������E_]*0����tw��ϓ�$�>Z���)�2d�7�}�s��U�/�����D��x���_I�|w�}H%�`F8Cs͡�J;vX��\���D�p��Nd/����޳n*�#��8	���L$����Ҋ%`���}aɉ��0��~"���,.�e><������
3 ���@���T��7�xxdjG@�0����6���>MņE��ּ#�� �O�	-'�;A�%�El�m�4gW$ڬ@ g�	�����o�+��+��sTy���8��J����<�x�Q%=z�������^�o�$�7Ԉ�atƟ �Q��2�1����$%��� �"ZU߂gۙ~F>��px���.�Pa
H��SρQ��%jO���N�F;��0^��6�pe��B����Kc��o`����5��`��GN�/���N!��.T��k#&��c�.��J���#�"�_�\3�t�������q�,`-�8��ũ�E7g2e�7" g����?����,�UvEv�]��&�g�4˄�	���-�����fѺ�$)?<ý�7'�W�V�Yj�⏦W0;?���|FgW���T|�G���6~S��ɺ_ ��.mZ��㺊�}I�Je�N���~)�2�ژV�����f��l�-͡�Z�g�)QL����r��B�Ɵ!p��P8"Y*��j[����Ar��Zù�Y	3yt�7Բ�g��&�lg7P�fݛəd2��o��<��������A��]/|�:��� ��p�QE���{�%`
��<HyhR
��(��wσ��Gv�3%��!�]�.)�f�
��!M�YW=�8�q�<մ�(���Jp���&�vnU�Mp^��ݺ��23F�ٸ����,�c�-���ƤٕY�{�X�;k�Koa�������@��6f��O	@]=���˷����)����`�2�eY�/��z�l��X�0��	i��F�hp���^��쁪v��Q��Ʊ\��hτᔇJ.�a�)S���)�g���g8@�\�uo���b �R�����ukJ�n�) l����_��M��T��T\f(��s��,�ۼsF��ܾ6l�wyn���K��I�J.6_4y�`*��2E���>n�BL/�,;H�;��b�e��?�䡇�S�뻲���04(��v��y ��<g�y��V�PP��+�Xwq啃j1͏�-C_I��<���櫍��h=`�\�K=�r�f=���&��GWrً��|ئ��CmY��y��>�~&�β���=����6$P��"�#h(��xp���>y�M�i�
��7ʛ3X3kHF�X�Zik�f������U��vBQ�y6ѦY��y<]���2�R�}�M��Y�i�:X�M�{o��o�f��(��xg,K�'c}c;Y���+Vɛ�@��Pyv�f��C������I�����7��rA|��0� ��@!�S��:�l�����1�6�L���7�,U�4��m���Ԫ�*�q�D��ݱ�F����q&�B\6e���pi�t�Cv�&��!�؝Ovf�d*(W�D!OBE�\�J-���H���ښ��ڔ`g�Ŷכa�W��.:]�f$��yV>?m���x?n��[�iF=J��#��뾽�'�m�����(;���Y%�z�;�>�Z�p֕�ԍZwI*�Y%�/�h�d��(���@WX��wQ��4�Nk�|��z��'ixĳ����u�\M}��i�i��}<5�3|����l��|'!�p�F4����Z��"B+qϲ�	���DK^&���PM�^fB���Ì�MH�g���H{��/�V{���Q�����Atט��h��u���[vJ3H��ĉ��S4��xS6�ѸL�d��D�S�̞��x��MK��;��R�&���x}i'hW�d��o�`�.����	T@������� 9�^T���b���q��kཡ���JÙ5��F��P����k!�CX�����ҩ�J>�<�nW7]n�����)�}�2İ:#��P����Wu.g��$�6��9��>,����0SU,��1�S����_�q��r�Ag(��O ��ֵ�C��e�|����`�1I����*=M�v�k�C����J����ƾZ�>ȁ�{7w���A����n�L�kȬ������揶+a��Vq]DZ"S�`D�c��y=�z�>E��l}V��:�?]ūU��k�%a"�I�e�恃�9WM��k���$ל9��J�P.ŰY�=M����ap�v � ��Ե��.h�Q���v�u�Vǁd�f5��h�d��xN��j��`�I�e���)��������ʰe���Q�&�@�((f�>�l��%�Hz�~}	�~�HX�x���e��\��]zrଈ�2J�^�c¤P����q���I���Rx�������"r�����ط��Nl��
 �jz��`�����Uz(\q��{�����T��Jf�]�����ܥg�@
��f㽸`����0�����;�"c�F:��[m�f�H���`O-��8H��Au�����3;�2�^+���4)[kFaFJ�ZJ@���������Z+v����y���z&/�����$/�Gf���z����q/�>�v�v�2WJa:�U� �p�+���8���,����ڸ3;�d�Ս���?:	�1�az��`�w*��>M5I�g	�����Ǐ<��Hb��s�O�c�1F����FBw�/�:����pk6��ܡ�Sj��>���-,�o�8�Ǌ��V*�sϦnלI6:��7e�#�&1�C�vIX�J]>gG T�7��i��D��7�2��Ycݸ}�Y���վ�
�s|oj0�FJUQ"�|���DGm09v>p�j5U�i��=Uӷ�˒l2y(q����د�'}f�!>�Ƙ�������tP�O��1�E!N\�]�Z��j�bC�;���Ql �e����en�����oϠ����չm��٨,�o�0M�k���}�Dϵ�~�5V��0�a�Ƨ;¶l�����~X��2xť�~2���7MMt-С��5�p���j��L�gZ��G�z��3�󶻻#��N���t������G=1��3�<���w�꣉wH��ٽD߂@�v�&�=.���{�h����Բo<�jF�%0q b�I�M_x��4�[�����Up_k��K���?�r��jW�����_�M���,{��P������oF�y��� �ՕO��=���Ѹ�;��o1Oƍ5n!;��?���tLCQH��:��(���29��Ep �����(��#5�����7�Yh�k��p%p�N���.+m���|̨X(�4�	ZK4%}��t����?��792k�>�å^3�N1�xQ���<�g:��!�d��B;�,��K@��7�+R��c짛;e����s-��a)�,��7��N�+㓭1֔��l�e�[�D&�2���y0�p?�f�%������ژ��,Q�᠁��Ws#�N|{;�U�w�)3�mY.�����Q\^��v�W���G)����V�PS5�OSWKmD�z�X(��tiUÕk�7\��3���J[B̮ջ��:��M���&l�t�]���9M�V����Yw�(a>��C���b;`��Y�m?�A�C�
�;���5�Ρ���>{��z7Z��Q�#�c��6�����=>-o����Þ���� �承���"Cw2Tz�܏e:M,7ɖ-&X3�A�i����S�\И��[�v�J��9x��d��)�Rk�c�c�swA/�ucF�Z�3k9Z?�f��0Zj��l�ɾB<��R�ڞ�q�@q#!�q�M���A�H����M#O��)3Vԩ��k\'o�Z��u���/m�a� F?=Jq��f�ʨ���m`y��*�_�s�\�4#�8%gDsqk������(�ǡ���R) EÊT�Z"�6�!A�gG���Z�3B`^J���+]*>�ϣ����b�c��M�"v�]��d�(��	q3eC{H���T��^��\$��Za����PY�HP�{mf��PX���h� ܗ��⦨�}v�V�c6����� �a�j��J	�[쑗�����Ҙ�^UU��J��.1R`E
�|�����C�q�%*t�b)�K�l�Y80�u�dS$+��+�	�Xc��QK�#_�hC�`���P�]��v���k2����Hs3�-��t���q@�4��f�y�H�lu�U=�[��
��(|�4lPث��Q7��%��0Հ*W��MY�.��v[����,2����4�5� 9���JJ���KiM���٣6�"ST�cv2�����`��4uᢽ^�8������?VL�U]�8jx������L��U����])q����q��۶Ŋ�~�[��p>��O[i�$�e����:�q�d���]l9���Z1-q>��������/�c� /i����˼f�ֶ��ut�)ϚW��g�h$m�W7I���16&Qr�cѪ�z(�ĕB��.1㛛/Θ��[�l���Y�&�G'��Mi����>/T���I7�wj��Ln����X���F^���qۗ��"�K]Cԛ��k��z5\���%>#�ĕ�@�?lz�De�tlJpL�HW7�?S��ӛDN�p��P)����kb��\qiʾ�qe�˛N�Z�����O���H�F�`�;J��_<m���ғ�[�,�#����J��	�\8R�K
-0^��mR��N�(��V��hl\Es��`�%�X��
��I��؈��h���J�Ֆ�������;�>Y(燥�oj)���m���F�(�f���7�@��H�� ���\!���FA*M��ĎA/���B<����:�.��K)Aa���p��TQ?HE}�[�ƌt;x�- ��������ޒok����1��>��tw@%>���Q��V�db�V�(�nܶqZ05i1���v��4��v�H��G|��ZaFxO�߂�ӻG�;�o��7�
��؟ �\=f�{X�%�*�_c�J��hm��r2��p ��2k�γ������B!��Z�b �Ǚ�$Ě)7y���:���x��(��;�NI�����e�'�`h��U��.�6��@�
Y�(A��ˊ��52�]��L2鸴�\��e�f�-����������O�<Y�@\�6F���D�٧�FEO��� H��v�3�Ȍ�D�㖑��IڱM	��!�*L)����8��4��LQB�V���ɢ�Ň���6��f�k����mŅG�M�yn��բ,��]}��$��a�_����~����N#������Wwt�T¾�������z��-�V��u<�*��/�~/����e��3��#R�9����~�:f~��� ����Hl�e�4,L �L�[����[�Z��o]FM�����`0_Լ�&��@��6���>�ֆe������6�V#E�7����H&�G�%ّ�@��������^���`U��s�s�ք������*�q��U;ƚ���(D�_^����+	�rc��'��r^*<�DTy88�@w��J �b���>�b�&����ul�2�ci�/#_#���ۋ���Y�ʬ7M:	W��D�Mu��|;ҾP/ .�����k5��o!V��s���W�)	c���?H+�� �{N��1c�O�`^
"{B�8KOQt�fO��ˏ?��e[9zF�HL�*�fj��"��jA�?~�/�����5_o"	��{7�H�򔱣��UV�&�+h( �\����ߡN�F�k��W�wS�z�4��vn��-t�����6�a7D��	)�'똲���2��J���H�E���h=>l9S��7�O<�y��TX��d}��5�M�.#�:4��1w�y|.�*!`uc�&I'Y�e�Yvv�+�+�'���//�<AJ(����>���	�D�����?���b=�d���������l�����J�@�5�Ġ�sp�����u��A�V,g1	�������]>R�ִ9�Sq��:�Y֚]���^��/^S�{`�A��������9R��u��O��������C}��G7������)�Qdb10	��L^9{@��2��e3>?��p�}�OSRd��{��K��:�ݦ��@�+����>Wa7�Z0-j,v-����4�����5�5�l�"R��7k}��DP�2�C�A�%.r8Q�s��l��J�����- �mlwϘ�M�u�Jp�rz6܊)�ѣh�(���v&�_ܘ���l�S�(J�8%�j��nڌ-e}��ف�&%��I�`�ؗ�Uk��P��3���I��P������� ,��[��]bhףJ��vX�X|X�q$͂�������G�Z=�"��Q����]J��-�L~��\}�WW�Φ��q��d��?W7�}ȺA��wV5�K��^T�@4I����Œ��j���d�{��E_�����M�P��F9�L'������Ⲽ9��@zoͬ��5#--S;�g��i�����E����	'���C���~}u� ��0`D��Vb�耱+�~�q_GTs
�_`alR:ǚ6�O������Bg�K��)a��!7��#�{��[��w\�_����W!4�j�-}�Zv�=�)ȷM$�Y1��A��^��{2ֲ;��Ƭ�O��k-�Ӏ�-P�L:�k��h��IXq�)p>��R��� 0R=�JF�ũ��u?��Z�C(/� �r�{��^C���� �5�K|t�W�&o�縴F�G�R��5����u�E��+E@0���^a:�<k%�<�8�L`0[v�r�>��/��
9J�K�&�M�d_�T4��7�]%pH�RR|�I�7f��J,��:Ү�I��
�;nWu��yv�|�%�1��/���W�Qg�eo��0D�Rez);1K�%X,c+K�$�eԳ~:<0�Q�	�˶9����<]��6��ٝ�4㣀OT"���T�R�h�ŌDM���q��@f�?�mD�a����+�L��b Ȍ��^��Xb�=z�cs]X�$����>�Z�*=��Y�n5Mn��+�O��Zc���[�
(���T)����ҾI�V�LO�z�3ۂܮ�,�{�Mi����p���O5~���)؜�Q��o�Ӑ����i�1�H9�r@�%JD&pjqn�l�J,s��#�͑ԣ7I�F�)�'O�W�Ndc����l���$�zq@L�xm|Ԕ]��)��X)�p)�r�9�Be�J��x a��J�n���τ��(�yv7V������'@5r�Q�~1w]��b�K��(�a׺�{�﵅�p�����l�4-#�,Vp���p�ƃ5�q�s���V~�;��s��~�3��zN-�(� �<6�8�Q�B�� �UӍ]'s�0X�g�(��h�ㆉ�����k}�gԋm��\;>~�ڕ�6
ތ-8e=������9/�|�רӘ4�������qY��������l�6�z���} ����-�Ë5��ɖ�iu�Ѹ���A1�gC8����vϣ����\b�����s�h��{U��UY�Bs�؜]����5�N�5�0����{=���X~�Q����~��v�`ޕ=ސ���s�Z���і"S.��,�A�S\��q��x�]E�EWn<�C���w�UZ$��1����o�Ի2-4_�3  �o��fg��=W���%i
aaH���'��L'	'�9XU�O&�Y���t�t�M&^�x���W黳����χ�w�s^Ԑ���7N|��cĳ��k��,�/���S�U�:�6�*Ӛk��䮙y0qRjP
*SG9�C�� ;h� �YA�5���i٦�T�\v����c-��,������B��`U"ken�j�
�L6U�P�H?������A%(_'��t;Rz|�䀺�w�ٺ�Gn�B��ų��y�����G�IoT��W5����,����u�i��6�i���=�������,�/�%ؔ�x�On�.�@38?=�~�7�`
�e]�v+5k_�;�T �Xʩ��t�hL��Li��~l:�vG\h�_NW!���=R0K��m�&�`)�:J�	�Y�$��ђ���}����T�^\������,���L>�nwp�(�t�������b��=��r�Zi�Jԑ°d�t�x6Q7'�Ͼ�ť˙�t!6.�{�Nz�O*a!<��n���2���~1�q�ϟ?��>Y�\*7y�^�i+\�?��~��°���zBX��)%A��jY�&�q��V!#�'�d>H��7!z�?�2�v訂^���h��d�ir�	^��r@�iN�	�RQ�Nѱ{�\�(�M�N�Y]�KQ+�z��K{�����Y�9�u�Cpe���z���^��n�]D˱F��2]i�����r{�H.~��8��,�����oAs�:3<�#&�`-~e���q��(�]j��a!��U?:+�%2�D�A9�Aj�&�����3��#�j�����@�� ����2j~>>�ii>�b��¹�
�Zzѭ��#ˏ�'>�1��^�{�EĽ�g:cm�u�Ī�n���m��-߬6�Y'�q�>*i��uܠ��t��7Ѯ��$��T�����.��{W����Y�D��qGv������NZ����F�eyA�U� �%�ɲ����0�ə^��0*�Wn�K����/m��ȑMU���gfw����a{����v���d>���7�jW��T*�y �@ ���#��1���3��<)`-�3U���_����V�������޿|A)*��us��c��QU35�G-<��^��1,U޶3�͹�����+�Ed�7�0�aHc؏.�=�l(�����JH ��qR���CM�4^�m�m��m����~�����?�I�)��F�ʽ���ȸ��3�[kk��v��̂�9��A��H`�R�l�gޏ"��]��y�ρ��LD-�����X[�j�ٍ���'_�!EJ�؍Iy�P޲����ʵg�wo�Z�l8����u���^��٘�:!��y��r�i���֟�<t�g�����V�KA'������6�2�G��K��<Q%Wm�}ޟ�x�ϻ�~�=w�$)7[���I�%Ze�}��Zd�C#��g��Q����C�!B������0���X=(h��Ҩ�V�"�Zuk��$®�)嘭�'��Ʌ�X��<Aq3���?��,u��)�Yg�vnj�v#�	!��x}��X4�Zyb���Bzy��^�S.<��BY1`�߿b#Fk�ی�ׯ�^��:�b}������{�����z&}��&}R��0�4(e#�5Ee�p@�����V�S�n��d�;�[��dي
c����ۯ�q����/���`"�����EB>ѓ?/k�*U���z���i
�ڙ|Y_)X<*T4H����`\.Y�4���S�,4wJ�g(y���SW���Qĸo1�0����}�^;54y��s��� @����&wO�4'�;���E�<c�*C�qq&V�е�������(���&��3#�����rm���d�`�j="9�vD>6�r�M/A]�Np��cܗڔxa����t��]n*� �+���["�Lt�X<?a�iB��C��Rق�d��MiW���?7��} v�
U����� ��q��d�j,([����C��K�PpU�@��W��B4�ͬ��f� ������}%�z�|co�%�-7w�3�����z�)|#���z%��{ŏ��n~�W>�*��Ȁ״9��[��%k�i���a<%�熀I�r����Kp�p"�y�:=*h��d�oKg�w9-̻g���ˎ��lz��s���l��fHW�\n��?�؍�o~���w#���?��)n���n�-O�:uyn,v���NؚtU!
>6����`p�ޗ����2�N���!:����(�=����,<�=+��yzF1�uw�}=��٘S�_�pftn7D�T�[Iv��v{�Oj�U�����ɤ�����0�1i�g��G	�W/,�!�|�M�lݛ����{�a؞q�qw�����m�#�vW������r��Wt�Z���¢�*��ȁ?��OQ��a�k(������Rr�����|��ND�3�����Ϫ������T�Y%�RHr�`��-��ƃ�����`Fˆ��%��	$��i96� �`|bA�g�fD W8�4�$���{d�'��΅�'b�k��b�U����[kX��,+��-6��������Ðz�Ӱ�siA�N�����e�� zf&��ؿ 3Z�`(
N�T��m�1mL��Bt_dY��6��ǁ}^�g�1q!��F��0o�Hq������/|v��2���+�ӈI�(��5P�j������yp��=C��qſ��Ĥ����G���7:t�%�`�9�x��.h�q��>�*�Р0'4b`� ��#*!�%y�77^7
4;�v��<X�h<��C1��gJ�|s��8s��r�>����G�ucJ`7F��AC���Ǻ\�h�>Q|�p�F���=i���m_��?w�P�E�h����W5:��0�4e�Y�v7F6�E��'����SM&�ϼ�0��^�ǅz��	;��-�Wȑ�'�I���Z.��� �wt眨`�����f������޽}j������mC_�>�}p-����N=县��;5�e���As���$����v�$�����UF�����*UZ�B5�7.y�+5@����,��,.E �I��ps�G�έ#7��.��mv���a�ipq������BݟWX���!fщ�N8P�Ѡ���c�i�>���>��������� ��o�����?���*�����G����'�왑,�ah}�m�Xh7����{dF�?C��@����:���D²��D��y�=�L6�g���V��ye��w����X�}��#L7o��4���+�����6�N�za�ݕb7sp6��Le�7>����)[}�[o�-�W*M��`��{��
�����<B0G����a�r>N���#��ןC&���e�3��-�,l_��ܸ�u�Jο^ d��Φ����b�׏�(���^������m�21�I�98-T0T��߰�:�$���7:~gH3�υ_hQJH�Ӭ�NU�X��%�m�ZӐ�f����&pdIW���-|��1#:y��7��t��[�(��B�ejx瞱y9nH������n�vb��6�������Y�+ۥ�@��9q���4�>����|�	|,�7�7�lV�Qy
��V�f|�_�O�|�M[_�d!+��I��ֿ2����+�k�)��i5
�%�i�H�B��p��<Sn��&��{cڴ>���}@�fgb��@��B�H���z+yR���cK	i�/�W���%ʐO��{��3�6^f������s���F���!��P��3�K�Y��8#�	1x��/��=Cq��&=����P��C�(B#�EW��
f6�vc�A�����9f�S��ʂ�l}�<��ȺXٵ����9����Ma�o��
ÃPO�u��!eg	�}"�Ƣ�;N�	!%h_�
8�<���̲a�+�|���Ys<l-���dZ{�8���m�M�Ġ�F�Ml��ATы��w��-������%�W���e�ģk�}z��C�M{�a8÷�J&P�#=�"ch���Ic1L0�x!��O}#����/ho��:�(&��H�)js	#J���/��ed!r<9^��"\�:k���>�6��D��]�O�-�g��q:m�R`}��gv1��� C�N�A�oj�n�Z�B ޥ���Y}$嬌o���ɕ� �c2w×���R�*�U^��/��nՐ��*#�<�N^���<:MI��8'���o�~{�[��������ް��ܓ���s:�c7`��C�	������+��|����sҘ�H։�kt1Z)f8�pb[/5~|����u����*���[`~�4��=� �y��mjWf�}�X����B��4Ҵa'|p���M�"�1���S���9)7�I|��F���^R�x���"����5�����W�Y��>��=���p�z@������u_�����i��,#5
f�=�����߽Ay���O�}t�u�ߛ���P4iM��<Fg
S�
�����e��oN�{y�*���h�H[Q�o%��[Ң��)0�!3���FR�V6��K�����-�����Ҭ�-�'VmL���ې!��yz��1]�	�}oh�<ٗ3w�����4��S�� ��ܫ5��pƆ�#3���0X8�������%m�	$d�آ���@�uԈ��3��к���T��N�f��ȞV�9��Y��ɍ�Qm`栭}`��A��q��!��3��=�Ep'���&P��>3�w��O�O�G��G��[��po!���p6nf�:Y���0���T�4d����޿{�m��c��û}�~�:���.�
Z�׺�:�u�9�k�q8Y�0[�&h���(�ܰ^�Y�P(a$v[^%7q̣��Ek!�����vO<I>�	E��ѷul��%j��9�������.D��6&���!Ltu�)2��Ǐ����}��}H�gWQ	Rgqʣ����>�ٲ���`����޿������޹�C���ݾ�9�\2Ac�i�x:E��Cx��7y���<���P̎/%gz3J���T��0Q�D'����%7;�wѵ`J�,�D��k��p�<�"��q7�9�aj�_Yx��$O�ps�s���a�RGy�g�%g���28�<���2�O����.�lz�o�B�"�T�缩F8�Gц�33j;d�����{��#ՂΩ�/L�� ����I�U	@�,�C-:�y�L��ϖ����y�D\zεt���۔<�#ܱ��ƭ�zg0P	;����^��p�F�vQ���:�ujFTl$8�"�k�pgE3n|m-M�o֟~��x]m���\�9�\}�0al̀{����%6ͧ&�^�T`c7�� j�[�����
��6Cݷ7$��&�8{c�{v�>�����j�ɓE#X%��^�qA�G?`m�^/�<q�90��mt�h4�N�ʪ�-N�X�9���t������NH��8�NT����c z�Q������Ă8�_�'����_=�����E��
*�4���5g�
(xݓ��T��^H�H	By���aP��h�Z�lG�Ոv����L�!�X=˩���t��5�l�h�����?�*�Dv����{�`xRo�-Ly����4p7��Ƶ�t�Q��ۂ�3:�jA����}�Ήu��s���I�=E��|�/�2hG�N�+�/Gf����
[]���@g��-�9{xk�=< �r����o]s��i�yb:`{ �m�Ĝ��\<�(�I���H��0������p�qlA1:o3�3�X+bDR0B�����I�w���0��Ȍ��Ó{aKp��;U��%���(����D�WEж7�HY`"������ZԿ&b#�>��)�-�2ڞ8gxui�y~`}�l1#T��^��^u����������0B�.7jFG|���G4���sim�}-�ky�=pR�i{�7��J�#��߯�؈��H��$��A8`�ܡ?�H��DoU	#D�b���[���@~��J ���e7�����g�Kpv^$�ɦʢ)V4�c������z���+��+y�n(Ƽ
:}�7����yF�v-��=B�����;�n���p�ݛ���π?4e��C#{ 8i1���:�i��c��#Q��M{=dq�@�[�&(N|�`a"w����96�NՑ��#[A?==��2#j���M�~�U�J*US�ΐ���x���T���\^pY	|Y	��xr�2���9��;��:GP[��� �-~{�'bkW����VϬ��L�������p��`%D־$�(Z3�s>�x��,�̵yТt�+��[c� r���Kx�H>9V�V*E��d���ب}c"�%J��|��y)X�r=Z2��?;����zW�[�]������ G�R�ݐ���{�0#z��0FҦ�x�)�*x�5�:���]�-q_a�g� #�d�p�hl�e!5��P��6%�i��4y��{���σ�#w(ͬ�Z���DuG�����<M��Qc{#�H2�SdWiw��a!�����l��ϤQ<PՈ��S��{��É!C�M_���0t��鑊� oQ�BKCz˲V0�2��L���	�V'?� F2G�8Hԗ��<�d�E��C43|� \0��Jm�:�[CM%#�dU τ7,����)��MyI�����j�Zq��mSgʱ��m��w�W5A��mK����:��ptA�Ul�k�]Fo���H:i92�'��(���>Oy��M�T�s���q�+��`�<x��@��IQ*;�<��!�!�v�i$���z�᧤�I�F[='�
���u(���9�������M���'g����̻g�-�o��x��"6�$�^[�L�	����g 6��+�������o�����^���eY�V�]"*�i�=�C���x_$�r��ॗ�h�ύH�#��K�b���3�b4<#�u.f�N�uh"i��D���mH�^�@�y����=d`=zΣ}	*�.厪�=��@'�2�ټk
�����]p�N�4Sx7G�8Wax��I�q���V�U��3X�\E%�l�-hpQ��6�
c���X~�s&#�Eb���	��N79	wD�F�u#�d���U/s�Ԩ
�W�5���Lj^\&�f���]�Kc���
�ӌ��n���T��;R&�n�Խ��x�H��!�N�1)F��R�#�Bh͵ḭ�%�P���8�[��#���4ȳR;(;�I���HN-
B�|������?0x�V&J�e/?�G��@�	��)@����h�������X����9X�yv���Jc�1�����i����2J��:�ʖ1ef~+)6�ؤG(/�v�����gc����/�i�4t�D2#}�R�<R�-�4Gخ��]�w^�i���M�SQ����7�g�yIj�jo�J����0�j�!u'�<�s�qH�C��\a�s����C�7��Ux.O������
*���7&b����3��l`wn߽��%�����Ql>-r�\A��~��S�}�(c�ߥ�g�d�S���u2a�-<����G����K�9��U	֜���-�*b	O�Y�$)���7�*d,P��DàmM訵R�y
�B��3��s�BR�mޤ�a�7�qg;�)	�Ф���(��	X4�-5��w���5Mم�x�HT�C��>�{3%)��>8�IQ�*�&�[A$1'�F�ĭޣ��7�Se����~`	��_��3C
���zr'�Ƴt���3�?���7/9c6������!+���2;��k�xW�R�h��]؝{A"�2숯-�<Ƣ��!	���$�FId�4ʲ1T��	�V�#��$��w�Jq���~D��ϖA��VO���S�>�<�2���4�@�|��]Ѧ��ww ��N3��R�1~Y��$ޤ-�f������C�I�L i��3����{xP�X)6p�fh�I#��܂���p��P�e���u%�[Tȵy �cԺ5�;�m���5��U])�k�=@	r�iD�xOS���$�3� ��S�4�C��hz�qǹ�o&��������P�^�?��(���qO�8�c���-�8T^	m�(b��?���b5^.jUn=C{�/����h�dr'���@t�x83*���: 4/���@+BF�8��	 լl�c$�!%�|��c-hR{O�Ak%9�'�39��!���}7�xː�4@�!���N��� �E8�(A�/�a��.��^ANsn�֎�Qy��[����;�p���B�����m��Y���J�<�%��ͳ�}�m����� �Q58սt�1�1Kg���8�����8�Q��2���)��$��r�vY����z�۩b��b�g)��yM*Q�����#�3c]tz�8l�^��)�����KƱZ���E4N�Vw�H2�a){%�+86��Ǎ������W�N�����B}�v�\�Z��DBx�~�IP�FM��Z���A��{�K������@� ���$�:NX����{C�&���9ZIU�^a�?�au��h/��cՂt`V
V{З
[*�$XMkU��A�z���}�� ճ�������?thB��@@Z�DNʁ����?��b7�J�"B��.$��x�4@���U,�!7����(9�qJ�%<��'u����I�ޗ�4�M�'{���n��ԾV,z��
�:JJ�jǁM����6�f��զ�yf�IoC$�tb&��l6[E�������&~'.����D&_�(�;��q7�,ȮdH�$�Ҙ
OU���^�u�0e�5��������5#I�dc�J����OO���׵�1!E��v0"Cs����n��#��4<�&C��:zE߷ɆCv��r#:�G�`�F¿6���~��`��Q����%R΄��d==��ޖ�)�=N����EY���>��|�>�?��!���v�lgL(a�M��J��x�+'`���քl�HeK�a2�A;02�+�H���Ƽ
`&���\.�L��q+���6Bq�C3�FR�t��j5�q��\�)����ݝ1�F5��*Y�Cq�&+�!��WC��B�c࢏�TV�#��z��^<
���Rq%�J́�i�<��E(Ӭ����rS����[�ҹ+�RcM*Y�O��<�<ĸ�@��6��'U�V�����k��������O<S��ږ�m�$B`H�Z��,����H�5d�����aY���;-�O�7�uO�^�����6��Q}��%
?4�0h��m�;��TK�̤o��%Ӣ3m:�{� ��C���Բ r��(��(@ˍ�G+�4�h��F V��=$���=ĎO���#T��a��3(A3�Cv-,�%J�[���%nM	N9@�ޑpF��i����n�� h�[�̼���GF��U-}����-��j&e�� �A�����0�����xH�8fì�T��ȸzB�8Q�AB�[��9S�t����T�觔?:E{���~��{�!��̆*a��"�- �,䏚73O�"g_^�d;,�X���v�Kȃ*>^�H>�JxGy>=�<S~K�=�6����Zp|s��<B/ �� �9�fԷԝ��������c�)��6FK��^�F5��A�2�%1��6��,T2��! ���b���&r�k8��vzc4���yX��TEKx��2yqv�� nA�=��k� ��(D�ׯ��?��B��@'�E���/1�G�֞�=#	�C��9F�D��	F�� (��l��L��Q4�SOf�'��|o�5���MWi8��rⳑ�Dɹ+��:YE�{��δ�׍�ajJ��nL2i�jj�{���5�1�����ݰ����Gvf�S�n(ڷ������{w=�$�Z�bH��Id�<��tC�N�(�|
C*��]Va��	*������}G�.�ą���F\��k���S��=1R��!A0�<����d�����P#Gr!w�ŧ�f�Sd�'ǝ6$�DAѤ"���l��Z4�ؤ��^�������X�v#�(#�F��U^u'�B����$��"c*O��j�8�:���C�� ���ѝ�ɮ����S%��^��%ճũg�a����~��D�I�sxB�<���sьi��k��`-��XDa�]�ЁG��&j��P� ƺ����V��v��|hNk�}evx�Ŕ*W�hS�herb�-*������h�&����բy2�ǘ�W=�����?�P�*�ݸ=c^"z[�⠇���ᗘ���W1�5$���Fz�7�G�a5xZ�Z��PJ�F�Ⱥ�p��df�B+��3lP�����恙껌�7�s�9�012�O@�>E+ZK�l���8��$�:�)^�� ��~��; jo��,A �B(��l{�t.����k�[f|��sy�6.�^�Dc
A���z��tW���k���d�:�^��v��|�Hn��	;G��c��l��5��WHә9�����E�$��Qk:��0FX/�L�򴭝�{k�/����GO�̱���� ('U���	��lTg!f���P��Ȧv^eա9��.n�!J
���,h �<��њ��DʖXC�ڿ����b��T���}��'����}��([�H���CKy�q�m�pf�Y�ʵ��	CzU'��B����R�f��
Iއ����h�� jeltR`������[��]s�X�A�;&��P��+U�A��W�BA?Ո�Af-H��Ha߄�:K���KO,�O��M@c;4M>�(�C3/.��Cg�	�5u�����������{����6y��p�Ka4��T��B��b�Y�į[�?.�s|�)��������k�x�(��感�ћBW���_���mI�1o�_u�_�$���͛�5[�Ki'2�!��7��p>��?�Ȏ4\K��Ʒ���-el#O$�7z�"�CUI�Y�X{��V�14�5�Fy,��EXG��2z���}�hG��=�k��� ��4�0x��ؕQG��W�20���6Щ��a�b��ځh���4���#y�à&}		Uj�C&6�v�l��(�PQ��	&h�"#(OZ���RS�B�>'����38��w�lBle��u����fQ8�2fs6�T��u��E�7�K`��9�U"?F�#�v�f�0�V��9K��f̈́��m%<�\jϮo����OȊda�?sQ�@����2���Y&�,��-�"U�s����ނ��Ʃ}ٝ��7�������v�L��?�P>���d��<M�`�~]=Awc����	��c-��� ,0M�NC�Tw�m�IS�f`��!6dx���� {��1��eKOk��B�qP�U6vi�~�}�PI�aǢoI��gE(>���kv�@�'�Z<Bu\G�|{!�֛B2�����3;(B�	�����zʋ��"�[`����A&�R��vm��V�s��7��Y���; *3�żj�����a�H�+�у�H/�B�Eo��|��*E�o�*[�'!+��ښ��Ւ0����*�.�fߟ}�3d�q��AL�8�q�!mgޫg�aD�`�5��s텈ak:x��l�;��8�m�z�u��~��~N#�Kl1w��I�<�v��ү0�ޙbY"
UN'�jFz�J��:�H#c�;��IB���m��E�U)8iU�ɕ����������]�u[�z�X�*̨�bx2麷&_�ᬩ�Xn�B��n�cxEZ�G�ֆ�X�Kt�;��&�B�ӳ��'m�ǽ ��\ST��ЈK�崧��HU�Dٺm�s��E1�	������hv*�IOlm�񬮁��+�sTC?�X��诬o��CZ��_�H�ܸP}�͓�N`[���1�FT�-���I��8������PÄ�AQ(�b�]ЉJ��Q�4�6$m�7|Ll�s¨c~|���!G��(��*�zk8��!�l����5x�4vu�n��L�Wf��1�Ps?�X]윆�|"�^�y�tj�n���9�{���HmM�Sb�2��\��}�l����'*S��ӲF��y���Lc�"y��Z��������0�7z�*���ƴE@t�:x��r�Tᗰ�Ȅ�@�:e�+��M#��j�<��h.8=+m.�O�)��N:n3͘`'Z/�����D���D� ��0�0$��I�$�F��da��ĳ�0��������|b#�=��R�����Z1]>6�� �+s��!զ(�- <*<� !�\ѫV�E��
��I�����uȠ ��KUіI7  ��IDATX�i���;l�y[l*y'�Pfpe$u�o�O0/f�Ϭ��}����M~z�c���e���,!���9ɩk�d d��"/�.$���qZeL�x:�I�5��~�t&֚k71D��A��	�')��u�t���Xɦk�b]HR9��E]�h��a
�^�=hs	OW����w��\D 4[L��֚����|��I&�o�y0�W���� q8S+֌�B~o-�U������=b3T�4,�`���zgZ�G��6e�E�PF�ɐ�W�c>y�w{wsj��+�Ѹ)ԑ'dX��m1�h�Cɾ;9ز�&��:��%�:��	��O� Rưr�6p�H`��-�s�t��g���,�qÚ:Ͷ]<��x��������M��&8A����&�`���!�P{���k۾=���%��Q�n��Ђճtze�٦��Au𾬋��񄐴�3����ɉ1�i"�'�D���G�1JhQ�|����;�q������1�u����$�qh���E$|�5R�*ML�T����HN��e?�.U4��B��yE1DJǵ���y�뚇?!�c�����S>/��+<5Js	?�']��^_�s��l`d4J�����u-rv����µ�9��lln��[���6*"���T���S�ǯ������s����5 ������䡆*��o@0�Ř��� ���֛����3V�.��%?S�\�����Ҳ��e�`�A&ë؅��Y��C�ϡ8h>PG��K��V>&ʓ���~�����C��ֲ�x��"co�R��� V�h\�2���C��Q(��?m�OJM�Wԛ�bÐ1� '��$2�s�;ٗ��J0d%�+�=ȳ��`OC�l6��-��F�&����I�B�s<S���ᴔ�����Fe��Y�����C�~��>��IG7v���zx�� @�p�9G3<;~ַ5����-_�7##i�#����Y��K��kp:O��v4��H�����o-�xKg��z�.��C�߾,�+�)�mM�
^,a�
7z]c��'�Ea�t�kX���@22�P�O��DDF�L}��m���������?����-O0�.�s�t�G���g����u�$1���<ٱ������P�F�s拶��b�{�ͤ/)��RTw�-�	}�a�����[���0ɶ1�O%�k�����Iy-��a�� �u���D�U�,��6S9j>��*�����fl�!�K���~������%F����sXn7z�p�2�)C�5�
w
%Hƻ|��2gC�0�g*�?;�ll�Z�����+ժTaT������E<���k8�Ґ.(��0q��8gba-��iH��J���%U�IF},ܭE�U,1����sx�)�T�F�")0�#�9����oL��?J
�%z=Ӡq��p��I*�t���c���q=*y��# �\� {4����2d.�m4��#Y��5�[�y��!lk�~����8yUC�Z�VB�W���ҷ0uc���`H��Bo��oƇ��6u������ZVǁ�#�����?h���@з�5z����68�H4y����.�ۭE@�p�<�HHi��_Z�<Ҟ*�p��"i��U6�ήI����5���}�/�a +��r�r>*1�	�]��� O�W��̓5����Ž�Oz3�/���U��u��0�`]/�gP���L�P���tM�PO>���-�pķW`ZBn��A ���M�a�杊� �]o�$k+��s�*7d���w\�-C\�p��1E�[a���֚������6��¿=d���e��~� ��
�ڈM%�+�,�0��$p��7��=���ū��B��O��Ao�煂�9D�;���s���-��_}L�0�}�γf�\k��;�u��qy8]��n�	���}RԾ;4�ԍ�9ᎎhf� c�m�N�2��u�>	˛G/�ņ^��K�7i�����H�	UG�2�m�*�v�S�y�7"�&��KV���n@�g�k��|�G�	3������ߧ}M]�����O?�N��^z�_�pb�<R���L̓�Õ�ɐ1�O�7�Bk����S��R�M^���q�k��=���D�_;�/��c����j܇�u�=�(��}T�����钺��~�hW*���g)ۍ�*�*`�|a��M�J+e�E� 5��~�]dH�4��8 )����YhZ�>4�p��	l�XJt�F�t�O��_�_�	}ޑImA#1��󔑓�r	�w�М���u�����S�2�gs�^y<\�؀2� RϨ�qxa4��r�C�q	CT��l�ǚڿW�=+�ҋ-OR�	�G����@=W������|]/t�j���(
�A�;��,�_)0����v���4�{~�\����Ό���~~��T��ӛG��"3�u.g��k�#������P��wnU{���5�k�;�f�D}fR����@x���;�i�XX��C���?��=������݉z�����),�m�ZfK�ݘB�BЏ�9����2_��1Ѥ9,`iz�����u��F�#�zuԳ�TB�xI�q��^���	�#T)�7-��v*w�:�N�$�駟=�8xu�]m��4�6֗�����׿��)W�"��F�:�������\e��)T�R�Ěf�>f��� XJm36�����"|� �V�#�4��>��w�F�*�\`��o�*��D� �
�v}��^�-.y ^3�Β�O��dz+m�GfX�gQ���p�*���uԈ�%44�Gz�`L�a����T�ދ����R�*��
#�O,���5덉R\H�����I�o��nkC����PZ�F�qh*�5�}}���ZJ$� �sp�ʻ.^����I����~{i�wO���Ș��12Cw{�	E�5�c��r�_+{-�5�j�������w��`1�2��7��Օ��F�0L��#�5և`����_����Ç��/n���/fK�pްQ�;�����������C���Z�$�x.�-7躙�����/y�Phnc�yl����y���}h�R��d@˟��^��K�a��X��	�^IC��yi.���ވ�9F�y
R���ׯ�a���z^��0C��<J3��e�C��OU�l�7��X�]x���M�3R�N�� ��^����܀���9��/7����]�,c�p��e%P��'����B�?)\-��K�]�~�Q��oYg=�1����eM����Rz�|+�LM�Qna@S��v�d�JIK����j򽷃�*c�Lxm�mG�/�'Qx���(�Ƃo=<�
�Zpd�[L_��A	n�XR�04�4J��>��'{6-�&e_"Yu��G��}�<{2����{=��(/UuYT>�C� A����*͸�8|��L��9;3��'j����;u&z��ռ�5�x7�c�x��}l��=��ĩ9L��~���K]�g�ӛ���a1!P�b��5�]DF��%��Ci��@�{�����P��U�҈�����GZ~,�u�����Z�zn����zߣ�xf��{��믿��Yϗ���/�/�y��_b�fVk ��99���~����Jr��a�����waM�L6������`'9U�D��l1�^#8a|��XsFï����w�֢0�Sh�<Ю�P�$�њ�g��]�����ſ�߆n�|J�ŦvbȍF���zl+�]/'�F�Z�������U����r�"�%~c8Z˔�Qm@�&%%}ٳ����>3��s-o��ꞡHT���\"lUqȫ>�HBs���0�K������j���z3�v���w����j$7S%��ئ�ac��q�c�i�&ܰE�N������D��,9N�ϕ�S~��-P[Ϗ�<�2�`N���P���k�-d�����kTP��I�G��u{����G++W����ٲ�\��a���k3�|U���0m~��Qdq�қ�н⺃(4��0�=�M�Rm�Lx�XU��H�SPVx��	~c�&�^����;;]^����^=%/]���F3lϰ����g7&V}d�����C�8v}����������w����F���mc�P=J���0>I�8$��pH֬�`d)����	�8�a��kT�}ߤXH��z�^�7�x�fc`��\l|�hH�G��&}�h���T�l��ӧO����ϝi|��э)B3`px�$ԛ�:����<+4DR���������?�I�+E�+װR�����K��MKt��p��e�g(��F��`7�-ɛ�\�?���G5��0���@l��q����~�:����?��%-Դ�s��kH��7��@M�"���K��"b�鑣*i	O��±T�M0G⠕;kk�<Q�u_��q�	�R������5���u�|�("�p�H��֋㵞Trk+X5�[������������e�SVӍ��yD�!�G���!SH6��GZ!p���;���.B
�?��Y�j��9���O��=�D-�f�4�=Rm���	��O���������o� �bt����]_v�?�6z�jG!��hS޿k>��D:5�`ߓ� �c�\5��Mrj�Ka�=��G���q��y��w3Z��ԖLPr�6�_��78Fy2�b!ݗ�����fs�H��j�6i1�Ka|;�G;&$������)�ky����W���PRN^�LOf���¸ps�!E���z9#��]�Bo����i&� ���G=��x
~&��%�ٟ��H�6t
�QR��\,�6B�'?�bnm�?=��6���(&����}���������d/K�(J8�QucQ�5-���нF�}�d��z���1} ����5hp6f�/��ze�9E�asCEC�?�W6>���԰��v��e{6;�?�Ǻ��ʵ)#)#�i�#�:�2R��?S�:���ϗ�.�v��1��2�U�rp��c@I����ռ{�#M���_={6I�z��î����mHi��*�7a������Ÿ�g��%�B��W
n���뿹�[`�^�9e�E_,܈�E�EUI������~>�r��(�˵$�m_D��ϕS5��i!�K�D� �lk� ��&c0�H@�QU�*�L�h f'�iM¨a���>���0��H�m#:������'=zMvm��|���>v�싿���/�^���+������x�dH�^�(��Ңe3��4�g����1��ȼ�� �	�k�2Tz��S�^jYݗ+=��d=����8E�s$���!<-
-�f0ͥ������땉�[%��~{+��^��u��(Eϯл���xE��`{�׷��y�O�����k���{sL��Vѧ&M�L�&��=������m|��Lv�i���:���N�5�~-Ga������� bm�Vig_�!�a	"x�ͯ���r0����`T��}�(/t[	�3����ڊ�ꆷ���^.t����M]��$��r9}utT}М��C�<�e�0�K�$|� yHCTGܖV�d���L����@��:�z0�D�����6ڀdr�Q�3H��B!��3���{�q�xo?.=�-��֘p���-T�ά�u��}j�݈Z+c��jr�H=����3� �Оg��&��D9RWό�~�ʡ3ͯ��Q�}Q�D��M�ߖ�{xs/�|�Y��+*p)l�^׆��g�0�;�t��%t��ل5�����a��D�V����F�VOgMRJ$��n�W��"�%� ���Q�\cy��.��J����n���˯�4H{5�@{4�J�g}�Y"���8���Q�7M��f�:g��-^��rhu�E�� ]��j�l^��Q{�ʧ���y.9.�dg���86F��U�﵃�����W�L�ފjx���7 *��{ ���Di�k@�J�����;b<с���3�����yH���P51y�N��>�!�	>�d�3��F�z7dcJ�-�HiFq�����;x���%�`�GzѼNYK��WL�M�1��&E�6l�~f���9Z?� K���oϬ<7Ǔ����*���<���fp�v��g������$~��O�{V�^<#M/��M��f�����/����'ь^e� �c���:�gay����:ƼO��_��/�+��g��&�!z#f��f�(�Vx�ߞ!�}y}�'o�����Ȣ���-�7��w����%�4�`(Rq�_�D�_y@���Zn�4���/~(��g�9h>nh�]���,���J1{$<q���Yy��0���K�A�ͮ[ʊפ��
����xeh������x�v�@L��<��m�Gm�)ǸO��k�A1J��phݘ1��[�.�A��):���3��%�?����^�B��������:_��߽�"l"��ipC���#[���`�M	�em^u�n��M告:h���rISw��#���=����Z�iu��]x>��k�d�غ����@�q��\��V���� �hQR^���]�,~?$�������"�ᚼ
UH��B�ֻz%���[HB��f*ʈ:#���#���U솰E��C�Ps%ff������B���l��R�kF�J�f�R���Je!�ί���;Q�⋝���y���gFv��+K�+��v���M��)��%.����no�}���EHףc*�k֍�#D�rTu�J
����^x���~��eU���y�9 �W�"�EGC�}�̯�53�J��>7W�A�	q��kO�0K� P�A��i�������Bs�x����y%�P��P5��mu���{֚ծg�{�)���D�a�E�E4j�\ғ��󢌗[V*0U���l��-��2��Ψ~���]�[��G/��H`�SW��?FB���bu8��������ҠNA�Z���=�\��sE_��\�����)f��=��RT��^S��ڔ�<�y�£�x+޶�N�d;�?���OM�<̓�K ���S��5���� a�虡��ױ��2����\�%��ၭ����b�F%N�pf)���"����i|��!��Ub)(�}p������1��{m�AM��[�������#-�G֢II���@O�젇	����tf�
�a�,��c$�������@!�g��a]f�	���8H�~
�����Z!5o�ڲk��K����%VJF��h�w^��*�9�%0�tK�J�9�nG*�	r9����%��@�q|�_L���(!��u,��,`��nٜ��O�(��>sf����(=���p�k������NB�i�o:�8�v��o��D�U}����⤩�8�R��sO��Pw��b�ѕ2��h����
��)k�O�\�2�[ܾo����ԝt�frJG���A~`O(�|�����qnC�w�a�a5F�V��hk�s�B(� Q̄��{)��j�lۖ���8M@�^�9��8�|�Bi�w[�
���.�Ր�[��T,����ܠ�ْ�^2�RwOc�Y�Z�ը��Sփ?��8�%�GC��gS)fXb���B�+�V㒅
��9��U��Ͼm�e��"��Yj�HS��{&�	%�	9[�/>9�f�،93��p�1�(K[39���[��4O�Dt�����6�ڸ�Xu��#�^vF�U� �i�g;M���V���+��9sb\ ]��4$�K�Ģz�o��k��Z1�=Ӕ�p��Z��A4��Ϝ^e����H�a���@^E͠��X�q�K'�,�2���QB(�����:�J�vC�ғ��������Ə���q Ӌ��k�R�H&x����y���iM�mv]��-��M�� ]*�Vd����u�j3���}�H�k��� LvZ?>2��jMQ
��Ή[�jt���Voy�(�&#�%�'��9�I��O�u_]~ϵ�ke�4��vǊ����K�	�FG�͟�Θ�v��W��&D��밐�
�k��eQd7OYJ�_�c<Q!輨ĒA�E� �$z�	�V}>{�C���~��Vf�{z���'�w��;<�G�*S��[��i��ѷ���S쯚?�s�%�j�z94�kG��� L[�8��;3s�R:�L�����/ѝ"<qFsF�b�NI1Wv�5��
(~�~�%M�&%��^K�����rE����^��m�v�1H�L��X'�H�4?����<ȉ��v����}�XB���6�clȊ��{��7��Ĥ����~>^���^s��p��!�¼�Fib�1�4�<�&�`&�����癉H����n	�>j��#X��t��:�Nćט�m�U:7���������<;�Nl�W�w=�d��Kcv����id��F,V�@�z)���HF��DWQzt34b`�+�E�����{Y�H��m�G2"l>�aa �����a��\I�fе���TIǳf��xk����I\���A�G�-�kK��]RnP�}�p\�>Q@&���5��������Q��:;:pu�I#a�U�M���ɨ�mm:���y��������
�1�)�7&r-
s�Cd�%A�Mp�][�����X�V\iv��ɱ/��g�z(��[4زMm!��CM���̪F����d�i CC�����nz.i8�ؚ���G�?K؎�{��G*�سm�_��X%�G՞�x�wϬ�>%~Dϲ*�(�o��񊗷��Og�������Y�8���3�	%��[�O��`����.K,kX��t�u�L�n\Nx����N�Ff
�bl]c�(<Jݣ_��\�Lu}m���� ����)ȡzy��J����N�ߝk� 	�d$����J�f�b��r<���|E����z�����)������D����Ycoz��
�i���՘�NY�G�q}
��E<�9���R!�g�i t�ߧ
܅�ԓ��R����DM�3�Z�u�q
���Y{�*���L����� 
��H�NG��o��йx||�Cv@�<��Z/��ER=�;���)�ڨ_>�}��������UDl��A�yx~H��G�L�����2߲�5� %_�m��n'��yT<L���Gc9�	���Pt��b����\��Sb��v� ^����W���S������"2��3e��N%X�.G� I쁈����c0=V��&X�y��Ku"���n����E(�]WK(%� N�}s�u�0L�k�y�<�J75]��tְ/���wWrŗ=z��F=�e�#���6�0���B�Հo[?&?��s��g|�{��ʒ�:_�o�9������ׇ����w~��g�\3n�%�>�/���q�8؄҃i�%�����)����X'eJ��[z�����`ֿ���u������F�p�������r��z�6��4�������gBQ�S�pc�}�m�}"d�P �w�g�tv�ѭ�����G7+ѵ��k9�'������"㋃�Sge=1�$+oA�pp����p��T4B��%:b�Sn`?y�,|șUD��d2K�pz�'�����dx����:��w*N�rё�~��V���������g�����}��'�PO�m��n�$ʾ[�n)������O���4�����:z`m�X�8p2t�xVz�Bu�Z�ў9�>�ث!���	+��Y�b�2˙���c���ʘf��L��`�3m��QB!p�4�����Cf��I>E_�{%���n	u#�ε *_�����Gf�o�>���1ƭiT�T�o��Ӊ��I���#t�L���?h�������G�r���� v��ri[��-��N���ƫr����!Ґ��ф�&UPϣv!�� �j�b����h�3��"��p��L��/��ɲ1Oh�-�"XF�*Ғ�r�y
�N�`hk��'�����Қ���B�����tcy�N���=y\��d�MC����*��0���%/!m�c	⟀u5%yZ�B1��� �2'&�.A(�M�kA0��B(+'���yv!�o��YG�µ{|̦hØ�=�+�����X�dA���-�M��e󨓼-��tHZz?�1���72���%��b�������px�Ej+B ��~�g�D��<Kz���g�n�q��{�����"1ha��̓Jx��G6�4��D0ڀ��|#�V{��s+I�i�}Vq�a����4E�DF�&|}��R� 8󠓟<��G-zC%8O����	����٘�uU�ގ��W�Ƒ��z�P�X
A"�P�d�{`�W�^��vO��y��{8^���y�n_,�`u��;�Eg��d6C��1eN�+�I�!��d˚Yx�0mJ�ʾ�^^�7�,4N�ĭB>���� ȕ7C��m#�b��L��4��Չ�M(��Q5S��(�[8YcTH�x*�'8�i�2#�p�+��D� ��D��� �Ao��Nb�L�W>M �[X�NI���iOz0�?Dj�8 nx���"�L�@R���(-�\�5�(0��{�&W�1Q9��Z;,؍ắ [?��D*�e��_��՚��'��uINȀ��m��ck��"9E����a��Q*����4J��FQ��z0P:���9��Q�]in<#�[��Fz�T1�3��d��=�Z��-9���T����@R�o�b�ʪa=�~���]
�����U�Ȳ<���n����
r�#�n�E�X�)��q(���v�R
3����?
��+}�6�۽I����gci��=�8�e�Cz��H�A�ˤ/I��u�`�p�v��@��0�cd�e*OpݶX�
��@FĿ�\�7s���	T�NWK��{�9�~o�Ǧ`�/�*��&e�;6��q<��	E���&)Wʑ�yZ�6�f����]��p��I�F�O��X��gT�",ϭwC�y��5=�X?v�=Jj�N���P��.
]�Ů�Қ4���צ�S7h=$e���y� ��H�� ���]ԧLؑ28�k+��V���\�5$`��Ud��h2�|eBi�k>n���l&L~W�\�?E����^��B;�ʻ"�DkpE[W��E�=�w���x�5 ���6F+ј��e���m��w��y���
��nأ��j�m�G�Y����a���x��Zmas����U�#+2Z�yMYs��}�ó��pT�Q�a�ڽ��H�A^���G1�ū��]�Ji���o}榋�~���g!�yzO�B��	?��'� ��<tk�e���H���np=���r�k�D�I��w��*.���=�,8�+Ac�&{�\������
����,�K#W��� �Ry�f�
 �޼?O}x�SRV�}϶�#+EfNl�@��>29D(�Q|�&�*�}��������$�
K�r%g&�G��{㵼O%��� �b(UQX��z_HL*�0��r0�v���8^;kK�yB#=J%�4g$3�}���^0�����w�W�PPcZ�������������t��VEj�5�Ͼ�o��&����U����R�"��z����Q��Ǻ�ٿZp�g��G?�F��[eõ	�/��G�oٳ�O��F{�U�\b�Xw_0��He_�����dx�ln�PQQ�O�62�epʦ4,eh'���
o�V_ؤJ�׾OlKb����BJ7�� C�F��J\ś�:�-�(*��(+F�ڽ7ڪ7:7NXTSRO�f��+~�>�B�H���$���Q##�k
�D(�{��f���I�Q�c!��c-�
z�2��s=���rO�AW	�Ŀ��g�CR��)ֈ�>g�����`Հ�Ƭ�+�H�d��W�47�dD
�5>ֈc��с�з�I=8T�%o����J���!�-i�[�����Z���=�sd�3V
RY��f�jFH��^^��:��5^46�W`Wn���#;p8'����{C:�ŕFT�?�u[|7�mWV/A�U�Mb�q�K�])�B���Y�P�YU�,���ޘ� P7|:�eZ;d�����]�T�B�W��
+ܟL� �F-��6�-'�o�rt��AAG2�f���5c�$�/��U���+j,���J�Na�Ě���<���k����m��7*���1*�&��J$d��/��#�{=���M^<�C�.�^�����s9)D?��m��jR�
�b�ci}r�#�t�\�S�0E������KF.�ےc��%�Gz���}�{��{=;P�A�JN0�1�{��[[��Ҏ'�T�T�Heü�˓E�B0J�ײv*OɳB��!"�nWBz��BgxJ��ʊ-	�g��!mMsro\��������N�!���z<�+6r����!�&R,=ڠ0-���K�J��?��IZ��k�2r��V°hLඖ$��56�}y�(7�D�V�0(٤���b6�A�\�F�[aP>�.��$�ɘ��|�%�6��
3uǶF9��W	��t����w�������Q�1��;
��;�,q��͝��L�lM�Sz�%�tZ�m�e�������Z[��Gn�|V{�U=�d�x���2������BG$�Svo|�1�Keg� ��T+��K�
�|�v��_��?��ڢ�iO��[����2�����L9Ӏ�~V26��S_�~V�h[5�!���H��16c�.f3@��r��&�+T�3�9�IkI� �qJ��Rѧ�0tS�y+ޟ����Pe��5���?�!6��	���	\ɛh>��8D�i�j�4���6&l6f5I��A��c\/)[�=[ve����vO���K�CL���-��ʲ6b��ۿ�T���^[����8\���6DS�����W9����0#��y���q���jk�|>���� ��O���L8%wQ�p�~'����t�9'��Y��dUG�	_[t���m/ܿ�N��n)8y��s��@�!���%+H�
��4��,<��T� �?	�c���=�w�KMؕ�մ�/7��ϕ�x�㛏U��]�1��\+n��VA��s%#����y�EJ�c*���yJX��$mD�U󥹚X5&ÿ4�<�C�VM�o(K��FaH3�;�������+O�,Fҹ�Z�~*��|1t���Z�׹E��D��$t-~�͘�3�>�{)����2�20��̀��[ԏ��X{[�m0��BZ��T?<
>[�W� %Ɛ͇R9�~�n8uu��u=�d�mOz�,};SD�=<��@������ocs�ʦ��q/�3UC��7̌�\��@����>���X���Z+/Q85���J��D�G�Y�Wx[�Ű�nJ�}|���<�շ~�{&�Z1�Ca4����ш�0҈�w���W�Z:���[w~埱<Q�x����c썭 ���p���������.�/�A$s�
�]�F��y���g֭�[�	%���Ys�T� j�����?�QXm-m��M�+�ȯ?	�7�������t�w�R��x��FeH�������xc��0���{�)����9yV�v�Z\>�ŐЁ<�Ɠ8-�a��)����{�%aW �X���hl�e�P+��|��9���=�D�?�c��·�D=�1u#�O����VH����p^�{��*��)�#{�Yb�eL-�{=����W#�G����Hc,�2��%Z��p&O&��:XQ:�yP�PHj[�!������h�^��gT;�AQ;��a��H��Z҃�i���Q��c�W1��h�RR�9��+?gb_��!�nI��\~�uam�5{��RyoJ���M=v���ɾF��	,��JD4j�[�YN��, D�T!o)=� ҅O�P/�M��h�Г����iz�%���^'.J����5��sEH~�N�or��X���Ky��=�,�*[�����J��<��縁8)���U�#�v�rduT��%���㖷�wo��H��X�v�Mkഩ���4b� �d.��שM}���8��/V������l�޲��/���/�ևxh�e�?V}v|��Q́�aS�[x��q�%�kO�䦸?�����(�?�_�"t�P6<�e�씚������Ȍ�` 4Q��Č���Z���G�P�ʁL<��'����"�����#
A���;��5������d��<@$]�:�ש#�5�U`]I���Ű�������4����o5��{[��.�?w�1/�~�܅�p(��K�#��S���AL�����Z�O�\�s��們fH��x UYHj�%F| Nh"kO��P����c�w-�s�n��v��m�E������y�s)Գ���M�S�ZJ�	:�,fW��8(�1È�g��]/�i{��%0�m:`*:��kD�*�)N��f�%�a�����B}]�B� ���V�hn�=L����Y�j��|P[@�b���9�c��T�i���z���^۰��m��l��fK��PQ�����dٖR�ڷ�mM��s�jM	g��g��w̏_�*�`>*C��C�ND�&v�[�62L�;{�q�1�z/���#���y��IN<Ķ��h�3"!��	�5��֩_�!�jwT9"�!�G�V!�*�T:��G�v0����oV���Y�R9&��$�'�>��E�fj����<p-*��g��[��+���9)��w:UD�͌��*�%ޮ��:ΧbH/Njwל�峲�]��ĄZ;jX��0���,�[��3L9`��.��k���<�8k)a�'��@�-F�qÑ�d��[�90��Dg7CH����Λw7fkR�&��*������zi'.����/O�~�=7��ǌ�8��uid��p���j2�-���]�fs�ݐ��J�x��Z���-��*���V�#�`y�7���V��=�%���R�l�ֽ�95�kNQQۀ��.fn��`�jV���59��%L�V6S�	�6�=E�ys��fz�����	�Zz�G"���XK��Ęסx�CJ�+hF��v��Ġ�[�f�3�ͻ�;���,A�Sb�M���BJ�^JI�;�q�#��l�)!�`��X��O��������5�.�	g<�%��`e������Nʃ3�'.����7��!���Ki��,��!6��@�GY;��r��-��'\�yp�$f*����6b,�[���]K;[�*�a��eɊ�~TfOC���OLS�_x�%�����I�W�<� 6y��s�ic�����mE�QW?x�a�$�+nz�c(� �3��/��$����s�x<(���z�7�ÍS��B7e^}-Y����a�y?PU���5�|��h�3�v��R�ul xˌ��4���l�e�QNzu��z�)�����j��V~�(uuouagw4\�T��ҹe�x��iD�labɹQ���}|h+3���v���s'�S����x\�n��������L�̑p��u
�O�ȼ�J��	%���	���CP1�.�?�EA[�bZ�מWa���u�By|@��j,����hd���ᾮ�>�*a<�K��l���9c��]ɧ����g_�6(ޘ�m��k�ɓ�6�?�p�p���)�=���Z�#mxy���+�SW�b��0|�Yn���gW���p��S���ٮ/5���6��a!�p.jnȃ|S��W�߳)՘@���u�TE�Q��ͤ�����bHÓ�ސ!Sh|���+���M��(�hdZ��]�ߪQs.����0�1؏d&���NkLR��Pޛ���Z���O�R`��S}L��hZi%R+2���D\ч�V#1����<M�˓6��&	"[�gF�g�pJ�˼��l��g��s�L}��cd}� 鱬�P+�A�f�C�-+�����!	5O�9[2�0�������j�+���ď�֖�ze6x�SQ^NJQ�'x�-V$�VЄ`_�Z�լ{?{cD�<od��T5-J�����E�+�1H������I[J3�6u,U�0@�r�HU�Y��3��b�Ʀ��C#
u	MF��K?l̑���f�%F�;���Wb<����Rh��k�7��$n���2����Xɫ��QRJNX��IC-.י��ƃA��Z=$������Y��LJ���Ǿ,\o���co��-1�]�9m,����-�v���H�J^���fFPՕ�¼��Io���o�JR�=u9,a�YN����w���n�Z����{�D�d�_uy"Ai圧��F�2�je�I�R�q\�r�����&l���1��u�Vi�s��0�O�a��Z6׼!���h�W�*��'�4���!����FU�oj���їB��ͅ���	A`��K~a�3R�P6Oy��UY�ۺm>���?Hhl��;�����x���d�Y�U'�xP��2*ԩڶ�1��w�A�%~YD [�ыW�h"[Y	��EkYi��}wy��*a}g�j�Z@O��f9+Jh�\8ĩ��{n��{#� ����T��:���C��,IY�������	L�U�
��L�Ł2NGY׮�[r�"��{�/��2���X)Ό|�a�A�\وǽ�!Z�܋9�r���qC��R��.�Z�ɃG��d����l������ܨ���-�}_�1�P�)K���
����!E)��n��U����p��[\�Q�� �[N��(Ƒ�e���cl��%���I����\���)Љ56V�N'�hT[�F�;sA��.jA�
�zʓ�,`���]=Pvu0�+�w��2p:H�	8��`ȗ�A/�`�y�jn�����KY�U�njl��x�z�
��n���Nb�W���/nEP�E����3h�vMo�^�D-�{8x�����!���t�OF��2ێF�!��#B�����в��݆�a�Vv�Uģ�Ud�{t޽F�.�s�ͤs�ۘ��"�ۺXC\F0K�F!�?��$��n�oES�Ác�<����j�TlT�K���C����DZE�-���g`%��[���7W���K[gf�#�Z5p��x&ws�����u��Mc �$�2A��M�����F�w���n�rS�DϒZ�����0�y���?�7a���O-�<�v1��_u=���������u5L��wLjddP�L�	�j���4���!�/��*~����/�E�Wk���񹃒;iH3��a�8���OZ���F������~�����X{�����z1��N���V�/����G��/o��)x�UW��yL���!\mb�"g����p@��d҅��Z��	>��n���\ә��u"Ｓ.Q���o�jW�T�!۳�S]ac��A�l}sJO����FBF1�~Y=��k�WC
�
k��Q��b��O�yl\�Am�ӗ��r���A���D	�(P�V^{-;�����5m�U�;�B� �u���ǅ��m�_Ƕ�k��'�����%=��H&PLX�	m��].K��Q�T�e�
�{Q�[&���U��s��,И�g^:[Ġl�1��cN���V����7�u�Uꖌ�P��@W"p�ҋ�F%:Q��T7p��Aj:��Hw�G|H�4
Ð��X�0���RZ��܌�z�3�y�Y��)>���#��CQ�훸�\��Lw 6�}��A�5���;��%B�I8�i�=u>�r�Ciɽܢ�G�tF��a�����m���|��ѐPJ��B�;�P)G�$������sG�����|N��?2RG�?�ߊGş��`+I�zў���VfW���A������6҉'m=�e�8"�r�)��a,i���~ҙ�x2�Sn��B�T����Z+�C�c6���n���4��������A�D޿p˲��0���Q�q��� ��=<����*���r��f�|?6����-�ؚ�Ҥ�e�����h2t�2*8 >8������X����P+k?�_���Ua�\�e�5zC��s�4��@����k�U�5�w��[+��tB�pL&��mwi@hM����|::��m�o:f�q��>pZ����ɛ-{6��h'�q+y����'����!������u%&�
��* �)�'Ӗ�`�E��n[��)$ת҂��~>��|�ѵ��>�.�AR2*|7�I��b-Ƴ\*2'�0
e!�^���j��o��;J�ޓpc�|O2��k�i�I���Ɔo�:�X�,�x�5f�HB!���6$f�&��0N�ʩ�b/u�9P���¬��L��`�������Wd��Z.�b u���	ȉ�)��vwM��H��A�,����ǁ�ʿ�!��9��y���<����C��1�L<�8w��`���0��6t�H!����ض���I�8�T�Y��C�	�-?:"�!���:0���+y�	rY���#~��a�!�{o�6�k�������:t�aԛ�7B�#y��0��*��� ի�=	+Ȱrb�O}1�&ߥ6Q�|��߭�79z��a�O{8�n%^�we�OzD)d�gik� �:8�[����7�{n�$�䡈z� I&# �8no�e��P�����}T5��[��PC4Пr-t%�������e� ��]��eN���������쿟O��!>ϝ�e���!��mˆl߽�{��xώu���5���������w���ǘ��A� ?[��2-p�ko8~8G�����ݱ$7��{Dfr�K��F��>����y���nI���B2��xa0�H�J�3!e����;0 ��}6���s#�g��If�A`JsSC2	D���o�W�8�?0G���������������#��:H�.����T�N�8)Y-��]i�y6����DL�ս����lύ�O=A�E�=�@��*��t	EzeD���VP��#��#���	�e��MKM0"s.�!� ���[V�={��	0�e-���T1�e�*�����k���T��$8F��Ze��ʫ�]��y�$3�]ɓ�I��M�X�K��K�3Ct,��;[%R$-���&Q�v����@��[ey�آ継�3�D����tx�ͼ���E1�Ϻ����o�i�oBg�"t%<��Z��M�`�3w#ބSdP���C�?��KR�.k����6�=�����(��O�<�r��^0���&�0�q���,�JB��6�Z�h�Z�^VK|f����*��X�q"Vb#�E��0�}��zX�2�.�5s(׏��$Bu�زY1�q��0�P�U�И���Y^E-K���󭊵/q>=o��c�oV�߸V���d�9D�3��,����P5�|��rtj�̾UJ*vuX�r!3%�b�}�L��l����T��A�E�����2�!~���eֵ��C���|��Ϧ{M�ϤK\���`�s՝S=�d����ƞ��y	٨5���Q_$�KI'��Q��f-�?h�0e�U����G[��U�{��<_��[�����?�g��4��]O�բ�ruE����ݖ���e)�6y�ZM���,)LR�����^AQ�N#U�f�XU2�W�4��;�IQ^*Ҟ�R�#��CR ��RΗ���Ÿ���<K̍��Zhn��be��4�!;-B*��|*}%"�&v�W�A�N��d�%>��\�q������O�^��V��������-
F�"dRF��d7Q��]L:�-�u�"���F�(�r�k�F��p"��T%�}�+���4����{�������S��;�w4��q4���US��,�eȹ	�R�rl�M�tk%.���Z*c�EȮ��<�3��5�hX*l=e�*Ӎ|9$��^ݎ9>X�LL%Z�.W�{(�@�a�ge�R�&u��!�XJukd����f>��.��
�O���&�����Gv�R�1fI�c���ׇ��%:�l�(�z���m�h�[wC��ZD�=������Dy܅��V�؞w쑜3D��@d����,�F��u1N�I���҆;؋�9?�V;eii�h�xo�eI�8d�J��"�2�L�+�����]�཭�-�:Z���sYE�Z3�{(8 ��0U�ԳL���|�ޒ;[�RWK/t�+ġ�n~�X_��*$T]�P����BU-�|��/#�ò'�P=��2�Q���j��#n��y�ʲ��K7��F*6*sc��%��B��v/���ܽ��<���_#�+Y�������WE��{�ZA5�h���C	X�]� �(�\���T⾠����6c�O�y+.��Ń��q���L/����i�X��%3�Sco��o�DV�W�����c��͑hWLV}I�=n��Ҹ��!�a�%����H�m���$7�n4�V����d��*�?�U���b��:��qR�֔�c��i��	��Z��ZG>� ](D�� ����8�U�p���	@���Kσ�wy�Ճ5�h�l3yY����y/�Z[��*����:�ׄjK���7P.z{4�Q��G2C���Zl����H��y��ǫa�]4�2|޴�J�nN��]bq�+
5��+�y~Hڪzy�e��g�)s��Z.�]¥�%b��z���m,[��7c�]J鬺ڸ�E���{8f�D�S�_O7}�b�lPT�c��ŎE��rO�ɺ ��D(g��Ʃ��B"�K�m��?Zt��A�ne���|ΡW#��F��D1\�����P|ٻ��R���M������J�ֿ��$�=��#/m��_+)U�E)d�Z���W�-��p�U.�� ]��>?�P������N@�7kx^6 `�2�ZPӸEL�ҍ2]6��4�3� �*��Eq��v_Ch(o�DpϾ5���9��銪�+�x��9	4U�eCo-�f���H+Р���%u*N�|.��	����9���ڕ5�֏��v.��~Y�Y|O� �3D��$�朝�[��&%t����T��בi*�HP����ޔ�]��"��oj�"����Kר��
�p�-V���O����Z�R͡���h�8g����iΡ�>F���b�Ҟ��2E_њ<�&�R�]�Wʮһ�$�e(��]S���h�D�9�j�Qkb��k���UO���x�2�آ���|u�7�$�J10t-k��MM�x��E���F��s��@��	���ƺ��wB��VV�qh���d=A�?o�g�*��Ik���dGPC/���!j�U�u���֘����"=�c�ɗkT�ӶU)�}��k���[�h�~��ʲm�^��Q�k�h��)%P8a����#7@���2^4�ə�k�Ak�\����2��ӵ����Jݚ���~RZ//�U��n}���aN%;gV_�]�a5WT~�2u��v �!�y�b��L%�
Z���-�J.�gm�s�E��U�dU4Cue�
F���狢k�|^���_����ĳt?�1�i�shM�zU�EE�g�}�b����М�D�e>�N4%��"�4"Ul H��Х���C~8c��$n�ҰҘ��H��4XBY�L�*��˸l��񔆽����k�$�w���I)fٖ�UԄ>Z�Ֆ������n����ַ�AP���z�!�����u&|�Z�,��MZ��OO�Ae*W���������v^�N�Xc� M�y�*�m=y��\�^�B^�gK�lE����������7�H�ˮ=�
�޴ٚZ&JF����U�Rs�U,99�Uiuz��HA\��,2{�]�D��7X��,��g)r�y^��q�^����؋�A+�N2y���u��+�OV��X2�4�b��_dP+J,�2�Gu�ɲ�-����רwݯք<��dJEl��(�f�=ǹK68�&Os�|��zn�<q�zN�2��H�e�� X^e��$��Mx��>OR���,[��e�*� NT+h��'򊂰C�%Kd��l䃪�hy�:��.~��m�
��׋�M��ed���FGuS����Vo��[n	�$%:�,Ua}j�_}�9+Q��5GA�)
��F)й��2�>��(6%��K�a�Yv$�3dU_ם���D3��Z���d���"��N���_޻X�ӥ��~���KgG3��6�<��F��R�Ȧ�Q�*��F��Nz&^�VW���_�hYkFH��0!��;���ͽo�M-e܌R�Lq�ԫs\N�{��\��^�x�)_�`v_W�KI�����^̓��ǋ�}��J�ni�"�W�����ō�U���Hx
�7�)����h�j�^3�}���1�����~z���k��ŭ�F%�f3?��YP}gG���﷔���_6ISj��%�%��EFe��u�=8�M;�T�<��w�ie� qn_ ������kb�m�1�]�ޣVjqȍ��yTM�My�B�1�K����V��~�z�R��t}C��P�j=U�J�(����ͽ\�W�/�!�4d*��#JW���e�
$�2�K����z��ac��fy92z�L���U#A�:��G��k-�q��?k���4�������ȉֵ����FS�������.-���I7d�cp��Ja�X^�������R�U��}�x�%�YZq��ma1�0��/I�I7��|~{�t�+���x�j+���AB~מ@xEq���sҷ���NOw0�z^1׎{ma��u�U^^��ҥ�ʽ�Q�#�Š���_W�yi�QK$��ߠ�Q���ҽ祐Li �2FGɥZjۄ������[��eL�Ja�w�9x�=�ߋ�2�/:Y^��W��}ͱ] &y��׫�K��7?_S@5�?,�yލH����{���q�˺
����y������cq�;�MۋUr��oJ|1UU��q�H+�7�n�	(>��=�$F=��ܻ4m�xM&2��6e�eN�(Ѯ\2�Q���+���@�Y�F�u�l�c��
��C�Pq���~gޚ�+گ�ՖP�*�K�$#ueP7ϵE��t��#z�N�r�pRn��j��-ׯ�|�i�N��iI�q�DC���,��(��j
Wu��gmk��OJ��t�K_��
|�o��17ܺ��O�?U��ԕ�ac�c����JW[��hʆ�ى-���{���gv;3��ɋ+��d�Ĩ���t)=��y#��/�����d��4�NyZ��w��������l�~�W�V�*6���c����xy��:�.��MG��c�"��������|�DC��� �nĽl�(8��K��H��i��
q���D��B������eLk�ZrNe47���S���V<�3iu��p�[�v؜�P�i�\y/)�9�Tf�-����1���[t�ɷ���鳾��<-B�C��cJ����H����J}�	a"b3Wc=pcn�����N�5��y�Ϸ�^<��]�U)\�b��� ��I��7���l4$�L��eZ|���lF+鲼x���ӓ�Y�E�ͤ�0'��qU�/c��ZkL�3]iI@Eh�"Һ��@H��kG���G��e��*U�w�u|�D����Mn\�Q��u����CvX����F��[�]�Z����7eu��|���{j�G��{p�0K���ϒ��Y�"�%%�7�Z�*䋹I�L��m�޺��$6��e!���9�=�>B�[R�$O2��������_
w���_!@G����8�NK��6덲īQ���V��3ͭ�Y�Xk����m����0gX"VDx-[S,á���V�=~��/�%�4�~����"�0����2��y��V�pe�hD����gS"ͺ��x���j߅7�{�> K���W���Ÿ��|&i��Zk����X�kh��r�
����BX[Sg��1�����6)t�t�U�ǧ���� a^R���Z,�n�����g�1�c_3 �J�8\�J�͞�o�S��YQM�1ֺ�z,q�ih5���D4�O�K��l���^�I��ۍ�ܳ�lpe�~u}^��)�K�s����)m���~�jk[�������"���ꦾ;	T��E��>��ؑ��wfۓ�YL�:��egh�^5�)^�R��F����)����*�M׫kP�`�ѫ�)�S��=�{%})y�T�l��#� &����g
���żS��޷��໗�~YJq��d`	���>��L*�2�o&��������R����Шȸ`e��o:��29�Ks��� ѥ�jv7�|ټѯ	op�b�]XiԆy�\7����&m�9�$x�}�rz�q�f~�����b�`;�x��),ukŵ"��F���h�ёP�!c��n����P*K!����fl���;ۚ�^)L)�n o��M�ι����4S����H����֍F0�t��w_�!ϋ̡2�y��-�:����N�d�#iY�9�^1$6ڸdb��M�W��՚��l���3Ou���}�|����Q�\�g��L��E��Jt��hc$r�ܮx�&�;�(s��0�����XW��\�a	���=�#TGh��jP�=����k�ҥ�oelrx��Ht�Hc�y���.����Wz�6�Y�mLV��8
ٜ�,($��f8S��"j��7������fzĝR�jw��Ԟ�-�Ԣ�j]���p�iY\+� �R�U�$��n����4�����Y"�l[ht��� W�۰GVݲzSRk������
a��Om�!R��?��Ӝ=?'�cK��J6�e�]�Z1�QRY]���H�������67�f{M^Vc�[���!������(�4��)Hc�
�Kk�ϩJ-(A����>iE�5F�\/��˒������g*_�^�Ȱ��EN%�,�����;� 2�w�S`��}y;s�-�6�7�΄N�����󳿑l�Gj1��r�ʒ��ut]�I�<�l��Պ$Z�퍡�bc��EHx���M�e��v�ï]t�����y+��:v��u�n�/g�pB������E�{a�g,i�=�7�Xk�s��I��A��u��ى��,��s���^%_R���spZ$4��X�� �d�X��Ms����ׅ��bT��k(���l�]{�l\7������$<�RW'�M!�%��[ěƀ�VB>C۸��>�R[<����4��\J��4"�"A�^8���X�^�)o_���`q��>�K��m��]`�|� ]nj��zl�zA�0�hf"e;y�� ��r�1�����ID��i]�u�U�5����s��Kl�V/4G�/�vM�����y�CC�SQu�+]�<F.x�@�o_���A٘��%�1�� L�w6�5D�z:wݒ�s���"e��e����NA^w�c=M[���2v���Tq��s����s
��]�f*��5�4{6�3�l�������x����"�d3��^Ќ[뗈�_ULR[��s&zL%�0��{ܠ�������Jt��;��OW��<�qɹ�^2��&������,��r����M��Ұ�{S_[Wzj�3������z{(^�Hw Q���b�X6/�����kkmn��8�K��X�Vf�r�b�� �M�7]��j���a����0������o��{����9ц�,{�.�@Ԗu�-6AC��
�U��qI�ƆAHt�.�<G�0[Z��+��5n�����{;s��	�!J�RP�xG�X����"�}���F�Y^Ύ�;Qْ
���rWEZ�iU����oY��'u��!B��N��Kkr:(�\��K҃i�B�W!�r^���pO�*�HS���bo�a��ѧ�H4/����+(՝sܫ�.J��yM_ob�.Qcx@c X뭻l������t5�m�'ä9y�ş�,�ٔ	P�*�S!�M8�����cL_�����<�<˖�t��M��r�IY�Ɖd>��M�kd^�B<�������**ݪ}ICA�U�.۟��Y��j��B(I��H@of�U���3{�m�̅��Ѽ����=3�*��r�t�òE�2/Ky�pGˀ� cRx��p<�'�P�c�H6�pnK�����oj�]��sf�s6����o[J�Lu�8�K�I^�+?|=���B֢�S���8�.0�"��kڛ*>�6�x�z�[]\a��µ�0)c�q��=��ܦ�fQ�b1H��8���!��K��$Y�򨞓<�h��s;kz*X��fhua���|����a����z hݍ:Q)�ch�x���"���'�'e-��1���1Y��*{R��#S�6�ە���\jL�ݥl�|����U�_�Zu��dMԲ�
�(�M����a�l=�C���%��z���{�LI�SG�=2SYR(Hۖai���._]�9ؕ��/��'@|�t-JQyZ�i�����H�9%̒P�����b��BƜLD�.��Z�Ǭp&�~xbWsrl�.��#z�}���q��mtť��"�+��1����E����m�\K�䐂��v�&�j�vyHbp��o�Cʑ	$m��"�j�(��P����.�6nC(=?K��+�*�dˠb�\`[/ ��5����aРuʡ/p+j(ni�ۓq�$P[�,�k�}	ۢ����$σ�m��v����x.����l�]��`����\xs���ʐ���� ��ǹ43e���%�&nm�����@H�[�F��>�j,l����%�Y���=ۙaG��s��lɧH�IN�vE�Xc����w����Λ���"��䝊F�~�0?�.V��_���w�nh���Ҋ"uڊa�Y
&����s���ΡdC�.B�� b�R��DϧS[l3,�v�����}����y�ʥ��ue٩]9C;�d<r����TZ�i��M��r0*�3n<�y��y���f�b����\X�x/l�q��ST��,R:�[�7@�n��;�R�z-�Y5-6H����!B�F���q��2��J,K��F!��p]��u!��"<�t��,�'?w�j�����	��ZE �)���E�=Y������MTN�	p�M!��\W��LzGQ�z�k+ `�"=��t�4���ihh��fw,!Q���b���)r�{Dz x*�[�hhy1����Ev�꞉'�\�s�k�ze��`R�G���{F��{Yd�=&�U�#V1� ���mR$�,�n�H���c�*"U�G"ѪL[KD�!���i�̨�\Qָ��ue�J{���T�n����%��n�xX�m���m��j{��P��0#?/�ҍ�}`!"p����K5W8c.H�R�g
��v�s���=���I�-=��O�B�RM~R_t��ќ+�u,��ļ\��Ukq4��ثMtu�:���H)"40
���I����L�3�A����!�C�yD�~���;G2K�?��ۏ��F�*��r9["�rvis|��g�-;3�� I475�'�����LK6�г]s,76i�Z{6���/�U!�  ��t�es�?u/

㾟��X� 4_�3;t"R�06J��b��@�mٔO+� �75�s����)T�!�s�1�x��5Kl��RH��f��R�p�І�5�ܓ��� H�����r4g�	f��8�X'"=�썮ȹ/C^	�^U�5�I&e͖�ߴ��ٺ�[2�U+����Q��=�v+t�V_�9Jњ��s@��TA��n@s{_2��=1kw>Q������n�M��^B�7\C���;C�qi")tL��{���+n���J�����θ�}���e�_W�&w��V�;��LYs�Lp�2Ae�9�ݍ�WI ȯ����]c��'�P�OɆ�\B6ۢ��F�����@�C"Cs�BZ�t�S�1�-�]�'���uDS��8FC�Uxm2�d꿇@�t�x�i��1�����74�i|:�:.Mͷ�^��o˘��|n���p�\&w�^�]5���'��s����L�#��v�=A�h�j����њ�5��K��(���3�L1n0��+c�s�P��Aw�_ho)���sE������V>�,���vI�r����K�:�SO����5���o%l��*�(U)�.���0�+NSV�^U���y>[SC�1J��~W!�s�B�F6�X|�����5š�}\��GB���:�� ����Ն����� �����D�}.	J���B���k�+��ɓ��rщ�%�&�m*̃9b��w���~�,d9��M�c|���G�z��x���存[�a�J���$w!͐C�2f�<�!��R�mn�I[c@o�&�M=��j�MM���!�#y����P�JU\��̙��3_.��%�-jޒk�(�0����Los䘎Cd�w��V�2�)��:���e���3Tp�5��=����etw�o �e�(�����������N[�]_�4P��*�\��	��	���HԳĢ������H)�✂j�V^:<;-����v��Xh�Ui�����}��l�3k"�mK��?��T�)�e�UA���c#t�h�T�/*y6͞S�� ���Ꝝ/�0MFky���759�ͅhLɅ�c���:n�xKE���{�AT�XmT�h������ln%����{����$eLJ��X&�ڹ��ؼ����]��^Y�.���إ���J�6�)r�5rG�z���~]�9��m=B��{�k'�z�s���Aw�f���,)Rq��{Y��R�dF���dR�A�v!xR覕��tĵw�����^Jh�_h��ο����p�fA^[ܺP���W���96��
�z����ѝ�𪫵�\�^��,W,T3B�(�N��%�P�Ew��{\x��,�W�IlK �8��|���:])�XǷ\��=n�j.����x��eN�Q G�w��@z=����=d�z��'󱇂�z4���T�R<)�.)��=�1�Ƕ��O�cp�c����;"u��a]۞���o�D���8T�$�8�kH�5�i��k�`�c��Y���%qj�FQ��}�����~���yW���άCTy���Y�L�#��z���	���m�"ou�$G�P����<l���y�'_(RCI���I����dx	�*�W�^/�bE<WV*�qY���S�{�JCq���=����)Ф�k�Du������Nܧ�H��f��^��8.�3�?f#�ڹ�|��|�	0��̩������1��߫F�n�g��F��Q9��D}�Is��fL�c��=�z�%ⷘ���
�!JR]�@����ҫ�F�qm����1b��D71]qO�V��l�j����Wg���d���#K�4�c�m�5&Z+���>,t!i�¬qBmK�x|��1����Y��%�ϫ�4��ɝ�z�5S�m����bgr^�)��N�*���^a]���佗�<�s�����D�%<�<�<�r>>��=Q�!��Uq��xA��y���}��W�z0֌<�3~5FJ��owww����~B;C���pյ�k�H�V�Hu�k�B/%�E]��D�r��K(�����Ӫ�P�6; ��u�4�G�Zn� �B7������z��ƌ_ή �Hp]+@C��3��qQ+�+�(C#�����(��l�Ce�{U6C&�,�]hZ�=9��9ϜS���l��'^�{��D�`��v%���W���}� SҐ�M_�ێX��C'4t�I�1�5x�K��t��e8K��23���*����}�?��U�q-�.+�(E>���tU1؃����&��׬��q]��=��5u��&�>[����ZY�o&]��3�g�qoX�݌a\Na��.T��F�绹��kd�y�Ǔ)Q\w�}��]T�܀�U�{���51���q/�rQhs�Ǩ����TcU��Eϔ����z���o߆"��/�Hщ������H�G(ͻ�T�0�T��נ�&MV���-��B�븄�!Re�*�
��$��ה͝U�}�m�Ly &y�T�(f�l&%;����j���x��*O���̮�[͂.>aBE�kیA��8��=I���n��a�!j���׬�(U��4L�Ŧ;Me�8Ű���܎����O1�.w�\��N��Ѕ)����[,Ȍ#v3^�w��(/�aɰ�-a2���>P�ސ��Hz�m�T�ol^�lw.JJ���)U_����o�Q���t�p�%�Ft7$��F�jO�c��5>�쨡�}���o�r9� �(ZKMdF��*lE���/���W����"��^1_x���%;���T6%Sj�@����P)A��H.OPn�&�lc�� ϧMx����� �S����y�1Q�1����eW�:��4�W1�+!ү��zU��HG������*�|�T��2��|�po����Ѭ��l�]��N
�:ȭ���n�H$HJ�)�pY�G©ʇD;YŲx����`� 9��F�;�Y� !T��0a�վ���/����s���Q	W�ǹJ���`|�1�6��
�O	�B9��kݳZ��ω+ڝcۘ5�"�;;:�v=�x��ۛt�"���K7�簄�-o���XkQI�n��ڦ���B |����K�&�nE������?P��B��0$�O�͓��������=@í}
�|~�qu��gO��I@����C������O.����)� Kz:�R�Z1"�\5��nW��V��דL�qo��^�tVR)� Ej4,$#��=�k	c�5��óL�?]~�+Ƈ�^��Fp(6Q�4F���Ӣ��``�n����Ye�dp��㊌��G��T����(N'�B���kD���2:�����Si5��Mr�l��7%h�GE�%�v�(krJG�.n)�(�j�04b���qL���x��PY:���j��'޷��m.D�V�E�`^��r�k��f\���$Q���y(�>���:�#���M����%��j�+������Lj$J����竲#@tg�)D���M���S|6��R]����@a[
�CYt�!��~?G�M
R���aۖP�����Ɛ�]Q4cx�r���Ux_��b���	��S!���?������(����qdX�Lxx������C�^�*�+��/h?�}�|�w|����c%��/��@a�}[�odX�2i�}�+�j-�P�����q(�B B�|�A}
G�pWZe�V�L���c� %���ֽf<+���3�5��s���@�J^�<ͱM����?�����+��9�]ʺ{�޺+`1��Uf|7i�т@u#��d�>����p��!�`8��Z�K�`S��9��1Ez���u����Y֧u@�J�������u�OP��V���sK!�>o�6�@����v8h1��~p~�Nm[��i��{G�TV$�Y��T��s��M	_D��6�o�D��<)�F�;�:�9�R�����Z�����:�X�xAyZՐ��&a�qѲ'O�&G<��MO����;��W=vd����,���0k���`��h� <�C��+D_��}�k��3(Fk��"g؋e�T�DA�H|4?��W�,E�p��a���fl�������O�!\o<;�H
�
�������d�C�2\w��$�}Ng_�K̞�KYO/=��v��-ۍ�%�o-�|�3�٠κ��&�U ]�H���T�^oV.�����w�T�Z{'���э��u�`H������(�!�)��JK��!�#
��U.XZ�}�D���lbpbL��ͧ��
��YdW/h3,�M�����m��,�fc�m����f�Bg�f�֑�hV<Ks��8�g "�*����2�ٝ�@!���}_?�/�g�ޞ=���Z��N��\_�K�i�3K��su��nf���I���*�(���>~����8�K'
�.��~K�yrJ(H�E\��ӎ��ŸK7R�GgF�O1�H��M��n�uE,�%���C.����>/`x�(ҡd��kk�5B�"�k,�a�ǻ0�;SJ�Xxl�������Xo�O�S?G�ʞ���p���9���aP��H��7�<��-F���
���9v�7�QB%��֩9�Ԃ�4#��IB��I{ck�ϐƧ��l�c��d���2����o�1Y2����<"Ż�ץ��Ɗ�b&�Vy� 7�;��mK��P��֤-��Q��ʳ#����l7S���~$�"8�EKcq�7o͊���/�Ç�� �! L���ú���u �ie����-f�>.N8.� �	eZ���72��8�ֳ5O��CQɝ�畕U�a*YF\삟g��,m�B�7���C�mm��P�_�8��*N�%>�]Y�u�M�>w���ڻ�6��8���Ap�3�������H<��Gs��Ї�7eb@�C���z2�~�����qëJ���m5ȎE�2�Lp�r�^z��/Śm����ؒ�'W�N�ꕃ8�������z>����yK7�d��̦˃!
$�0d��1���OxU5���dU.���`�����������N��a�k������c�/�fgc���b�8� %@��}��ݭ��$O�a��B��/	�L���0�x�W E���>⭶V�g��A�`�ݛ�!����G�� �9����h�����
��� e$�2]bB7�c��!d�E��\�K(RQ+4xh@������&��Ӌ-@e��^E�������;���������O?��aU�o�e���⋙�/W��>z&�q2�"����׊
�:��4�B��g+��ȑ*��PR������z|�R��(�`A�Į��U�U���x�/�VxV�Ʃ�%�"�٭�[����	��(Ct{�r	�3�(�#�Z�0`.1�_}�U(Q"���z���.����)�sO�����ɲ�9f��yȤژ�NX���=�JXA1z�nq��+�j�?;��U���ܖbZ1�Ȓ�*�]��ݻw�8ܵ�����==�s0��oq�+�����u��B�����۷�L�`�t@�1�R��)y�2���䝡�J��.(�O�?۽���9`}f��0oQa8��*�;�0�b���gH�����c��axA�W�Ŵ�aݽ����->��a� �Hq�Cҝ �"���m��5�>����_���҉q��1?��<$�ب�N[
��R�z��@ִ)��+Þ�0T�	<&�eL7�����Í�����}�bj��"iqCh!X�����}�ȸ��?��~���U����:�m��Y�T���?��zC�#�	����}�����r��ŬiA�������f��ȖYu�٠�!�N��`��ΐ����u��ݝŸX�ؑ�\I� p�0,���(�����X�oL�qNSP��N1��ި�()��1@�7���7��u������Psko޾1񹽿I��hڊU��@�٨M%���� �wͶ�н)>j-�J��>����גަ��uL�"F\�iUr�;��#���R��`,a�/��~�~0y�}��dTن��V%�*b&�pN(�Z�Fo�{��a]g��=RZ�9q����?������w�f�>����O��fw����\� b��,�
�3�B�\���<=��)f�;���B��sךԪ]d�eH�H������C"��B6�|tgi\�Ǉ��K�p�<����� E�gȀ��q˴�}�"w��T��_*�Ɠ#>=�-��%�+�آ��1& (D��~����cRޯH ��& �t,��@�*`���5�B�z3�+
������kQ_Y%�d�\z��ص.�㰉äU=D#c�?�*�A���4���.��!㞮�`��-�.XkYE��ňq2tW�M*�P�&fWVo^����U�~5��sB��\�)�Y�	�\-CӗP(X���/#��
(��=V�!�`c"�ǖjO>_��~Θ鲄��Y�Z==>��y
�����BNl�q�}�,t�h;�9!o?���B�����*@q@[�y�e&;�qQ(c���c��V@����_���8�5���e���ƓR���JJp�Q��Z��}(XR劜	>�d}ǳ?����w �{Ý/b�Q�F�� ��1'��ޮ����2T2�8�J���u2�S�Y���$Ӣ�;��c_"��&ܕ��_���+����"�[)R�0�䉩�\ɬ���b!�_~��·�;����_�$�3h��h�,Ѓ��:���^�����tr������O�����D�Τ|Q�N��Hҟ��)K�!��{��e���\���L�nDD��@]�p>XnX��*#:y�c((.�Y��`���U�]q+{�C#��+:��v?�����f��/��b����=��Y2k��^@xP���Y��"D��)b�ճxa���S�	M��Uqb3	V�A6��ע�=vW�B�{��������x�XJLW�6@COD�0^S0f{6�H�ҭ���dn��H�����^^:����$�Z��E^d��ԕ4$*{܋2�_���3��p �Sb��IԻ"�=e�����/�����㺗�\�lМ�%�)�Q9S�0����'e��(;U!,� �CZ7f ��*(}�-&+�x�i:o�Z2V��-M+Y&u���4,��Ev��FN�'-�V5��H�>;�>���oG%�P�ל�>�B9�_���0��Z\jU�O+�� �e���Dd�po�(L�ϨD:y���*P��x/��a�(����Ǘ��?!���!N"�[��f@_��]i���bx��ɔ���NP>.�'�.�D���l͓v����VK��X�h9BpS1F�ɡA0b�pOE��k9"4�s?8�i�1�\���}�[��5~⚘�_?��I�3㭗S�$j��ӟ�������2Er��UiT&�x�������:�ό/����qFk�$�EF�rV|�P�}^���7_[�U+J�a,q~��-~?M.sR��-VO�x��w����b������c�]�ڳA��2���ra��`��E~�uv}�A͈�;���[����x���ft��޽�sclqN��Q��'w�l���ΏO����0��bxG2>�(n�0ח_2��@%��ט7��Ֆ�%	*���R��֝3L������4�8���P��e���[-DԲ��t��
��㺴S��f�'��&GJUu����K�,.�ɂ����O�?�Ы�$�2�l�ᦉ/)�عP��s�H�͒3�-���N��U��i�ЛE$IX|��T>,i�!�0/,��.�=\��YH�>;�D4���r�ĉ$��K�O�z�}(1���d¤$����|q�'^#���{�gWlcS)#P'��-�@�X��o�ǧ���̅"Z��[^	k�v_Gk��p�$mjQS����������q�~?�_�r>�5���J�$s.���q��:���nYcs�QJg�b�����mF�1g��4R�GM�Ϙ��Fơ`�[��a��bA�2�<Df�	pL�L�&�wβ����=V�?D�&�R�Ԣ�nF�����P�%E�g���Z�����K��8�;c�-in�ښ�t�
�\!nz���� ���(�B�Cܧ�қjʍn�W?K!����o���o�ұ�p�����y6�X�z�ÇP8�Bt=n�}+;E�熙^�Z���9�l�19۹p�Ϫ��0����7���_�/�6�z涮��	4ג�X�rQ��W0��U�}�d�6�e��㧾��n��@���/���EĹT�1zW"�_�ɛ��� ����E�R�_�J�/&�ޘ�5OǷ��zk"�����)N%���U�S)|t'�����a\��B�??�4?N����a}�>�}"�� �D����,s}�.5b�G�ĵ,��x�]��-t4�w���++�U�CC@�?�����&Vٱ"3�'�!|VqE+-������(����!}�?x!���d��X>�<���@�h�U>���y��J$}����L���ɾ�q?�ThG�n�M�2ݬ�QZ6}&�E^����u�$އƩ�I7�d���N�¸4/!d��h����&b,l}������E�].5~V���&�6&�+�T֚��v+����s[|n�W�b��TRQ��57�¿q��R`�k��!�'���<0㈸��$�){��!�$f/��� ����AA�-���ظ�Ȟkﮈ)R�p/�qYk��=,c�5�G���%�0w������?��?V�D+[��,r��']F`[����;�t���&� a	e!�Y��q�[|4��Dɖ=8�_Q50R�~���=���Od5|��l_�n>�A�ӳ+u�ÆDuw��`0VV��9�8[�u�����z����c�{"�m{�Nɘl�Ȯe��1����@ō���F'2��Po�CR$)UY'�ϡP�%㼃�JHE�V�^�)J�UNL�|狖�U�^��!I�ǋqM���\���1"�#�?���a��g����M[޸�PHt�W�@�̙�Fw���Ժ����
�����(��¨W���J�J���l�R�{r	庶W����БYt���JU���z�v������(�m��Z��BTQ�X?OCS̧�#�f�{/%�b=�<`�pb���&��!+q<d ^�-e�H��4^�/��dUѝ�%�P1�������4
����;xv����qa(��S���p���Ѹ� ����/vN�O�A�B�H~�b���Ѕ���;RCF�w�F������PƔ��)�8�=�K4O.� ��RoW��X(�����n���7\w�Kܻ�ʍ�o�>b�1�k�BZ���]�4�;�A� n6?<��~��_}n���sɤ3��?�����;G�^=�F��crO� ˅n���GK��E}0�D/������|ë�X�1��s��x|^߿u����.�1K(D<��t�iwWy�Rj"�l�W����]����gCų�8��í#��� ����x�i�<_���*�*���_�2�����ӯT��|�Z����{[����I�W����z:U)r߸��6��o�=�y@�5BrB�f��� ֊�h�~d��Wq�8�z������K�����^��'i��� �L7ۚo�����A��h�H�sܜ2�p��#ӣH���/�;���5����u�.�E,<罻�8�n.H�ѳ����ӝ�K`(,���!�q�/�Z@%��|������X5�OO>��%�K�4ј�9�#֌�f�b6Z���p�T�\t��;�v��@�
��.��<�J����I���Qߠ#���b`���Z,�m�'Ɗ�E
c(�L�?�6�￰��0Ηܱ����5�ŀ�;�;��<�G�ޟ�Cx5�^b� s�q)�:}7R<�(F�ųܘK�9�����-d�l,[��0:�R��Ce�����O&�޷&˻�bޛ�	o
��=�հ%�3׷��)���UER��5�u�M���=��k�i�2Z�P����µ�aD1366Jo�k�g���P�t��\܇���R5k_u[(ّF#��Ͷ�^�������׌U[��+�7���XE�Y�Le(�8[����[۰Յ{{��
�	��n�ܯ��u��h�CZ~|F.&GM(�U��;/����b�X<AYq�kX�����?9O�C�)N��d��a,���3����,���ǟ��M�-�r����o8f�`q>a<�����L|p��vz(R�8�Tԗ)b����|�8����}祧�JX�tq��������w.�%�<>�4U�]� =�1�
k@f�[x�x_.w�0bE��yX��\��q�#|D~{($ݷ5M�g-�h��k��`���.�'w�ob�����#	�d1�=r�d��b��TǑ(h �Ǩg!�M$��2Wfh�N.�S�|��Iw6�"��qB<�Ь.e�ay3j�S]W��ɥE�X��m5_p�P�d@�t��#�W����.0���9n�W��BJdg�^��ւn՛�fX��ǿ�����3\����78�����]7^��h�=g�䩹��0�${�`KT�s퉨��l�6fBp��q�~�7���-�ƞ�B��g6�I4>�7������ x��g>쐈t5��.��z�J�� N���Q����$Q������ZRN�!z@��om�￶���ovO�|�M��߶/��2j���^X����F�R'%� <�0����-h��f����H´�n�8��{���)Qܳ�9]*U���CW��O?�+��=�iݭ�:,�/V"()k�] �A<�{w�(�ÝO*�B��b���r����Q����φ�n{�c�M&9.2l/<�[���yrw���S�N��u�q�莻S{�?9.�Oœ�G��'ƣ��\#ɉD����M�W������sd�3�Z�S�_��o��e�"����T�j��ܑ��F����8�4�zw��Fz�ɴq��':O�}�0�^֌y�(�)ۄT4�$ܹ��&Ej���J}�q}�R�����mA��� O'�K�AW�Gj�����|���"-٤���-S���+Z��Tk�a�ٶ n<l��N���#�-l�*�C��	 Z�F���P�Bj��)���8��7��3n��Eh�5lv�Q���M@��j��cq��Y	T�xR����.�:�Db����>3��v9��7`Q��,��r�������z0d&/沙�u��๕>���˷7�����Dm��deеg��ήO��4#/N�qҹ��aάф�8����l�c������'��2cG����2w0d�}#�|WE��?Ի�;*�Q�_�,2&��s�)�y�|�Pu��D�/xc��0�}G-N��&&� ;���"o�vc��G�X�'� �6�B"@@ٳ��nrS���W	Y�}�FB��B	�]�K�j�U���L O�������;���ͳ�6� q��*A�6��x啌Lm�r�<u<�RURsm����I�I+�擇�����H7�'����3��J`Z�%MN��1 ��{� "�n�*D$���I�V���������d�ѫ_p?IE��frHI�WuI��)w+ȘX
��3�����YՅ����n�:v@�����i
��w�sq�\4 P��L���u��ۼ���S�p�����1n�S�쁬��W%(�V�8N��aR�[裓�w{�b�'���t��T0�\Gۣʹ��-��j!���ͳ�֚�%��?������O?�x��\ͺ�xp]�U�=*qZ����%l1�[�>�ʠ�!���ҍ<d��<8'��x����U���a*Ҩ�h\����aI�dN.kU�2DH�⹕������-�g9�6�S���L�>��ZW��W��{�� ��17�ߋ���%/R�L�ђ�5���*o�yBV��Œ8�|=��γ����"��Wyj�ㅱ�a�=��S
��!C�,�?a���u�����5�4������g������&Nq���أ5����}Z�#Ăb36׊!��-w�dFRM�] }��C�$��M����U����4��v���^	�0h˒ƶ|��A�R�j�JU'Y��gO>d�]���4��N,�V�1#Q���Y�g|H��X��a�3���?������	b���|3w��ث�njj��K���4�ME�Ɔ��Ο�1�;e޽���cg�R�����K��뼖$Y�Ż��_��T#o(0>zl�}�]`����@lϬd����ў�|~::0IԠ��N�y��%9	�����z�=o,��t{��^����2�09��w��2]X~VJ����;{숌��'�5妑��T���:5�b{V_m7�����(�g�;*4UF�����M����8�}�`ct�a!R)]�c��a�����`�P�ry{���QT�E4��'B�0��Rk��cc-������?Y�<��zz��T�+�z(dﵲ%��=��4���������ɃЁH/9a�X����(9�w�&,p�q��0| pVYuv!JƮ�ޭ:(W�7�������ˋň{#!y���5G�S<+���gM��i�*	���ؓu�Iޞ,���C���{���Ǫ����5��gvɹ��l�i+l�H�w�kp�����j���m\��%{����)�⻉^"֊��D<m�(�%����ԃU-���&җ��ϐ�{�x���H�v�
�#)D\|0~�7���?�bW9*��_}eJ]����#x� ��$�->��-�&����(HGn ����m,������|cq�/�� i_Cd���k��3�qk�Y�Cdtq����#�"Z�!�er�L��yt���ݳo�A~um�&D������-5���gӴXǸg�2vIER�d�|2�Q#n�>�"U�}��?��"��8�O��",�)��m�Ⰻ����?c��+��"��������1;�yM��"��q`�KR[�'<RG��[AsYz��j~7�(��J���ܵaZ& v�s衆��Y��W9��ذ���a�����vAL�߾��<Z�f���m8�Ư��s�.�/^��^h�;?jk�1�x
����'�1p���;�֒]�G��8��1�jP58��j�������
���H��t��i��m|Zw��q�j�k�](s2�[� �J(������5�}R�D�!GQ��T���N[hfU�@�
����s�S���DCOA�"+� ȇ���s�}��,�����Vu���]��Ũ����K�I&d���}(`�-n��l�U�L���~�bƌٗT-�Ы���ØՂ
��QUD7��>E������<�\�"c�bO�2���F��Ѝ{b�O<�m�Ε������s\_� �E
IK�h������R�ݷ�{�~lbOZ��=���{���s�RhT%���.���K�|��E�������X��
�Nd�2���-�z|�"�B7�?o_�Ba�)�j�W(N�����Nŧ�E�+R�]�����_عH������+L�8 .�sxVeNVH� �9�hIIT@�5)s��Ʌ"���{�P�+�vp5���jy�ث>=>:!�%�f�NL�(�����ʀ4�[�����؆xOTH^ Q-��'G����w�/Z��H\$WS�����He��VE
��T�yTB}r%�geOT��=���"�g����zlA�m5���bq��g�?������HَRк���5�d���66�BIȷ���Ǫ���L�X��i*L��o���O9'R���]po���̿5����s&r������T��<\��L�O쎛��fU69�f�c��*�OM{!�+Jz�'��h�^��[M�.S(:��Crn��5h|Kq���t{씱��#�T�W�JC/�����Cª��	�-p&��~~t�p�&�'�"ǝ*:Xc�N��j�V/�G
�����s�b>XsƇX�C�K(;�C��h�����sW����t�Ϧ���	h"�^��ݞ���!/ >����`qP�����wW�(q�l~¹ =��	���߿��ד�]�e}�~�w�}�!�7�cB��	��Ǭ)���Q�σNN�����wZ�e��^K(�RA ��!]k=�������������g����P�k�7ǵU1d{�Y�"�C��A5�wN�BÂe/�m(F�(�ڄ� t��� &�D7��ʤ��˄�y�Pj� ]
�V6�`Ƶ����A��?����?�Lַ
6C��m�E�S(,�{8I��M(�~\��o�Ka�JV���"�``��7� �H�׃��5��ό�����4pڠS'�9��  �vN�ސl�n���]���{���hz���)
)6G���D�2յ�A�W��Fl�#�='��Y�F�\���KK�jY��iN�ڻ�����Ҵq	J�-��@{.��=�Xoqͳ[E}E�Z�E�]i�g�E`=�����B(�R`P+ƭ���'������V�)�e�C�j*��1�5�HX¹��˟-�޽p��._������S gܯzEVt"!�g �#���Z��q`I��ʬ;�cqw.d�Q/c��@Y��⮐��	��{��45ߖ[�0���U�M�}������+��"����&[�E�Ě�\)*{,φ[��T�Z =׏^�k��ֈ<���C2{m}��u֖�ֿ�6�U�]$�{$�$i�]d=�9OsY۪p�^'�@a�)���P w;e�S'I^�%��#7?�,��h2.h|..��ȴuL��^e�C�����V��<�ZH�q���潗�k�F��H��Ԥ�<�y��������G��('���}{��	�{����n �	�:��uڅ��{�/�ϵ��>糺m�2BC\����	�����X�FT%�H�ݵ���'*����G��1y������b ���^U%�J�.R[T"R�ڜ���n/�k���j�T��������w^4�[�MZ�sR|�����6�~5R���ف��ڳ�f�Zm��?�2�uѪ��dfR��9���Zat�\�}�_�80Q>w�?���v��L˵��T^��r\�==*g��'L�AZ��W14$��J�1��֤��9��-����O0.��!7�H!㪤���8"kE+N��y�jZ��,.��*��H +�=��=���`�6���i�LŊ&�ٶ����y��r�Ϟ2*�J�U�ܝ+Mzd�J����X��ݓ����+ � m�'��J��k%�Z�t�T�?	������'z��'��r1�$��J�$�'��|!^&�X��=�ҶRM_�t����)��g���r�-���}����@����|���
:D��	�QPO|y�n����Hd�JAYB(����*�Z
|K��9�dA���BS������51��{�c1���,��P����-��`
Jt'�%*/M����@d����N���}��ح��bc�ڹ�����qKCesnu��R'�o����سqLl?��S��BruC��a�8V�әat�TSe��8�_z	�nv]G�\�+dB�f��V=���0оS�N�]�Ձ��K���0�J����N�U<��#2�7^֊Ј�ܠ�_����xm7_�� M�4b����{��ِ��!��㆕)������NM޲GK\� '7^�$�2�]��?�Ǐ,�Ѧ�*)_Zҿ*\^�|�@_K4m~�(�Х��*m���	�T����bp{Q�Bc�Ȋ���g{���pa���C}�7N��y� �H>��0�
�b����q�����2ˌ����[�ekNoai�ު���@�����v�ɰ��S�n��w�r�1���
��i�� �Jj��e˺�{�l4����wn�+� �]�n�l�.�ώ=��nn��T��uj��]'�]^����=�.�� $����+�	]ԕ�K�ݾ-W.��}��L����4�
��}{���'n��h��s(Ѥ���n��#���}|fS�;�j�'C[�R(���9�-$�b��H���FƵz�~���j[����6���{K��2gm��x/4��%b��LGW��)����8i����)�S}ie�d���j��Y���1~�<��S��G�q*�)�)Dz:=�:�U���6�1�ρ~�ǣE�m�\�XS`��dU[�HCq��_D�5,���Yd�8!�ɗԾ�j�M��b�u�ܓ/(5�9̒C�A����n�*��"p��oCv����l���j�E� W3���6B�3�%���O�l�yu�0Hn�Y��(��N�i�a�R-����%�h_���" �s��.<`$52t���F-��� .�{��)'KRA��V#O�	�XUKM�HW�=�#v%E�k����{d��5 �9D�
D:����y�f�էS�'� ���7��?����K
�:&�L:�#�[&~��'����>DR���x����ܳ���D��|��/�\y*c)�F4,���$��tk�X߈9��8���mv&g�+ �h[O��<�W��S�C*�ը��]6��{���۷I�R�P��0�PҊ����D�*��M)y�:����pQ]Ĭ������"���i�F1[=����jK#{&o���>�i���{J������ ����4㣆|<�i�<)��߹������jYm��n/*%����QZ��{�+�s�
�����3�e|��d�IǸs�򥡺G��l ��g�EH�j�P�v�e����5~U�b�¥=F��g*��+Ɠ3��=G/�gS����w�{����~�IƗ�D�w�ΓY��I{8Y����
NYnm-����u�d(�'oF��BJ.��o��Y�8ȅ���	���:�iC��pҞR�'wpXA�/B��L��W��ʘ�$�ԗ%WKha��$r�u#��IݤQͮa��R�������
�eb�� *�98��s�=`\l���q��W���Y��Do���'���D��:.��(([_���QZ[A��{�
���Iq́ܩ\� 3�<�nb/��	@������ѥ,{���(g�*���Ԏq�{�-S����g��Sŀ.	z�h�-���<�3DD�s$�ΗdU��/e裄���z�t�_|�����ض��"Rf�TO�O����<�{v�����9��V&MJR������b;/sRu#��m |��@1�P����)��&�{����@�r5ɰph���ѧ+ў[1Hq�b�2��
����γ]�W�L��ۃ]R��� �������G�.F8� �ݶaq�|��l�|�#R�Z0\��׃#��Qaa�U+X��ַ�\� P�bU��6�I��ӈ���V����UH�11%�|Yj��?��A��R��b^���/M��]_q�Gߙ�6����h���q˗��A����z����������پ�
9\��3�a �"VW "�k>ll���}���#KZ!H� &l��>&�*�J�� �����a�����>�.hj�Y�:*K?�T�R���4vv��U�_X��F\�!��/�#�X�l�$Y5��ۺ4��Ge!3���f}��U'��������
��K6��ի������Uw��>�8N�M{d\E�]
�h�JxH�rO�n5��:�	�\?�͔���ל�
S �˩�ߙb) ���g�7�>d狄�yur��\�l[6[�$��BoR¤*x�s���j�x� �z3ܘ�1��^t��i�P���^s�nqځ;��(�����-[d�Η���|�>�*ە��-w�\5Q�<q7��9����	�y͋E(BP��w����	�w�|�R��������Yq0�MZ�y>���y���B�9�g5�8E�����qÝ��]p�Iyr�~
�h
e*9���xY;>6�:K�q��5h>x¤mb�эi69���n8i��IQU�	E�Eݎr�81�Ѯ���� �v�G��.�వ�xd�r�����)��<��%�!w��=�d���M��.��BN=�szfY�IN���ʧ\/���:��]��?6d�*p%@���D!R,�h��S�pO^�� ��]�"���g�x��P���8�Bʾ5�x]|�7�F�H�"�J�[���ܴ�Z�ظ���@X�5��-�RI�6�{�4�%�;\���7��Ƚ~�W당"�7��$� ��Zu1��]�U�C=h�o�o͞���TՊ��}����g����0+L�mev�i�<�W�xR�B����W��dwܒb=-��ޥ��w��u�0\����z|T��y��[Pdܛ��PZIR���D�\�0��ה�����#]�bE&�ٷ|&�<�@� M�L��S��ڸi*'e���Z�A�ùŕ���*�N]�Ll�f�V ��)1�Z���竚M�j��ŸY����'c��Ԏ9�u�K�UW(�%&��`;G��ϩP:?��wＤ����hZ4@b-n$$;��f����b��W��e9���O;�׌��o8���Go�|�&��D�T�J��^z�K��dm�����%m�=b����Y��A6��$xs�#��`�H�b	P��S�5�����!>�~�ۤ�''�ʲ��~.{o+&�d��8V��
\�����2�
�3ÙƤ�"7Q�Ce���(YP�߬J�޾��}X]Y	s�VntT��Nʕ7��^��ۣ�F�p+�]~2�/���������n��J���h���$q:R��?��3����D�"5>+*����(Q�yts��W�~~���~�k��G���㻦u��]r�+kB��Ç�gH�iPM��8uo���W�Mff��2f��f�0ؒ_�Tx�����}�si�YV�A������Θ,�l��ی;+���~�9�⦪2N������U��}-�1T�F[؟��8��̃ws��z�nĨ5�	���܂=���k�6n<���՗X�Qy�HO�ܽ�Q#�H��?����/ވ��)Zұ�F�TS?���_=~�־_!�q�mH�^L�77��~��%����95E���g��ҍI�WqX��L���ɮY��}�mr�e!]�}��=:���$w�[�~0tc� KoM-�_�h�Z�Zf�r"���ӟ�d�tn���u���EcB"��qS7z,j���÷�rq�S�*$?��C�n�>�0�g��C��/��x���c[�����s"CR��{��-ka�	JV16.b�Sj�}�h��@�b���u��Vp�R]KD�$��%���A�B��������%c��ۏ?N�̈os{��T�y����=��^�l���e��0nvHn(� [;�D7�d������%�J7�j��%K�� 0T�{@�0C��=C�����o��u�0c����9��7ߌ�/��j��'O4���)�+�v�9��E�����,����� !~p�g̞�,��Ay��l��[���%x��/��;ǵ��N�``���������o�7[�?$b� �B�o19���o�F��ʔJ�w�朊����t��>gB��q��p�� �Ɓ3���GGi��`i��S_��~>��]�={v���Rz�������8�X�� �`�:�/J�g��h�>&R�� Bc�VёVNn'�d�M٠�C��+�"� kQ��<zB#��aW�O���1ceJP�[��R��'�vu�fŨ'Kk�!� e���#$ג�烳�L� e!a�՗�*���%����@Y��+��˿�����{n���s�'t��|�|�-�|O���B۲h+	.T���6��n>y;�v�jȣ�]7���v���e��+T$z3���,��[�(qn0x4���õ����]Bi�H9�������
�Ϧ�w���θaRV!�������Y���c>�Jp�N*�V�G�A�Xz���z�#�!����q}Əv�`�b����"�1<���<iǈ,M�-=�Z|�[��k��?��>�L����Dh��wr"��♗�ƙ�"KHɝ�����Q�'��a_��R���`�G��k^�J���[�V1)���"��sdH���)�@,�\���b��?H�$5İ$Ѫ|��p�����pr4�T��\!����b��:J��P$8��K@��zA��>�q>� ���s�KxȽ����b|��ch{����d�D>�5�W_~e�Ol	ۖ���8�6�����{R�*J��F���a�^N���������c,���:�JV��I���=����*��R�K���bIhW�q�Ap:�{���T��yWiq�m=��֛[��]��/I���u����)^��]�����8�*�Xi%Y8�A��x��;o;�|��L�g��_�k�q���EIRS����nY(P)׀8�
�T}�~�d2x��ų����	kGr���1ҪP������mE�l�QWqQO�]���"��L�v�-�yX�K�؏i/���pqe:9R�L��1A��)`�"*Ū���Q���UҶ �)Rc����6s�=t��cr����������^}�)�Z.8{�Ԓg>��U��@�����.>����&g��0j�bX���;���1�=Q�:$1S:�1���}�?'������`���*-$6�^�.��?X#�'�!9c���kـˎ�����JV'a쭦�_�U�O|��Q��V�"��T�K	-*�l�A%�{��k8��������b藡�7��[��ۦ�)f����Z�����8B[P�7^j��v��v�KŮ�Q��L=y�喸WŢ1��E�3�@�)c��Å���8���+Cow��<��>;<������GשOG�pA>(��x�R>C9�32��]鷰���U��h�*�w��K��Z�9b�b������F������Wh����te(�W�����i��;1y+�i��+�����[�O�J�ҥT�BE�*�&q�98�`E��ܨG��+s/0M����@��T��~ٗ2K��E��O5����K��n�E�ͬ�[` fY3HO��'�?�X��!�2�2��9>�7�5W)��C[��Sr��ңR�:�{]��Ѳ�H�=#�j|�U�Ɲ��؍���ֲ�B����;:�1�O�R�9<���͹Yq4��`Ht��Ð�n.��<���jՙ�-ʋE�Y��,��P�Ns���k��c8G(5�?�Gۢ��P���ߣѼ��m��O������*��e��[�#O���]�)e��E>nr���q���# Ej
?Ш���^�6O��u�v+�a�\�U�"	՗�~g9�a�V79%K(�*�<dH�{^��w|���h��P���������:|���W1��Q����@�R�ኈ͙�Lڟ�Af��-A���q��)X�9�~��R�r��*p�L��p���C;�;m��U JV�^�%�Q���%������MĻ�Yz5f>���z�/� ~�(���P���u�4")s�u�|{(a�  T�8�����a�ϛUa��>�+	Ξ]����}��nV��#V���5���?��ܬ��̕���'�\-�d3폎Ȳ�E���NO(fp�����[�����
�P��bØ!��P@�8��K�\����JF�KW&8��њ0�^��]�Γ��<��Uf*A�k�v���)Yy���s6�|}��Ɓ�6������5�A>>�����Z�b�����B�{��tt�0�
�p>�;˖q����j2��Z�d	��~�������	���	F �x!ݰA�vC����H��c����N���6_���{-I��X4R�h10P��������9���.䈞��n���{d@y��+��-��"#\����CVބd�ucC�y,��"���
�~	�T;8l�ʭP�@���n���7�wU���s������;Rr��*�j���q��G��T��ʽcHJ뭺^Ê�ѣG��PĠ�*�����4F����J�q����!�� p��m�*�Q���<6;��xԠ>:qj�ٍ�62�7���smVR��)C�X�1,��n(��<ݾ��n!�LG��P�w��<���s=b���0��/����ĺ��+5���̆{�f�uB�vu&}�x��59W��:��YP���4�) K�+}��e���vE�g�e^�,���?�-�w���y�ggZ.f ~"���\A(6�-�p���m���k���I+b�(Mڧ&��T�4 �5ıu�1l..���dbmHպ-N����9�̴>���u���9M��Z���Vq{q���|�8v�L���ƀ��pQ��K���z�:��}��0œ1��ºN��"�k�Y�d�9�S�4���UE��`�3%�'�`�J���:j� �C�C<���O#�U1V
���MI��hʨ�HiZ���������_y^U0�U�6��=��=�h�`�oN���p0��H��} ��hs��>hkEu*�0Ћ��ƵPt�4�9*���MJҖ�U����
t^ܢB��E C�ej�=S���?+�<�FR��#��p����A�6��Mq�ap�_�n���)ֆ{HJEX�y��Cj��&��6e`5�0���z+.��/o���=4:��@�^��,�.�
=�1M�|L���g��;��i��Z ΒP�Gp�Tjb%]s��w�K��1�o@1X3��z��jU�a�m~�n���-��BP˧}��К+���@8�k��� �t�8��{@�HƔ����A�zE6A	ni+c&'f�If����ڟ?�ؠ.�ݍ5ej���j�{��xO�Q��M��G����h�MA�x=�T[�J�������C��)('W��0\�#�QDki�J�O�ll��h}L@m� f�gN��a�B�5��cn����߃�l��@|u�
�c���_��mӖ�+xh��`E��i�^�ާw�Ao�>G�4^���9q����-�mU��J���~�ņ��FuV��qzcNTb,�L8����?cx^�Kt��}ZK��Na�tu��
KbY BP1����
A�:�T]5�"/�.NS!��Z�z�8�d�c�r"�Y-����k^�z'<��w�;�)`�0D�T�G}�N�.?��|≭�Q�3zԝh0�I��Y���ĵԓ T=�!�uX�#�G� �Ǣ�1*LB���ɣG�n&�F�E�/�G���S��Q����C�TY+� l������4��+���g���`3~�7���=�,�L���iU��0ҍ��_�����Ya���T�����U�u#o�d�v�jդY���� C]޹��j�v�a����Ӏ9���͡���-�9�`>��W� ^\m\�<��W`�vpgbauT����-�� ��[q\�Z���ɉ�x���������]D��˜��WB�o�k�ޑ�t�b�Q�<P�g]C^,�6�E]f�4�[��*����_
U�WWջ��H(FF��S9$ba�}I)6F&R�ד�5�|I*7�W'��8�m9I�m��}�a��CM��zN�->��h��&��*Zu��a���W����:4�)����]~�	��D��afW!"1s�%՝�$��}���^���k�ixG_mXl���5�oyF�P�4L��_~a�x0"��o=K�C0��̏i��Y��d�CFU:�xd1��k�qC���a�^$T����1d'$�~���{��Y\J�<R�%�b��Ҕ�?4��`��R0��fS������7�8I���$GRI�\�L�,D���vE;p{�/���:g��L���4oyb�{�ݨ�I<���ͨ	}��\���dl����k�\mH�UO�t7�=��js}\�.[��q4����F��OKl^9��ذ&g�R�Ѥ� �g?��$�1#��z��w��0����R\�*�#�^����w�s�#�8�^���8��tn��
�����6	�����ӏ?��C!��([F]:8�voס�}�
���9�W�m}`�t�,�D�h��TvU�Z_S�4Y{H�^㚳�2��Q%G��ϗTZ�]�pxi�P�f��Q����H
��pASC�&�J�����^G���������j�<K�ZعK�q����������8p�.�>���M$�ڴ���d�(Sb-�f�ܚ�^��~�)���/��Ž��Έ��1�*$ݖ�����K��U�����zU`���Uk'�*]�`����&BE"E}9��#I�>���=<OUٍA\��#b��=�bb(n�R��[�jP;�~�	5�a ���<.��t���0�{�)�2ڼ���u"�,/�6Z�3!�*���\0cZD�� �R�������{��*P���ȩ7�\	g8T ~+~�V�_+J4��&��8�Z�6���k��gvms�鲑��gN
T��46���6��˲`(zW��j���-�>��1(r:���v�S��D>2�$��&f�4~[�LC�8�E��K�ӤHuڅ%�X҃��P��9�<������g��x�%'\��WӦ��Rc�T�*̓$�����Ȗ�l�
�D�+�k��F�T�)���f����s����s�Q��e�5����j�K\CP>���~i<��,l�q�ya�7��b�8Z���"�ش�!�q���ru��X�乥A0�B_�I�P��w�ͨ
�TbGj:=���#e헟�t��я��S)�j�������k���	�"�wE��?��Z�%Z[O�Γd���;��yZi*:H]O9�^�!�;+���y�L@�aH.�qrq������gp�p��yx�0��)/� Js|�r$G��1#�ya�M�'�)��DID�������sL�,Muj/.��M�7mD4���:~ľ���M�3@���6���R`�˳�XSv�D�(�54��*�hZ*�r�&V�L���,(�sV�+*��j��:��"o���#%\1Gڟ�z��%��a�Kk$zsD%gk)b'�����χ��|<�H��,�&��'��Uc�T;=���6���`v�C;|�қS>{*�����t�}���>ֽ,J�(nں�,r�#̨�Ћ7�)#REWaPeL�FH�������û�$ȫ`��eC�7a���Ts�\�ү�������u�o<I��#�`̔ɣ!}i��ژ��C'e�Ee/�}�3�n��x�p5�)��#�!m9qxaX�@� �:��$�3�=Z&~)��1��9�at��0g�n�5�>{�!i�*R����{�*�]��V��������Xd�-����4d�ԊYҐ.7s����r��s��M������߼yW޽{���n�v;�1����U`����d�ؤc����o�]2s�c�PBЃQ�a��G���M��P�}���U�KU�sy��^�2��R8��9=9��&��ޏ�M���u����n�=�r�4�D�7=���!՞Qg�0S�O�{�1O�!"�B!iq�YP���������{
��2x8O`��ɑ��l��g��=�E!�z�M�~������fF��!T3�m���)�B-���<�1�T���)<g�S{Yc�Ve�n%ߐؘS:QMS�G�uӴE��w0��YSc s�D��OEP,��ż#�$��	��Q,��`��X|rk򆬚#
#�*2z����ݤ�8�wX� l���׍�bj�GD <k?&�'�	u�P��7��d�.H�D�Ti�*ir>�<x}I���ZiI��;L�{
�pѠ��x����j�e�&D�@݈�Є����n�Z�Jnn|��S�1a���4�F���"����fJI8��,��g���Sm����u�I�i�����b��k�Rv�H�)G�(�Dѷ�(�Hڮ�W6��#�-i�0f2�08�b��j���aL��G�j^�(֬4NS�Y�n��N��m��KqKm�ܓ�����V�fJ����",)]h�@���`��sS��,������O��3�an��2���>j�,�7 ە,?+�l��Mx��h���TH�ӣU��.���!�.�A�v;���hW��G��lB�P<7#�׏(H5F�Ɖ�^�����"���W_H��5�(����j�6�>���Ԋ��ʭϷ����z�� IPWU]��e#�ֹ���>��╊2�(}^��=o@#���R��A$d �`X�y�ɕ�x�C���u�zY�~��7���FZ�,�t���/^�V���ܥ/�����(��8�"��.n��j�kH���v�9�W�Ţ�MD�tt�Fi�&���F�?)�S��"��:��cv�]#����%��m��>,�S˶mR�`��	eS'@�4�us��ɩ�:�ɉ*#?xD��D%>?5wy��w�gP�0��a/`_��^H���ui��y�Kd��r�;YHӓ� hR���E]��~��B~�c����oֿ㐼i��2qm+�l��Ş	��*l�a�+e��.�E�r��\E/̐rF�(B2�����3���ߒi��[����>��GX��~F�)��䆰���#�4X��\���s>y�>�E-�u:�~ly�&�����n}���7ߚ`�w�}g�
*���zy`�֟1"�l�_|��Arc�[b+��'q��7��ESt���W.i�E��>�4C�ԍ��u2<��~��#Efs.��$C���YB�����ɉ��V(5	E*��Bup��i�������D�9��h)�FW�`�+��\C��Z�c���*c���R7(�%/�/R?S!���,&� �_;ۧ�ŦN$�{�8-Re���&���eIU l<��v�i�p��t��$ں�<y=��?C�4�a�����ԍًG'��й3��x(�z���(�SSW ︁��U�蠒3[<B3�p>[�I���ûw��T*8w�8�}���@C�s7t�����Լnj��=�W=m&Q*�����:��V	��H==�*_�rtu90Eh�8k}�vX��iܤe �8��6�F��^��������jE�}x��5&���*,t&������z�HQ��6QΖGF�/���juX_����ܐ��C'Ux��*�s��ѐR����(�J��j~����F	�!C��(|^�Ф4'm��N���.�5���)wj��g:��A����iDo�w
$����ِ�xc���{��Rہ]O�Ȳ����[���(W#sXP%.[���u-"���7����"�\2+e�*f �����9FD�3g��NMΊ)9��6�x��\�2</
�R6N�b���=�Ԑ���ċ�tV��I�rfxD5���V���j��o�:��Q���� I��_.�H)C���J�h�&��*���	�Tl�JQ�O��Ε�����Nޮ��3.E��z-R+/M%��t��ڸ��<�u����n���.-`�;� KX�$��6ý~��.�5�H#��H��֍��&��ޱ[��,�a�R׵�P�g�Y5/κ�i�)fŽs��U[1�|b�j�J�� q�6hC���60*�-T]]�wk:�Ť�9��k2D��J�p��X�̬�k(�]S�#>O�ugN�|�<]�<��K��d��·�PL��0�����mp�`!�U��I�	,E��eq�2>s^�=��H�'ߧF��u��5�;����5�Kma[�X������z��̩~�O[���4|���5E�Y���h=�ͷ����K�t�
�����9��c�*�9~�^�]�j�T���F
�oJB��.{�J'?`�c��E7���5.�k���k��uL�Zw�~��Ee��9�FVv~��ܥ�(�Yr�th�y�C���:�{}�2����kae���W�`�م�ŏCtß�}m�;�Fѭ+���*����X#�w1����n��yCJ�O�A�kt��(�0٦�['@'�E����6����M���2�Qt�(4�scQ�q=���#z[���G�fOC*��������B�,]�r&Z�t��8�I�h]���T=� ��Gfsj�AU���`FfG71_��(	n�0Mda��2o|v6�� C����>9�����7��5aM��u/�Lf>V��9��iۀpp�m�4�v��D0~�j�3k��it���Iy�U�	����U@�&���>3�ɚo����_\6���?5"ޤPXŐroz����w���]I��m��}Sy����/Ν���b��\a��t���v���;W�ñv,�;�C:9�>� $�4l�,I�K��ܨe!��qyXS��t�n��ϑ�*���q�$�9a��!�����F�+�	��v �I3���͠��w��w��?���������h��At&fD���6�f�#"0C�ۯģ�RJNc3�w`���Å!��?��	OXQ�h���^B��`R���vTP����g�	0p=ۂMD���2������Ed��<���ÐJ|EІ����߫7O("�g8XW�v�0��L�¯S�T|UF�]��beh4	0{QA*����o�P�Q���,�����tV���\�E*��O������
�짳���8�%G?�\�>`]-
Kd-���0C:Q��9��^��mH�N�YٙhH</�g��P<S��V���Z6���wCU9�g��	��:і""������e��l���tM5}�>�sC��i$(a�����x�K�V�cDL��ؠ��T�T�¹���#�>�����x*=�t'���IC������vw&�l�-��:��\�NG�GS�_S�k����u)E@=������&�L����f��Tv��}���%�T[A��bbQ<ĵ�����&� ~G�����ɝgm=:�KE{�C�.+�=�Kr��GQM��8��mOO��8�߯��5*�����{	n++���������z.\���Ɯ��T�.c���MZU�3��8G�5X1���ZMoo���I�G*�a�OKy?�F����k�8�U��z�qΚkh�j��w�%��)�`��JQ�c��ДAm)L5�Є
�Hgj�sxP��H�ƿk�2*-�kDj
(W���IŦ��|�C8���ۼ�J���:���؆/`�v,��Z�r�Ar���w5dK" ��D<j��z�"n<i=�F�W���8�]xU��H�T����+-sN�䠹�oa����hm�
ޅx�4&�{�OPT�_�v�7���9Q����SdL��&�֩�K�|�9�:T��r��Q�\%Hѓ�kFUK�K49����%�&��v�a�^I9_�-Q�O��[X��f��˚�L#�F�m�sV�y�m%�V:�4t#x���'&~^1��Q-H�97���r ���l�{�])J{F�<��۷A3�uύԕ�H�A8�gkrr!y����\޼}kFgS�7J�P'�y�c��ɀ�T��0�x����Љ+�)f}T�~Op^_�������ޠډ�u`v@��߯����˥s����s�r6֧ع���܈F�:&]>a����!��y��F��>u�I]ʍ��ϼr�ɟ��H#����5EH<�">�.Լ�`���.�f�D�z{ĉ�G&�� B��!��6܇�gG��I�P�����[��4OQt�������QJs�n�X�zG׍��߫�՚���U�������J8d��v)Mᐁ��k�a-V���>(=u5����d�c9�)ءt6���F����`-H�i(N;�2C�}����יS_��jOԺ	�����Ë�R{�ʬT��lƴ������'�����l�����=�SoE�38E�6%��2�$���`*d�����C�M��+�K�jB�u���i�lL]X-�=���Q�u0�oo?2���#MJSt��e��n�T�:��M��&E��i*D������Mx�R$̞�����>6�u(�����L�unң+�o�܄�HY蘣�&#R�p6K�Fb�H��yp�Sr_�ۍc��.�Rb��E�`�pY�H�a\�A���7B"��Hka
���0k��}���-�W��W��Qh<�v�"�:�ͬ(T����:��`I�n��m�x&"YTt�����������훷A��\]A����﬏�9�F��"�I�K�\Έ�*��ˇ��_ߛ�Tt��a����������.�\��;��=e��%���d9�ַ�{fN������eLy 	e4%G_�}��>�;ƸǠ�;�r=$����Bm��~�9Q �^{��믿�b><Q�����mo�>���z�J�sAD���u�W�g+�s���8M��z�xI	��#l��o�L��j)q6�x��jr?�uKo"�E$�k{�fE���zw�{S�P�d+�2���gt�қ�k��^}?��Lj�i&.����hty�_5V�,�����7m��%�ϩyi�n��;&Q��%������j�E���'��k�`�\E�C�>�JO�=�H�q�@����v1ي;'�	$�u{�C�բ�yd�qOoh�M��S/��hT�K����U�p=$3�`>���1�N�?ygx���&r���.�I�M�n]#��u�P�3��iZ�N-KC�(�"'<��<p���,�Y�����~�������60���5q@Ιm�HǓ7�
{ݠÒ�B�~�c�Rt�<��V����.����(=����ڥ�����{��h�y�u���Vө�>b$f[6�I������Xk�3��0x+wN5���v�5?*X	�l�z4�SM;��j���a���B����(~9~��'�4�����?%鏀�(Z	#���=Baz�0�nlJ�8���n�,%�tK� ��a|��h��ru�Z��aQ�Q��� ��� {)��76�ҵ-ʘSM(NC4v��dj��}��i==i�H�\FV����զr\Dvn��C����E@v>��B�D`@Es�5 j��q\��HӤ8%j�����/0�����՚�,���ѽ�R�_u�\�#F͡g,�"����^t��O���q�ށ�u��������+�"g=F0d8�QzM�j���S;m!�9�YB�W�o?TX�p\���o�����z�zF�2��A�����N�VU���[�9��T2����Sݟz��o�����|L����}�j��O� dJY@M���f`z����Y�Lg�p�D1.�wTJ����G��H��,�E%�
Ye)�y���K�W�����o5�o����ٟ������Q=#�s��rY�����<r�u���$���!�GO!��Մ���`%� C%`�D��u��E*��M��SʞɳQ�f�/�4��w��S4qPt�ON2�~���ߣ �۽��0}xC���,2�ϑ�xo��� ��E��&;[��Dn��tY�9�ay�*�&�02|�,�US<a���6Jt�Þ�j�틗�i�:Dw��`�\^�o7v��wQPI�.>�*��>�k�9��!���K���E��u�{YG�E{Ƣ_��lz���8F��C8]v9�X:�}L3�N�GFቧ-Q]�<s��2���*~j��E�h���)�&�j����Q���:���VD*��Kij�*���~?�:���ו��$5h�p[F�h-�ߡ�V���c9�5J7CC"���3�b��R7;��������N�ąz��g�i�!����Ϫ�Yy����|�@ߨf�^�&͋/I�(���� z�zIW.�W�#��&�9Q�����G���q�'7����D�D�Y��Z����n��Ɯj�T�^��q�[��hX�^S��}��b��MQ�H]�wRJ�H��z{[$����h.P�G%��ɚ��ڄ�ňj�NC��06"��l����ײO��"�R�4@A[�����i��5�X�_�*�ީUT�G����o�%ǖ�g1����{�L�<<O���,����<JE����)i55M)�,x��l��\��:��q��4��,�s�ZXfaH}�� k��v�x�XO�&�g�s�68ǳm��r��NٴQ<2S���DtM]w�:]��q��X�3�63{�u�?e����F��垭���\�-��B��M/�d9�Y�s�t)��]SqƖe+��')C5a�M4Z�'�Ƃ������M��%~���h��� ��%�9���C$���BUY4�)1��铞��[�x��MDjyӺ�Gc2��:���=G	K�
���^��W�-_7@㇞���n��uD�@��OܹRmNimf�~����!(F0�8t8p"�S=��n@���m��}V��6��\�"#M�4cǽ��w��K_$���!���,1G�.�Rd�Q}��'�N��x։R�}�����Q�Rؙ��|�)FO(��i�@߬#%u��3c�"k<�N_�uu�4�ù�����Z�d��8�f֬#/R�r(�^K,��P�gp��� wL��J�b��}�ڂ�i?�1���9�M6h<6��&�53���v�;�7SZdnuV8�T� �EMdQ�yƵ�k&�±�Q�����H:���٭���>�-w������)L������?y�%�4��c(���s��9"U�[{7HGp��%�g��Q8�a'�ǖнύ�h�cڃ�Gm}g|��A+8����Rlo(�?�R�nLU�Tj"7�lz�t�ٍ��!z�h�<;��bw>K�|P��6 ��E��Ř�ym	� ���nh�N׀dw�%D��^���wvXLKz�t
����Xt4�(�ag���g���]��Ro\����XO8Q��9G\��EN��&R=��a�x
N���SVz���..N�G]��7:g������5� �Q����\�W�V>���'iڀ����Y\��j��޳���l���oo�ѡ���S����-��4%pu�ۄכ�Fr�y��~4�ޭ �ܺ��<��B���ޓ4�t�e�4�ʻ
eH�Qк��H�U���[����jC��B������T�4܈�^�ʘ*������"����M�K��ً*0(�b��@�!"�k,�@q}&W��Aw��mnYq��u5�� ��Â��8���<}C8
��VEJ�F��ܘR]h������G?���&��'p{�kC�8՛�m���$��p0VF�3�!�5�@��`�aP�T��ϱ���)�����$�"@�` 8����iNִ)�7���B�HB�k=����-^,�s]�v�g��'���~{���d�ɌB�	�	Eӑ�6�{���Ģ���=�j�8o�f�F�Z� �K��Z"��]�W�QG��X�f8�1ǌ0ҿq��G!�E�J�ܫ;6�8i 2����V����u�ǜj{�QM�1Ѡ�i�:�9Px�Lk�ۇA�����dkT3Ar�_�X(�$%���9�0���~�H������_�2J�
f�����L�M�wM6�|�F�xf:�l�_�@U�k��	�t�n��������H�$�1W���2�R,�rI�_�eĚ�����-�6�����WKl���Sy0��i��o�ug��F��^�i��bG�<`-{Ӂ�qн�l��K�Z�VP� ��OA���o0F;E�s�'g��5 L�BQ�H���G)��"-a��'(���-��{���9��g�*�o���68L�Y��&�1q�o�yw# �,�㜪p>/C��-:���u����$ڽ���_8Ċ������p9�.�$�����d�
b�6�WG�ZO�#(	G�SG#���!����;p�e����ं��5�����#)y�s����L��7ERM �{i,���_�^�j���C{.�U����Ft~�����3Q�v	��ȤaI�ß��kŷZ�7�vG�{Q)?g2�W��ƶ���_�v����m�\��`��P�G�w�q�h��.�[X�� �%��HE�xE��e���b���M���B���x�����ݾ��
h�OlU�z�x��Q� G
AD�SF#��q�}��;;h�?,ת2�Mf��B�/�
/C�7�r��~K����]�'Fp5��I��<��r!����)�]	��ީ��SY9��
%������&x���wC�ʽz�Ma�#�������ڇ�>���ѡ
sϮ��l���Q\��V�vJv�L#��$�ڐ�@� 6���	��0����~��fwއ��g!lp�q�ǴS����n����lE�Keh�Cʂ���F�h�L�� �1�V���J��֣Ud]?��c�l+����k2ٯ6 �a~�������#��%���O��MR�y���O]ǈB/��F'�"���%��t~��.
�9|�Q!������f¤�����$�3�t.�ն� �5��JX��{w����UC��-����))>��cH[z_�Η͍6��J�KvO��%���{��X���hz`��z�;/�ᰙƦ3%x-��y(U�����L�l�w7'����ZL�ٮ#��:"a�/���Kͥ4�ML�$����d�/įս��O}p�˾hb)�s��ud���.��a�u�S��.�&�#�·��{��F˴<�^zZ�S����]"�bRYک���%�%������ A��׫N�� 7����ԝ����L�p��.��Qg@4%8g\+֛i�.����K�1���5@��3�I���N�u��}�3�~F0<��X?��i��I�1z,�2�4�G��j���#�GƮN�e�j�>��T�tY>��T�풜8�K��K�^�����|z�ҵ0~���W������H%j�8[	���n+UQf�8I�5%�s(A�֖_�}�%�L2哃��}���������߲���^j�M)�:Q(��I:l���i�TJF����w���Q���m2g#�i�Z7f��8F>�<a����ůA�ۜ�o�_��D���c�f��)Uw���(@�V��Oc��n���:EI���������3�?�#�>�=��Z<�t��D��?5��|~0��$��QG�7�ԴA?£��Y��>O�<ԑT�i�g��r�����QpSS��Q[H���d�y��T���K"PЇpe�"��:U<aer5u�뻈�Ek��:y��H$�<g\�g�������o��jޭ�LJ�4M# ��R��h3Ϟ����Q��u<�A�Q<�T�tC���P��0��,g���@��CFimt��B��vpp�]�z����`�l}e�ǋ�r��(��)�cxwp�TT���%�&��z����H���������b��� ���ާ'�8��UU��Q�]p�$d<�)�����o?��E�~إ�ZD��c(�_.�s���T��"�NDp�H��j�%q������j�7qΝ���]lQ�*J����>�='��`KPx�}���	?�����c-�n��	9�������.+<�v�4r9-����������?
J���Yޝ���Ϯ����G����`��u�!�c��⣵��3��vf����l���Ƥ	�V�Z���4E�\���պϛ����$=9)��	��\��Z�uO`��;����f���І��'���O<j#��'�I�s�	��Z��g]�Q����)�I%n\�L͑�M���F3�iDJT����B�mkH�Aj�л5��uU%�x/�s�66W�6OD�0��!�,��)�lE<YzϹP�0�����5�8c��D�y�i�J��ڄz�
���0Gf���[� kPo�+1"�.7�B�O�&#�E-��j�� �ZFΪ0�)���e3l�H��$�b-5,u*���%�Ȱ/&6$7�� �!�7R��=ͳ��6USy��9�1{|/���M��y?�9
���q^°��&(kj�|=eH� r��ۃ�Ꮟ��o��7v�9{�~}]Mvǿ^Vߒ�l�7��m+�~��_S�z�����<;C*To�u23��a���n�(Q������ʜ�N�s�s�F՛�n���Ҁ���3�Ty�>u��R-R�	��a�^���q��Z�c[)����nw��9�8����Kߴ0�x� Ȱ71�%�,<����܄7Q��a5���N)�N�\�hK�Ϳu�O����z��3o�|0�O��������!r�3�F��pF�+�H�]$��������Ǐtalp��Y>d�J#	�-�k�}���C�/#��;�Qp�%��9Ei�FS���v�k����T�h8��8��4���(���!�9}R�Ӊ�-�K�7�(0��O%�gb��R]��~��4�&��ۯ����T��ȏ�?QyB�sۦaf��o�n��J���9ʊ��6�3����&���6��0�Qh3�~�z���K�L��+���>% �~y˶����1"�q�ǽ���c�����y1�͛K��}^�^"@��"�t�qj/���J�P�MA��ee��O�w�����g��Ŀ�*�@U�gWO5��O���;ǒm�%#�q��w)>���s}T��{]E�Qׇ0�%���9�	�*3}uq��fT�-�Ґ�MV���ʏ�.��L��C���<�ɣ��*�"�7i�"9���p�
9s�g�7�8��WE�*�ܔJ��ٙ*�TϚ���q<K���g2��A�ѝ�爵�`+��Z�P%Ew���	C��\w��#&�xj(Ǡb�al'���.�zȂ��<`Xe��T���>tK�,��~�Iےv�M�-ɳ���Mq}LU���0�\�-�g'N]g(�:u��.�`�0� T����_����N��J\=P� ^�z�"��d3����#�/Q����OL[82� ;���Y�F�	a��T���	��;if&����-���3�Xp�����4�`���,�2<k.S������)�*�b�{FTPmxEK�U{u)L^�Z��%��=|D��W�qP|�'^6�z͆��e
�*���d���PK7)�T�kէ4���H�0���o.�ei��UZ�Y7!��|��3{���P�d�DR�_U�W�D�-�M����[lVK����>'"�2Z�s��B ��J�i�Zoٓ�}�6�qW�-�N��H^��Ud�T�9�;{��5M��b��9>�0`
ҩjI}��E�A��z6�!���]t[�
�C#qev[�I;��_�εcw�p��=U�l�\԰A|�$��O����:ͮ�����瀭x?���3�F�p?��K���u(�۬!����R>ru�^$��j�����8@v��j�d�TZ���h,���Wg|�̯���{~B���	'%,��麇��Y���R-�[F��������޴��h�?2>��
:��:��A��hF&��s{���A3�1��ʐZ��EҼpy���Fc��t�v�`�#e��C¤rJ�VQ]GJO:��T%�oɶ��{}T��J�(u��'9�M�J>��ݷ�Y:����?��MC�<FE����պ^J�<�s���q5��y��KF���:h@r�:RCNI=���j%��ؼ%��,�4��11�n�,H)�Q"��g�����H�U���i܄$	3
�Ѽl����É�ˁg��wx�h���S��&� !L5]�i\�ͱm�Z�_jE͙c�{g�,�Y��:���ј�����KM���¡T���M��ދ�"��:7���:�k�F�uWזĎ�TZ/����k�kшX=O����󽋀{��=�M�,��s��z���OG!���ɮyy�dޓw}�=�+j�գv:�t�/��ܝ%T��z0�?����z'�@)#�%��C�G0����2��R���P4�B��.��9�����9f5{J0N�M�Q&�^u+���;K�I�
P��d�H%j����m��I���Eё�$�n��#/�8���ީ ��N���I���0Ҹ���_��^~n��,��a4�����3z��]"r�F�9�˿����8x�{�6�w<A�!�w������>X{�ٮ��q�5D":J��l��� ��WF��' tmU�-/�aQ�ܸMj�hZ5T��b��  ��IDAT4��mk�ŮJ���k�7BP����A�Ǝ;ͪnFׂ;����6-����0a_-��j%���.iM(����*8�Q!��>�8�b%�L��"u���H}�-���'��q�q��]W��#�T0��y��ѯ�랍aO�;>�%�������k߅��1$
jd�Ց$�2��鰧�^�s�T��0TA]K�8�Q\b �T�(|�� ���Wm�%�����.��ܲ��i,%
0��b�{�s�;�P2pl��k��f���|�dۙp�z�M �.�a���H�N� �韪�}��<��~~X~z�8^�y��(E?vm�@������?�`���~��A��ң��7}�b�"m�n?O�-!��:�X~������ǋ|0\�O��[s�'���ӈW���[�p\u��Iő!R�\Rw2�pp������6�%�7��}ui�R���
rⵊƣ�B������n#��,8�bŏ��3���d�w0��W��&�2��,�iGW��T�C�]�߸�J}QɗcA��#�4hN�62�Z�}����|�s(�*�)5X�s��I���}����E��@j�RĆ�}��.��*<��&>����}H�'���1a���`oj*��*d�����|z���2�Ri=5I!m�c�B��A�x��!�-�Z�B�ߣ��|6�9:�8���0OG,�m��cr"qs`LΧ��A4.:��x����-߸	6��)�r�n��0�go���33��ݠ 7�s#�|��Jd /;�:�0� D-�����?	z���I�U&��H����!y�����p/�R2�)Q^ߛ�'���f;@`�%�-�5)sq��F]����hb�-�^�R��fs���*�/^ܹV����qP��♍�z�%m�Ѥiq:ǵy�k�iF��Jw�d�3��?�S��L�zq���w�H;I�[A`쯓G�Z����\�qC���'�~Xm�R��W�t�X>A�hu.�7�7b�hm�4jd�����~ľ �6T�q�^0��c5�2��T8R����x�1�*�\�ݰ=�!��:�T��EZ�~9�"E���S8[��a_����-N'=ͦl`_�64���E��R�;7������!�V�RD��o3p`�900��8�V��q.y︙[�7o�2s�A{�6�6�`ja�7zt�,�`�ĈdP�9�8��B
��`'�m ��I������Ui:���s��3U�<]�ݙ��~��T�JQ�ka�����T�b��"�3��}�2��Q����޺!�3#)�)��gg+Up��q��FV$y���?Dz�ͅ�U���sBYp;�=���P��w�W"Vqi�4V�j�K�fR:]rb1�!h욵��Qvkɭ+Q	��B3�[;��B�ukFO�S\E�u�pJe0�˸�Oe���Z��l=+B�tZM�Z�ި!J>v�}�d{��+*Z7�"eFԴFO4Tl]M�c�o7G���c�gm���~��:G���E�wqI%U��^�~�L���KL@�5G�)*T�S�~�o�N�kj1��umH���
ֺ*:b�q>���6��)"њ�V� ��* �'���1�G��D���S-�*\<�G��uYс�m�����{��=�1Uꖔ����y
�N�<�ͫ��L�	�:� �`�'�x��G���8T뾼~�:7��f.)h���'�!�X��O:E�`*���=��S���n]��j���<�ڳ2�,8!a3,�H)}�T�x����&�>���Rt��0�	{Rt���p�g:��(d`�
���4m`�l�uE-�#|}�Ā訚(:c�*|^�_����n����=c\�=�#���7{I���xK�GNn=X��{��z9�yt^wA1���E�iT�K�����NjVEZKY��S$T���CP����߸��XO����v��Q�tcϧ(N����P5���{5�(�Wǔ�6;����N�Κx���K5���J�?�1��cp[GQ$ڼ��j�:�LҽJ�_]��F�"�ʺZ��o�)���h�Y-���[����2� եs�]�a�nXM�O���=p���׸����w��h��!�ya��Gћ�0�φC&buM�a[<��'���)'�yL`0�H��X"@P�4<b���Z�\L�e�}�ͳ"#�v��S)g�$a�d-������օ�лX����F�C�>DǗw$Ie���ޮ���?�bUo#W߈v���3��f��/�Msblո
�'}�Aբ��m��M�t�6�-.������e'�E9�>�����y�G��֜(�T���)̢�"A�&���1�[r@``��W��!C
c�lAJaj�Etٵ��L��`_�-*���`H��jjt��0��U7Q��7;��/6��Sb�yA!i��x�j��}�2�]=�WVC�r܇�\�}�{������[�]��^����*e�I�4�Uw\��N�����L��ij_{�0�S՟-2��@��"�lϼi{¥ψ�>K=��ԜeM�EUl, �L��M���J!�X'ۨn���'�����o7�rRuو�YS��R����7�PЁQB��f��NO���&A��?���z����=R<���)6��\5�Ŧ\N�X�4{i̹8�G%}P��4uE$``���?�aF��_~*��߽y�3��'�w�u�"�Sj���k�L�:�����/_���ֺ�@�
�R_S��៓����7��4�D��,�A�U�,��%d�}ں��E)N�3�q76�*j�LN���c���"�Dr��NG�f���C��{i�T�p4�PE��[�}tlT�*:1��
ĘQr55�[�q�3�u�����O?�lq�hf�Y��$�W7'��W���&�p��i�v�w��a�D�/&:R9!�TZs�X45U�'�^�vA����3���8$����+�����c��+&R���r�:�O#�����4�ؐ��z���o��䇗��&��!�Ȃ���}T�=�fZ�~�QR_��m��'�.9o��<e�g�'���,�&�������ތ�Gg�x���H��ro�?��QY(^��4
/��Gd|�'&�x����ޗ\��Y,%�u�%:5���N���Uiۮ��Z��o�S���-u6�ߤ���S���r\�(.�~�P�`a�4F4�-�6�Y!mn�]�G��ꞌC�~�]�%�,H��yэ�QՖ�,k�O�9]�К�Ve�0�����}-~_���+��Ql�jR�5���s�!��ZWMw�τ����{f۶��ĳ^{�&C��*AթR�X�$�+T�([k�`*��7Z3F���?,>��+�3�5^L�Ԟ�;�V�:���M�^�&�7o��a?���Q73��K�Ö�����C��2D@p^D�m�|��Tڿ�G���-�E}�i�%���:�➀�@/��F3��Ci�����<e�E�-5 _Mx��zm
	��+��S'1�=Ǌ
Cw��.�4q��mQ�R<]Lu���J��)oj3mn��!2/�ƩH�xC�GڈF`�j}T��)�n,z�3m5��
���v<�?�(ڍ"��;Í���[��	�k�w���#*�Rv)'>�H���4�(��oQh{�^�)4C�L�5���POؔ@Fk�#�<,�'.ȑ's6��"{��cО�,9�f��G�YzK�ib������W�}Qp�
Ք��a�#�P����T�u���A�V���g��S�k�6c5�P��['��Q("��4�k�}�u�>��V���>�s(���e����x���:�5�3�`�nn���>��0�^Nݠ��˚U�Q����ӏ?�
�"[U��EN�����#ҚF�����
����	'��'͵�G��Uj��# ��պ
�����&�P����kX6����)��asӐJ˓�MS�0o|.6���\���@�x����t״���P�,���v�cQ���T7	6DfA�u��EQ�KL#��ŭ/_�LT\�|&�Zq`M�V�T�T���aM�ؚ@�z=Q�8q�z����o����򹴡�Ak�l�%��F!i;�X����c�oMcN���74��
#��]I�l�	]�5iђ���q5��My����
���w�}�^ue+�	8���ׯm/=X�gp�y��=�;���gJJ�Z��~�����(d�E���������\��3.N�K�vY��������ER��U"m����s��4�Sg�D���u���� �ޑØ�v8��O���u���΋�3[��E�M8H܇ś��u�<ؗ�;�޺�-v~qn���{]��"���Ծi�Ѵ�u4�{y|���7�sCZa>5�<xW�B��8{I��i�3�ɰ��f����PK gO�D]+2y����I8QV�Ii����}vW<8�/yi�6~O���=+�鯻gi_v����b(4b��0�-
��_�:RHI��1�m�~���������x�Y������)K"�)�I�P�F���$��߿{�j�N�Z���o�[��X����Pn��4Z��U�-��:�X2}Ed��)/˛�~-�Z�D�0F4���AiFw�0�LGiԳ�w���鶺|`D������3kX_ԕqJ\�"���dxd#���%[�������g9D�3��|��Df�U��_?Z4*�[׾ꖺ���i��${W��E6N�/�ۇ���uu��(W�NJ��(��mHVJ���1�nHA?���n��Җ,���X��	�8C�|h41:��|m��U�W�%ɹG�H�S̓����4-rp��2Z��cF�����Z���z�i:�2̈K�9D�>+�FL��̱NS��k.3��B
I|\�����H��񟷈�鍷F4j�����_J TSQ)�]�&T �� o�兄�T]�X��AF���Jŋ�w��b�`a#3���H�X �)�o�FIr�)
?���#�յ�Z_��r���(T��� �C6L}ˍ�J<M�Z��R�Q���
_6��B�a�G�+.���n5l��am��i��������Ѡu�;���y`�b�t!h��� ��a����f�����:�n2��6�O�%@W׮4^a)����}�t�ڟڣf���I\:�e�UsV.H��E��Z��������\�9i@J��1rX�GZ��ҬN+��ZJ�;����Y/e����~�)�	���Wb���cI:"#4:]�K0	po�yΩ@��@�4O>�j}]�7��BD�Oe7�l� �O�Y`dQ3]/�{�]��7�8F��w���	��7�U��W8+���X��>�ɵ)��8wW6K���3�[�+���1ϭ��#�X��'T��M*#��e󅅃�@4&A�q��6��ӣ����<&1��(��c-����r`/�j*� k�-Gm����:ڇ�)�'j����/3�5���h��>�m�ׯEc3$a�vΫᓌ�h�q`Y����kQqS6�)c �~����E8�!v.���R$�lֿQ���ه��/�ص�h�D�j������iR�6J�̚꾸�su�OJ�!����y��A��gZ��nQ�X�{\�SB�#>�����q�n�c��g7vX��9��߸����+!���E��{Ҁ�O��I������������M�H��jL�������SJ���F(:����17p\ѩ#6@`���>�n	Q���\{~�Y�ѵv�cipM`Ɯ�%�[�BX�����
��?���0�k�X�c��&~�d8�9� �9���!H�ɢ|��H_���I49�thA=C4,gn�l��A����{rt���=ˌ�J�?��I�O�6M��+P�y��+p�Fx�&�a���t�ibEX�j=kZ�M�J�R��Q�ޢx^��>�3�b���95{���B4�ǈ&`H5�M�;纏q���~�hk�2��� �I׉�@T�߿_�������5H�%T�����B|�p�tɣ�����`J6#
#��%/KИQ<��K,��a=>��#�Y���o�ѨMsN�-�B���n3�߅C:�$��Do=�ų�&��&���'�Rk�Q	G�2;Dg�Q�|�:�h���� y��p5�	g?���oY��L-��	W���áVXb{7��I���=�zX�g�֢S�;�棋oc=�5H���0^T?�b��X
W�����'�ґ;y��č�����5�(�l���58f�����3���Raλ�j�%	�a���XI�fc��X�x��,>��ihx�}LQ9F�;d�|}�*q�#�gE&�I?ɔ6��~~�\�m$A#�D�i#���Ȉ���ȨV)5��H�T���,�գ,��%��"κx�'v��"n~7�N�nð�FǄQo5U��B���Z쳶����M��(4^A��S7�	s8W��W��o���HE�	_S�u�����`�l�VVl8lr(��5�^�C�jd�ihV��&���л����
�m���	�"��m����8p-U43B���[���,��A��x�	��dWX$��ɱ"���j�l]�@�%�0��)[M���p���~��ƻ����֕���:;�T�J%�.";cq� Vc���}X��V�C5KDB)
Dd���<�u?Κ�K�N�f`���1�Y*NĘ���9������UT9�Q�}UѸ%�'�a�Ԧ�"����
��M�g���.�2�(~`�C�m��v�9+u7�-$�����X�%nov,�>����z|"�)��&Q��Ƀ_c�!G0k��~'I�5-�kI�0��0}|��|��󶍍y�,� `U6�r�wC,gP���h�����y�$2�DT�J�m�Ź����cP*�Z{f+����'��x� r�vFHU���C���C���9q�MZ�=���,�]ʛ�o"W��u�������[Q�Us�{Y3Z���`ׄ��uB� ��y�"�����841ѱ�X��Z��a�H���V8r����i�wY����`�k9��) ��5µJ���{�#��7��������?��\)������LC��j`��f ������%|����pv�:��s�UTC��בbӲMV�XW�Y�)������U�P�3|�;ز�MC������Xp�S �CSJ۰`��G�����`��͡�)�Q���,�Q(<W��+�X�M��(�8�*�(���xh'b������})��nY���!UT!��FԖ�j��7�\�w��pPb������ ���C�ޑA�����´KRs��K�@Tĉ����1U���Ｐג!�Za1�~��y1^�<�C ��ǟ~J�^�8Z��6n�@.��(`���V���߈{aN��>Z�]_��SCy>��}R��GB狫�_9n��!{��הs|K6Y�I��{��*���:�\HCSWvζO���a�MU�J[��#�K��	�I����g�}�����&۸��ԩ�fܟl�Y�����G��$�i �EPU���m�󶰏`�O�S�]���w��)������eb��d3�j�;PR�ޕ_��k�5QT59?	��|\]���J�C���p��cm7��W$��lJko�-R����8O|�lJN���
�Y��?�������b�ܖ�h2<vޝ�I'��yӶ��a���j��p�W:�Y�E�1sY�*b�XƠ�yI����+��c*��<"%olr�x���r1��K\Dm���$���Z
�����|r�nQy��!:��E��X�Kfٸ��<�ج�+��:�V��'a�) [��7_S���F7	I+UV5?�;!����Zı��W�Q�!����ȞK��]��_]3@"(l��i��	+"�X���,l׳� "R�3#.TWmmY�ױ�OXMh�5j~o��x�!���>��M�&�>l��T�����iמ1I��|�6k��t�z�m���lI�B�a|PZ>^�3ۻ�>c��|�"%�a����#�*0��b6 PI
Դl?�f�mVp0z{�`�~���2�)�8�k������iB�V#��c~m����*����e��]��qT���4���<4;gU\k��f%�%����0������ �3k�X������Hq���#0�g�FVc�Z#�3�$�*�#�3��Wr[ M�S���(�qJ�8������{g�>��MSo�%�z�o7�<o�I��︑-�G���-F�	�MmeHe�j�U[y�l!L�G��v0ݰ�.A*����@��mC�K���w����`��t�G�+j�61,�AK-wqȰ�~�����'\�x���(���l���'�*u�S���I�\K���I�Wꖠ��sr�wȤ§G��p:�]ﺱ�o)]�ma�Ǌ�G�8���#�Cw����{K���8�5���� I?����S�5E�Q`jRR��;��N�H���g��W�DHm�6�����M�����M�^�ɲ����z�2�d4K��r�(:N���x�7G(��v��*�
����Z#�_�{��*%|�sV�u�9�� ��!�����9i�������Qݡ�"�Q�b�6�{�6d�V�B1ZRC��ep�=�#v��z�P�z.�t��h|�����u �4.�h�(_|��s�W��?zH��l�����KV�'P��bS���m�ҷY�hsC"�%��sc�ti����y�YC�ćƈ�ŇT�����ͺDa����GU�gF����bL��1*����H��j��!��C�����~��M��1R
)�@39�9�,*׾-*��S��%�}:�uȯ.5�9����m�d�ם���`�|V0�ѣ�ǆY<rE�Ml�p~�4� �꣪��!
�x�!	�����7? �ً�2�Ͷ3��[������7�����
S�uFf�S�7V|B�\����m��ʐ`��,U `dwWh�=K@G[0�hu��^f� 8���6=R;3Dhx��'c@�	��]2Ua��� E�N�� ����@�)�<*��x=
G��ĩ�(��@Ӕ0l�o_��^ߔ�8��3��B,�	ң��t�Ā�_��.�TI]��U��AR0���isȈ��6��c�գ���?�|n���󈴭#�6�"d0բe�[�h�����Ы�&�/J�p��f���hc�����1��4��}i�0�q������A�(̬�7������TĪg<aS�ۈ^O���z�*6���;�Do\����6��=;1l&���,%�!��W����ɢv/*Q����7Y��\>n}��!��DFa��^�z��1B�b ��} �q5���6g�9w]\�郭���0�Z�����Rl���?'wxS�]��\������5\�9�u]oonܐR	�k���v@�_x!d�(��}�'�ˎ<�xu��L�d��
u�X'c?�i�0S��VE?1�RPPCF�݉�FOb�������~�߇s�����s�����{rA�!�)E޽gy�\IÊϧ�2���ZDH��4����vސ����4���c�qc��u�ڦ:8�8��~]q�uV�nP���aːj
)���#v�=��o�F�3�p�# ��.Y�% эIUOJeL�f���ː�EL��R�>jn?��4���X�?���ǻ�p7�.F@�P��&0�F��B�*T�ߚ���`���W����xs����Ӎ�,)��y"'`
7���-XBl�BɽGcχ�e�$emX<,]s8i��߿�Ap27���ԓK��*��˘
��H�['�g*e�D��T�6����]� �iJy�B�;�*tKF�˜\�R��w\��6:����$�v�ǭ4.�׽�Q��7�&��DKC$�ȟ}�W�1����	1꒩�g��ӝW=�fwh\
ۆ[7�ZΡ��k��V<Gq�ٚ��G��	���k3���D��Ϥ���y$�"%��/Bip;7�9v��;��H���㝮�wx��t�=6�����w(���=ԋ��%��
��9�٦uc��Z�� �Q-��N����>_�������N�3�EB.�%����M�"����߿cM?��f:X�P��"�J�5Q�H��&��jOTTx{C��6�bB��� �^8��=hc^�i=�O	��sԶ�WmD� �]�q��L}4uR�R�'Uc�)ܮ�z�y�����0(����`1�s}/D#�$�ñ��,����Ԫ�r����Abˈ�S�Č��X>F���9��A�� �[a�U�OF�gK���H�9�������Z%�R�f[�M�5q��Z��O�h�m��ڽ��0�6��Z�zا$�W���T�
;��u���
XE��%��auS���c��燑B6(�a��h�a `#��!껢���@:��d�N�q�������~oYC �A]q���E��k��/����OA�E슋�:��mlLe4��������&}\���=�>f�s��"o\�YjP�P�U��SbO8�M�h�����G̜ A"AK���iJ����Pz�>�D��M칥=���?��7��c�����9tCQ�=��%�dQD֛�)3��/,%���=<�q�&�%s�"�[�̔o2���N�$�,���t*Z�9��9:����i�y3�q�y��~x8�CG��D���b;�yg���]�M���i5�[]'����~�.t���$���^}����1as=.�1!g��Dڐ��_�`E?+��	q_�=�_F� ��Q~\�z�I����P���FE�٢ \��M���zM�홌��_�Ck��N��K7��/�����$��Έؼ��sv�ᵎׁ��'��y]�ជݸҥ�q\���4>��q)���&葺����*{�v�&w����k{8BY��s�2�bWw��^�W�BBA�2&s�r,No�y�D&�P0dF�O��,\Q��^�'\�u�{
�c��Xq��*�;Up`�F�Y�t���PJ�0_vN����{���b�\Wֳ�MPYա��'[���)��|Ύu��ba[F��s>103K�a�Xt�6���1��$օ;'%�#	�PN�ϣ)�\.'Sg���&�7�s�pBmH�0	�S!�6��Re����
7���/M5�.6+�	�A�
ԖhH�����7��f��>fL�av��t���u��u2�aUǛ�X�\:y�t*3����������~o<QPJ�ۈv�#|D��o�;U�|��'"R�Q�P�hkxb ��羿���~i�����9e)�4�8P��/���Y x�S�3�h�0̈JŨ`�Qֲ�9ED�e""}�^r�0JV�p�9B��S0�|����s&������[ߏ�&�|�@�$��8#
c������+�JfM	�$��r���TR���4n}4M�TT:��0w�(�%�6��pWP�P�������v������;��>�=}tMb�y��;��GJ��^~��֣iސ==�k�	���5FZŢ�ʧ��Վ��_�Bը��8�R)D��ܥ��E.�Ns���"EHIX��2GX�y=�Cu�
���j���UŴ�H�6;�u8��b�i����ʠ+2� ˻+
%D*:��a�/67�uy��D-F1A��J|աg���N���ɡ��9Mq�¹���cgѪ��^ฅ�E�j�
Jͧ��-�V�Xa/q1�RlB.�{��_��X���ͩ@��5jl��ã�
��������$غ�j�Cg��q��)�|��(��!.��#*���8��2���ǲ�Hk�>,����E��b:-�/w�Ւ]��,gjx4"i?�g:h<���p��9��1ޤ9A�?X'���8����|O�6��4"P�c�Hgfs���X�3�P�a�����
��?J�SQ��s������{��|<D}�j�}:�P��r�6�$���Zim1A�� �h�Y����LJ���0�n�}C�	ָ_m�ܓ;�ٙ$J�&k>�:$x2���󣖥��U-���S��Wx�[�z�wXUf!��)	n���"��/v�C�1���4__g24�.�|��1Bp)�Pp�EhyJ��n�b��-�c.����&�uq��v��)�g�A;� ��:M8��}y�F�H�8�䃍�Ib("�ӣ����>'iO�u�a㷾�,Es�D)���t�'OUL��Y�Pr�=�}ai�m���X����oo�FrcR2|�`� ��(b)��;a��w������B��k�磳���R��"���]'^v��X�0.�����\/�x��K?�1\7 ��iH��3f�]@<Ț��Q� P�W֔�)����gqȫ�ۀ��ڥ�YcY ��O�A7�~��,1f&o�I8���pu9F�׾U���0��X��C�:�R7�� �p�ܮ��=�ِ���1t83F~�o����Dۯ�x���ch3�WD�H7�B3��f��:np�n�b7]|��]���jS^��M�g;�=*'�8��oKH�Q�:\K�bэ=���.�QJ���ztC)i���F[is��h(�H�V�w���ȓ�2�SP4k-0����֣��V����W嫯��4Y�6"�GO�mF9�8����3R^lVu=1U��,h�b=F_�>.59_XdE�����0��.3��fX_�x�<��Χ�R����zK�pm��,�W��Ӝ������Nmj%0�z(9���:�n��]'RS�Y_��qE�9$���e����=�ɢ!��hWT�ii� e\��۞�M���6�/�u�T-��=���gá�EU��"ņ��+b#J��ڻ!xFT{VԵibuX�_M{�$J��� ���\o�m}�Ѡ�!����_F����ώs#x�f�?a�a|2,�x���$�c?c?iԈ�>U��پ�!�N�ә�����������_�`���ć#'w�S
����zݵ�hd�)"�:�櫔�(�"k�Yt8!��&)k��j@�T�Dzҽ��xX�[�Q��!�F� ��?d�Do�h�@c�s�U�m��ۊmD�GMo��ɿ��FF�{�ٹ�DJ�0�\}߆h+>�QFaY.�zY�hn���l��S�M8�&'�;W�O��
͖�q1�>��p$�J��UOŜ�MN��
�u5\�w5�����;�X �dMS/r���R�٣V���xtm\ҶMϾ0�5ޣ�-->�m��.�wo���D��3��/� C�
7�戀�3��*�~PL���x4��J�QVi�^����mF6����y��Ce�65?��y۾�rx��� 9nO��3��9�0�T[�^s-3�3�	-U��""��6�ϤHI*��Y�f��Á8��ό�~�]��s���
��<[}�䐁��\��)�;-�����3�)nT�1ҕ��|�p'cJq�'�,�Nq��v�̻fs�dHe��O����͙��	>Q��m"�Ń��!��eʠ�m�)�Ti�-�q����nM^QM(��A_d���4i&������ņ����7��l�����3Vh7�����sZL���)����֙��}�bS��|����uF�z%UJ0��Wz���s��B�NU�,��ܣ�HPBX��֩单Q��j�������-�Ьl�}�����읾�qƇ��Ba�:�/6��zk��6��@e�V&:D�R���y̡.��*ǀBLJm��3��S�px������x�5�+�7��=Wx�R#eT�&�7�wEeë�w��B7n^DoF�[,:"���I���*��Fs|kd�~�u�~g�[���J���,-��֛7�>9-[e)�v�3lTWz'Ƕ1(D{�Eܱ��2��Ǹ�u�B���z�>�ds~�Ս��ѓ�fz�m�C�����_��"�1��z����(*U^��uY�!���t}�j6�p)�M4��^����T���-!�e������^��9�sKx��\]�TMv}n/�^���;'�F�W�$���T�u#��BI��M�]�==�v�
5�VUHPt8.��:e��f\���+C%�#�I�]����w���!I�ΑE���%�O��_|����W��OjҐf�����4�H*X��s]E�#" D¯����/�o^ݼ0j�����X�E䅆�!�񔔩�Qb��xf�������S�y�&��:o�;�S#31UT�
?��`}�����{�Z䆩���LD��c(������}�z��ʴ,���ept��T�Y%�Rx�lK�ሓw׭�Nc͡W������d�W�x��X�� Ԣ����w ���*���Y+T�j�;��������S#[4FE�D�q-һ2�S<a�t>Ť� ���y�q���ZM�h$����2Z5cA������5;LR���@���(�j�v�z]��:�Q�d���"�MD�ܘV�PvI�u:�N=�T������S�a/^U��]��PO�Dd��mR�X"В��i2��yY2��>p����\Вv52E\7��)6��7�~kt���֮ׅJ�/��HZ�$�w�."Q��de��C���P�WO�|�-~�����=�I�#��L$P�ը��R=�����ܷ�w\1Ӳ
@�7���#P3�偬���* 32���?�Ǩ��i<v��F��b!ߒ�Z��c���M�*x�ar1�I���)��m�
���1�s��[�Hݳ��K�p�O�L�����*X��'m�tu0bbk4vT|_`�@�K� T���g��$�p8���}��=����㗨����wl=��?��<>]AA�C?��qo���qqc�Yj�1�h����eCt�]�0"�U燤=�j�f�h����l�`M�E£��D���nӜ-�mg��W����~>��!�#rP���R)�������r>�T'� �눴�����[T�yn�]'������3�8E�zw\V��ղ0��4_��Q~��H�C���#��#9h^�iA���c���8e"�L�Qiske�-�1����:z��$*�*���v�.�IbU�!?��3��f�ty(�{OE�aX�̂P�v��v�}��F���m��wv�W�U׀0�eUs��n��xx�i��|\��@d����i��u(�B>�7ǈ�GNj�y�ff2v��Eu�)�� �o�Q�!hd>�Ǖ�[������YZ�-�-T2(؋d>$�JA4�k,J�c�G$!�9&S�RAH�������	9�CrI���1�WP^�R#1����|���?N�ёCl{��-dU�����FFo_�����RH�p�W��8e�������hum��#G�����U�!�8:�X$�Y9� lsj�<Ys�q�)���Q!�g�ɇ�4��uH諗��>sϫߍH��Y��T���T�?s�����i��a�����UuwYU���}���5����#R?�lB�V��^��\���V���V����M ��T,���È�����Q��ǈ����%��%��U���8��jT�H�a#�r��u>=�$ڏ7�r���>/Af7u��hׁt�\Q��>Lɨ�D��,�w��晕ToxE����~иvT��)�?u �Z4�/Tп~�hc�����LL���}b�>@��C���/�\G �껁� iF9%�: ����<�h�]E����~�xh�*J�ǲ�4O6�"�e+�Z�ʦƲ$O4(E�L��d �/)h<��N��pL��YY�S���_��R�-��mXpf�fn�\q@���|���(�s�$�(Z]@a��D�C�����[����U~N��b�~nE�m�]5�XL-��h�4�B;S�ք�1���a���5:����1���S�5�k�(nWѓA���F��}1E�tY��������e���-M7���j��������Q�_����hP����E���G��z5��n뻽%IނN��gF�x��)G�z����
8hU�ӧω]R�L��sv\��]��F�>�C(.�@8��	�+RT��T������wR���9�	0J�g�������z�~���v�cRV@Q436�� �����>1����x<�q���?伣7aX�����SUܡ���q�A�v�V"�9M��4}w����v���	���z`��F&������,zJ�8 �0�������&mE]Y��9��VT#��j{��扊�]_c�f���"o�RCa�sk$y��{��H
Vb�^\a�2�H�7��:R\�H![�]�F�5bw�J5�c|��X�Ε_��֚�s���y���$V�,�g�;�Q5S�hlD�Iu��r��	�mw$.���;�o�:�c�0O.<-q��]�طǏ�jYDwzmH_㺿1}�1��ڭ���!�[�7.���]2.X�E<�8�Z��.��>�-<l���v���z9o��~���|��.@��h�P���xy���ltN2�?d�u<�o}���r
��Ym�QQ����
�)��m�Q['`��}���F=ޥ��Dt�*r�,;"'�����>)�����UU>#L|�6X<�>���x1�V#��.�3#��`{�i�M��p8v��9(�+���|](�%Lxw�DV����1�!j>`q��]�Mv<5��|n���~��{=�2Xm��{w��=4��	�EN�Q�x�q�	�NSCxY���&�����fi"�,�6\Z��-����]c�~������Bvhx���&�sp1���|���b�زn*��Q],�og�Dy��6O�75f�T��ɐ.M�!�xv;i��L��+9z��,C���P����r����*�����x�+�WH�ݪg�#
�|�ɿ�|{Dn!��;4z�.��9mc�M5�յ����G��O���{�_Do�bW��X���N��������X/ߟ����pJ�
��S�)<?62�X=�s�mre��Y8 S�=��t��8�����;bL�.[%�H�6�9/|63`��@������9x�0KG��*����Yl�%6�vд�b�܀14���if���a�	�	�)��������y�]qX��b��Z�_ "W��
qq�m�k�4
Ǽ���ߍ�_ݥ��Z)����ف�E�&tネÍȭipY5�G�� �K��R��n��0�2�oVt��>r�q���3V#r�	����Ρx���o�b?ڡn�a�6(�I�8g�kպ;skY3�] �G����Q���u�K�,ΕQ���3��?�0I_2�v����X�L�ʃX��н�u@�u�m��ZԐ~��n���g$M�W{l�ǆ>�b~�s��j'���1n9��3Z0��)6I㕶e�/���% }�F�&Fa�į��$�����FI����੩Pyҥf�Ħ��s8����)����#�r4�U�$B���!�.W8��W|���m�{-I����)�F2&lk��/�w�Jf�b\0�W�OnTr���Et���������o��a*;�)�f��r�d��d^��}]�����[}��/�jj��(�Z�jH��sJ׭o�(z�kv�c����p��LM���hU�O������
���^�;Ӝ4)�y��#Hj;G���eyz��@���Χs�l���t �λ�<�S�����Mp�{'��Jk�.��s�J	��'ơ梅�) 9c_F��
E9N���_YB_X�����X���������w�?v���@�����ҙ�9;��j'4&�Τ�NO�Vc�P��V�p�l��<����]V|m�L�rO>�.�����J���Ѧ��p��>�J���s:j&�S_K���R��6�~.��X�)R� ��~v^��O��yR�2.9��V*�B�����:�ބr<"j|���Q�n7&-�YEG�Ƙc���dѨ$�5K��P�v�v��90*
x@cVއ�=�ѝ:�.�B�h���J�`=̈T|H�z�z(߬�]d9�&%
�ٶ�)\Q*Ν΁�Ӝ����i�~��l7{�w����4�=���/��Ic�`�#R��߾{�Њ#�V?�i5-�uQ��QV�#16��}�N�^3�e:�`�[F��BdƎ�|!E���g!S\����l|�p�PC�(.����,��B�:�YQ�M{� [ř�ې΂�Ᾱ�V�
�f�_^Ā��n.&�W�I�U�V�e�^E�՘Vkx]�����!k��b�v�ՉQ1a*-�ߤ�J��>M���IX����Ӽ�p�!n�X���7�I
��n�G9�B<��;�Ǯx�Bp2U���3��Y|��3��}�Z��]����i��Yj;�;
��C��S*s��ta��XN�H�US3(EG*�;b�Cr[�@q�)��6�]S,1�oۦi��s;F����a��i`>��ؘ�/ˉ�ա��f��>U�n��Ͼ�-V�����i8���=y����u������Ģ�Ѻ��6J^a�U��c��/��f|��h//x��|�p7�@�S��J֊&y�2���PS�0��b2q�OO҉u���eM��3��k�*j"ts ��5�9IU���^3�"��v�d&Uz��w��a�y^�������s݉r��h�ZT���oݍ�,%6fh�.ၼ#��{��Al�E��'�Anc��l��φX
 �,�̤����u���^S�5�]���@�����P�y)k�[e�_ť8h���`}fOxwƎ�9r����IL	�;�}���P_I7Y�����c��q�e�ϯ�ε��r��G�G�Y��dX b×�����XZl�Q�ݝZ�u��8�0��H}���5&:IH!$����	�� ��������*��:�����>n�*)��w��4i�.��]'cU~�
���˄�\������0�"a��WD�l�M���he���0��-1>���H�4&n Qt��t���Fƛ��uӰ��s�����rО��(%.|�����85ː�A��J�S�lp���Ug��f���N�	N�&j���*;PwO�I�T�w�F��fw؍2)�� �����_��vт���Ye<�!x-V�y��۞=��l<���_�1n��Ykt4��p�X�l��.�����̍P�:#j'dPa�v] ��rM���֠* ujo��U��UqR�]Y��n&w�r�c�y����RT�Wva<<�������!
���������FI�ƭ�&Up���fFq'�&�^~��p;��}V;gr�UCU�}Fۤ�\8e��0����e*��U��3��c�۶�"Ӂn�2��(O8�û��É?�=�#|���>��5��a�(��sF�~����+�:h����x�g�Lp��ºĢ���>�s����U���O]�T�*��޸����(gE�OyOQ��U%&쟣& DƤ�J��%�f7�xp���Z���4[�F�V���&y�!e�e�u�A���#0ȱ5����c]c����}�`�m������sG��D��g6�Cm�6v.��L���&
�`���x���嶜�����4��kE�/��{:��a��56�J�0ǳ �۠�A�
�E�o����Л�7���^81�����1�����`@ciJ]�����NI�v(��I�w�=W�������ujoS�w0�5M���������6"n�j��k`��̘�_.$���zӑ�з�B�S�� 9��)]7�bwi`�bn��I�d��k^_�s���V�������9 �'id�Ԟ@{_��k�撞�S١Q��nْ���:up�Yq�X��g�&�OK�X��P�{�eԍ�h޴b?�U9��l�0�����갔�z��9t��}���P��lN�4zU�T�������F��8W���p�x�Ð��A���Fذւ���eո^b�3�_��4��V4U��;�G�2��`�q�*���N����Ya�����r����{ŷ�,�*Wt1����(��o���(�I�#1"2%E����i�X����q��>�s#~�s�fv�l��f��`>w�EČs؏�~���k�YhS���V.�1�L�jZC|�r����Mͺ�V��J8_����e�
��%0�����3�2���LgGG
"���89+-px+?1j|j��U�������{��v�+�1�_E�a[*�5G� J���/��� ����ۨ��e�=��
)�`���!D���aq;�7+����2O�Gd�X��F{��?,��/�{;ѓ�J|P�����d4r�M��oR�z��w��7���E����n�\gqCa>4i隅����ne�~V!���%��|7ϝG$���y��ޏ��]���zz��,��a{΅���T�r�, �P�z�Q���� ��ᔾ/�"s�Ύ,t�0uQ�k�2��J�oqT��+�����Ο>�b�<ާ�@����L͌��X�b-�3�0���23��Lu_��N8�ԵM�Y�ۋ�����8�DE���	�>�j��"*m�?�q��|��_�:����E4H����:�������G�#B��t�,oc`��l�����1�|x�!�B�P�Ez���u�Ϲ�X���.n�����rX�'�J��ʡ��5|w��k���loC��6Sl��I�"��0���q�nh�a�����RT����3�+���__S��cbf6n�z���p<v �v{�5���.��	��%ػ�z�0���>K�b3������u�Yo�4[k/L��`�Vq�X`p�[�m���%�Q���}��@A�pY�Fe�
N�}�i~|�f.i/|���9-n6�%�)`/D�ls��&�o��
o�ڠ����wa$?}�T>m{��ki��������'I����=�S��:�RQ8�~(��ܧX�)+��	t`]|�ϥ��w{r��_ԣ�Fo������p�
�1�Q�8���o�7a@�//n��]G������I�����) O��e��F�i=s�|Q�Z�)��X�kB�+���G��z�W�dKf��3��P�~:,7��X�䩟���C�����a���ka^>�&��K���iH6ֽR�v�3၊�;��L����8�dE�7�~�X9�]w� �h�`�!�����]�8C_g%�bΟ�.E��kr����#�QY�@��E�H�Y��� ;s�DQd��`�)>��`"R�}��)�g����!��2#.�X��a]I5{HC�C�,��/�(0�:�&��Ո̾n���f��`�R�r�p�`|>qO8���)�K�j��/�K�hg�xK�H�u9_Ȅzg&_�u���J@C\�^mЦ�����n����������6��E��l�z�ܕ��.?��c����?�g<��PB8SлD���ě/U�$x��̶/}�0�!GK��7�Vjb;40Q���Q|�r������� N���&?s���5&+|��sf�9%��ׁ����P~���X��X�����]�N�g41)�E�t���uߗ����"l�������KZ��i�U��X�&"����]���T�;WK�n�G�8ͬ��2�22%æ���GFQ	�8h��E}���؄�-�$�����H��>����T����)������I������^J;҃�7��� |��t�TBG��
<N=<%�Ņ���ValA'��O�:�)��uF!M�P�:�U�����03;�� 
�FH�A<��fQr�Ŗg�]չ��#E�È"����+|����
����((i#�����T2����H��Ut��ɐ<FR]%Kv���{�����wUǲ�#	J�cW��&`�\XC=I _�����x�F!΃뾗��e"����cjCD�E!)�흨%l6O�@���i��b����=����v;�(&ng�$�~��b��!q9+���3���q�]�3�M:�5���FnX�����id����#�^�B�z|րlЌ�}�q/�zM� �Ѯ2d��,��`޿kd+��P����?�w��������Q�����ĕ�0�Pj�QC:z���q"(�� i�;���=�>�L���x^�qXp����ύ*�-E^�8����+9I����i�<�I6��V�%��)��s������	�;n�8�C�̩�ʡ\j��x}Q��l+�Y�of��#�+_��㔅�.�r��x�n�+Hۭ�c}�l���?IpeR'���UA���O���Kd�f�3�(REA����0��M�`T,��͈o�֕p��ƂEP���/�l�y&���k�������Ȼ.g��{�Í渏L�/lB�����_��r�RD��hH�E�1��Ǔ�Mx��y֥��4���S�:0`=�9�f��wfY��Q�<"�h*��!�s9*0�4;��� ��5���/g���N�`C�.��Ҙb��o���Y�������^{�.��Q�Qj!3�D��h7�l��Z �8�p�����Ok���1�W/=נ|�w��m�i� �IU���lF�:Ԩ4�N�E{��S"n���@s������HE~ݾ��A�G܄[�������q��4�K���D/~'��P�׬�ë��E� �Kz��}j���SL�L}UG8��-��I�|�ᨊ���j���_�K��_D�A��C�����?Ʀ�
�f(��l�+e������Et�Ӊ�g�����	���4�ќ�q	0�<l��m���8|_>���?�%�����]n�ٸ2�k��q��	��RG���Ѿf�x�C��)B�"��ʉ�6���!V6�XV�wF�KK�r��^�ws*a��c�
���pDN)?��s���?G ���oL���nBo����Q|b\�ˉ�XOo�t 6D$-
��I��G��n8��	#�$:��Ӿ�����@)�Ѣ�Gq{�P�{�S���sCW������sF�4�k|��� ^���B؋�r!����?l�{NF�y��k0c��� fW�z^ӛ^����M�jO�"�uW�����SU�Tp��o�EjSXY#vG�z72��8ȰEeK9oF��t�����n��cv$��7�s=�`Hl��$��b��U���B�w]ġ����+� ���	�'.<{i��z�JŃ�Kx��ݠ��T�!ժ>$�G�Ѐ{>�7�i'c�|S⫋�V�"(
l�M���>���n����>X�1p�QuE� �x�yI�N���� �y�V+�@�R�3��EX/�.sM�c���'���#k|(b
�v��ḚJ�UZK�k<�]]V&
��w$�� �zS��a�7�+U�T��J���p��g�u�e-�V!)�׹F�cFSYz?��ݴrY�"݀�R�v��g��v.R�H�\Ea����W�c�ָ_*=�g�0r>�G�X��m�0E�cdE����Z�+:����\�$�W��?g�m�K4���ځ�k�5����7/�<Ґ�m��b�ki�����	�'��1�6-à���V�1��`�_n^�R �EL��xJl�7��)��$�����&�u �������E������>���8�� On^��D�oZ�_��9B��Ak�_�e����!���|6""��d���g|�{�	��@�>��D��%��xE�~x�Plڢ%T�]���*������=����}~�EW����D��.�˔stb/�3��e���GyB�a6���Q�̠�.{�Tv��k��Q�Y��%ӮM�h�&��]I�67��v(�C�;��Z�(����ݩ ����mYa~1l\�N���\��E��a/Z�]Ϋ2���ꭃws����0l�����\ؽh#b�`�5��[�Ȇ��#D��b�F���M�M�/� Fa�A8��ѻ�F��?�vlN� ��J��O��0�����w׆����#lGͥ7�0[�i����M�o�%���-��Q���/�9����,���FzG����&v�t��oԆԞ���F?y���M�:�(��z��6��öؓ�z;N\���u�C	#v������?�����א�c�TM<�1f���pU*��;�O�|�<�@���ys��IA�Ɛ�#u�j�f�G�o�L@��xH�.���;���S���Q������ɝ�x>~����XGT�q/HGQh�!6�4"7:�ϱo\�u���k�k����J�P#A��E����m� �-����]�}��{�5ۜ@��\K[���J��{�^c��sT�)*�n>d5��M�Bլ^��c^R�����)eͬ�s�Q9�#�y�£����RY�2�q�LTݫ�3��V��  �s�>��F'���;�1&�*ru��L�4;rP��J���H��"|�48J� �b[�k�	�Q�|g�m���Z�PȄ��1�,5K�!�SDe<�[��ԃ�*xk��Q�2-��牎No"*U;gz��]�Op ����A͠BQ��U%>��y���pJ���o��X��$x{�2��a9G�Dt��C�E�WАަ6�F_���_�%x���o��?���
%`S|��q�� !{����ZӞ��pЁk�(�j&�ć͐���Р���+)L�*
xN;
{6��dq?��_
ǳ|�h2|4����Ѕv����O?��d\�v�!B7r3t�!�������4��r���3�qG����;��k�f*2<1{��y����`i[4�b��V�
�G�{�(�t�޲EU�5�,��ro�T�j4�b!���	��4��`i#Rub!�2}��|N6��||���ޡh��Jt��b2��"o�蠣���T*�����!Ea�T�=W��`���h����j
�^D�O���x��<�>G��p潮��r{�:%��yZ���k����� �F����H-v䂓4G�m���s�*�������'g� �B�.i�&Z���2��r��渉H�/����ɘb3,ul2^�I���V!{%D�` ���9{�M�N�^�Ȅ)!�)�?\Uཐ�춛�� ���q��s#�؀��eꆈ�#�EtD���)�+�"��*��o@4�Q �1G1�aՑ���d�Q��Rm��C�z�9�_���(<�ȳC�����!�@�"`��#ٷ�$�ً�S;R.S`�������$�q'^�slDA_��f�>�3�X��3u��?��|�E�4�L���xVq����0 x��R�NfY�����4��|f��Z�՗)4;��<�@��1#�q�h�>=1"1���ﮰ�0�F�ј��,>�H78�����.��Ql�m�����u����J=�aa�8��.3\r�i��2����b��j֔�a��e�6l3�(�|..�������(�y�4A��U�g���;2�m��ʾ���i1mH_KEU0@6��^̳�5ђ�
!��Ε�˙)ґe�^)۸f��T\F��#E�2��/�����9cm�͕�����?dDk~�!�i�w�P��}�/Yr�R	���0$���t�%6r�QnlP�9��e7��F:m��_J#����F�Bz�50�l�a�I��:��*J�G��B�}}�#��n,�ǉ�_a䤤ONfm�ͷl� l��(����f�c�O|��JLǞ��C����mT亸��5�����
,���(8����aHmX���Y���s:죰a8��L�\�&�{#�[��P�ʽ3�p����<) �h�q��.�h���{����N8��(��(8���M졯�ti���kvR��QIV�*��ݠ�u]���D@t"�}g�"Y�!2l��q��2(Ws��B7�he��!��m�`k�Q�%�����Gп4z��S���dH�ڽ��d�����fa�.�Iy�]kD[>Z�S�I)�GCU�A2=����tV�������g�dc����?����?���9ӀPOza�!Da��D}���JoI��=��;j��;��^9$�\�Ke\9z�Cј=6���1���C�5�
:�V.��^���ǿ!\AR�s�.N�=����x���H=s�$�����-f�G��;9�!�KAad��ܫ[�>Ԫ�0��?��׍�F�T4"����ȢY�I=�v�ϭ�״�N��#�����ݶ�����_��_�l:9��6�|�ݐ��!�֡��\�E�ֳ�FBN�2��Y������
G!��q���JY�]�P�^�7=뀛�ݫ��4�2'*g�i���R�y����(C���BQ!���c�yD;9��B��eI��Vڟc�gD�H�5�.��>G62��������5��rD�ۭYl㵘�?+@��]I����E��%���Q|�}F�-��m�.Q�����OGCZ~׈:��W0s�7�-,�-x�5#d�[Z�����$�k���]{!S/~Kϸ��uN�������h���D�G��TՐ�'��,K�ZS�I��}���S��KL�ޯ�e���a��a����(\G+��tDl��h�z 8�bWT=�R�Z�����z���r�����Ǝ�h���#��&��H����F���[j��$CȗSزK�W�*���l�_�F���D�%��F��F��ؕFM(��cT�}�.���ؓ���U�'6���t�
��}K��\�H'Y�m���k*k����Z�m��m��{�|iy���ಋ4/�Yc/�.&LU�X����l�y^��&+y�17E,���ܘa=���m�#D�C�jB8��LxW���\x��Z��I�������<:�m�>���H�2\�D���	�M�Emb���:尵��| ��'\���D�g�j�s�ܞ�3MU�ؑ�EI��3"�����9��ѣ!Y���AV���Ї�.�_��n�^.�Z�(v)]F����u�sSv�X�
�<�T���u}|�Ȗ!��[͚:)��zEv T2j</u�O}ya���х����Rq<�+*���P)�&�Gl��{%�U�T�-7~IC�H��Ydp�����q��+oo1��#P9Nd�1I�X�RGQA+��l��=�9T)@.p`� Z�y�=]�q�u퓦gV��f��QxP��jpDI��������s���`n�nC0>����t�.�}�WDʤh�l�3��窮�=�K�$��5�35��L(�Tv(V�2s�M�kH-����ڶ�h����>�g�pʄ�I��p����𷆴���Ɨ4�5��)jm���B��A�-��<Nh���;�f�Ζ�xc��N"s���m�wN9��@9�גl�F�!���Z�׸DJ�
,�uF��-�.2���$�Y��r�iܛ�s]C_<�#��$v�b�,���A�1� F���,������'��G*�
�w1����6�BX���|DY;���0�W��/5
�^?Iy���RU����h<*4�f�9`��JI>7j��_.z�q�D������P�=�ѽ�&����Y�#[l��|�w_���l�"z� kd�s\q�h�=5��Ҹ�)E�fRn��PN�@JU���J:��C0ӼK��(����8�Թ��(>�1�����>k�}�.<�۶�r~���mG�Ps�6Ai8�_�J���]��`UU6>Ϯ��_۲��������`��WJ�g5��\��������!U8�5��:�ۘ�*��Ԅ�Jq:Q�R���8�U*���8�A��7dcg��N���R����mק.$C	�t����)5�6��Vc]$�b>�rC����B'��r�h��H�>_�15|6+��J�n��Wg�gv���(���(��a��I��/�K�-���F�F?���"�F�0��U��W=�S1/�x�#���(�L��?��ާ����}*�?<k�'���t6�v�+c�,�B6C��2%u	X7�����"#E��ų�j�	{֙^}��"Rv��<0<>_���G�x�(7t��	�0F�{@����c�.'I2Ml3�����ԩ��8*����ݩ�Mdq�C	~�1��T�uU!�t�v��xiJm���,�͛>�J?n��s�L�oM�q%��~�n*�.��S4���p��|o�+�sF�/8��r����6�`q�R�������,:�Q��,b����~-����G�i�f}E��w��\����پ~��u+�, �]�c.,�����Z�"՝��H�Ý�f��g�n l�N��7n�n�~a�z��:Z)nx>DSa������kf�=��U�)��L��*��_��ѡ��va��;���M*��uP�@L�Z�7�n��������wQ%�^Rx���9B�t1|.�V0��Y������׿�sj,���$�=m�� ��8�(��:)�UQ�.3e��22u�meV�Cd��95Gk���E�t-�rR1�J�@b=�^�d�CR�z997*B�����`>���l��S�oR�5����7%�l�r���.�a�1.T�Z�Jbfs���8�Y��ng���T�^>��{�}{�/�{��g�kF��zz����0	GG'��y�g�V��萙�T�E�Z�2QڥZ#q�l��\����:�w�ŽN�sOS3�Z�mj�%g�����t65mM�b�������B�4�j�����=i"���'��d��cl>0����w��6��bg�>ϊ(f����{����I�*��9��mDt�����}@\�o��ݪ��`��_�dɿ<���뇁.Ɣ�x1F��4X].H�o9>i#*�!T�=����᧟��<P�}CΆ��7Cz�ro$�Wv��O����9�_��"�p����q��kC�M���z�9��Fx&S���t��o�$�
���c!n�:jzh��x��SU�P̜�u�����1GQtzԆ��c,ʶU�igDM�H�먔5SZ߻���N�~/��MS��8�,��敓9�hHG�6�\��)�(ڒO����:���9pp0�v'5,X�"��%�]0]xm5�L�!�w
�H1چ���������c�׫Z	4M�cQօ�אeT�^�`�׆s-�АVc�0�z[C����n�q[K��ʘ�)�uX��F�Ge���a�":���%�bPҮ�H�Y��;�qur�(�����g?���StP��SW��?��gu1Q���D��nݽ\=��V��(�T�H�� �9ђ�ަ�='��ip�H�(�!X�5���-8�n�� ��"��P��aK�1X�N��%6:���	�T���Ǐ[4�׈� �1�ʎ.�acA�	'��wW�5b�<�"n�EE�����0� �}sb8����@��y�5W-5舴a:b��!���������R1�ڡ����8"vZ '��J���GE--�t^�#t3f���}UQ3D��"�5F�_�U�4A� 	�s�cCm$�`0��:,o�>�s��l?�ʀH��a�=L�Ħ
������#��:nu�bC��m��v�5�;�65l�4��J�A��Ym���PV�`�)�Fu׆ϵ�ֹp**�!�
���ZC��������kXiS]z]h��-�T�ƫ["��T}����h����r�0����WX�s��Q�@��W�Es
'*����� >����K>W�	�"�SO/SO�a(	�Yxj$ �nȞa㱌���4�m��G���*��W��kN���Ew���^��zK��T��ZɿC�6ܛ�h]��r���ܣ�k�ty�4��:�;��bR����3�)P�q���J�x�߅!�/2�K�/v�?�le�z]����wKK
��h��mD�Pe@DG�XE�����`��E}�1��P�=��DL�o���f
An��Hs��@��AM��rM\��ǿ����|�@'�m 6yT��d.Ἆ��uy~� K�kz����+#Y���Jڒ�f���)jKhB9�u8ڭ��ud��o�G�<��5���-�vm�Ԭv�qi��b��K�����H�1ص* 9�����L�\*��"�O���D��"n�!:�F�a���}�#�;�]o�h��qxa��~��7.�k���ߍ��X���T�5�H��q{ߧ� P�t>˾�\?EJ���"���@1Lµ���9O�e�脱FS����r���EW|5���=J�7��!"Q��������Jjւ9�A�A�S���I��F{a�n�����Í�w	(Qj�f� ��0�\��Ҳ(W�
32C��E���27>�`A	��H�zpA�R�p��h��ܸ�C�u�$�q�����Fq	�����i�rN9t�����o$�wT��!�xk�m\Lgb��.�z>����p���n��,�L	�\"cq�4
|GR������<vb�1�P|�$x�A�km���e������:J�'��Jj)Q�,�������P5�Kc�+絭�8�
�`��X�V��y8��3W��q�Պ�:c��ν�j�����9���>�8�B��>��m;$�W�Ҁ��W	��ϔ,�HZ��8>kx�S��%*~�]0:m�(*Ǔ�ɹ|��Cy����)�=ƁG�Z��!Ҁ��J4c�%
PV%ꕶ�bָ�Q���%���bHL�#)���b�����<�s����n�^hJ�9��}:�P1�N��oQD
��CP��U���h5u������L*7�t���/�h�kYׄ[!9������Sa���E����70���P�%��S�Wi2%c�1IT���>;�@<���9;�n'}�N���p�1����[�f�3Z��c����%����z�s��[�ä|�0hr�O8'}W������Yc߰p�|-��Il�H黔��5�5�����¡���Q�Z����Լsb�����a7R~�Q��q��3LC���\���{���]U�ƈVVɫ��s���aLCCuI�^�%p"U�cFN/�f�J����;�<��m,Q��ν�:�Wx���)i�R��-=f<����h�k�K����|�%~��	#,,�~������0�:EdgC�CjH��?��vc��8��"/�匋�5����oN���f-a����a
6>"/bV�F�C�a8���O��U��lH�6�JS�ś@$���>���0<�n5�i"Q�l�Z�=0�g��*�2t8G�����)#�w\G�>i`�(N��cԼ��1&��5��Dq�T�#����(��
�d��ǰ�"��J��xg8���0J��L~]Ŭ����Nb/-�A�
�����V�˵5�a#ص:�x����ا��B't�4CY�Cn>�����3۷�g�=CcE���|�5�j��lyJvm1#����s%���*5��Z���z�r��w��s��m3�kb�SlT�yKV�甇:j��r���1�:��.	���<]1�qPtQ�X��p���c�ǥ�����Q�rS�UӬ�B�9j�����EЉ��b/�1<�W`�2�{)�*�$��d�5����5}�WD����Ƙe�
����������mh�z���ύ����P�f��ʄ�\4�ё�e���e���'����և��C\�1ו��"�Hgȳ���z�~�6IO~��o�a��L���EMF$\4��ҍEy����Θ��5'e
+��p�H�w,ʌ��<�N��᠊��^G�}�u)������!�+��E��k�a���Y����G �0��(�e��3��<2�u��
g��aB~�g�M����q<Qt���0�T�z��g{�N��V�X6����3떵 d\����(OL��{ ���PE�wwb��湫�x���N�*Q� �5� F�7���H�B���U��32βc1Ѷ7َ��7Bg���Y �_Ү�$#���e4H�`�=[?��a^.M�_XEc�Y��;
3�%��}]�6/L���t�P����샧!%�yP�y�1���k�t��������KM+q�P����c#�2hM��Ҷ�E�H#t��cY���0�Xj�*]�~�t�4 _oղՊx�)�\�#e�(}Ƶ�X:Z�l�����4n��|nq�S \�s6l�Q?ߎ����a_2��?���TK�)�(��%c��Q�~��[��^Όt<�.��ƴ��$��=8����bةӈ�o���q�Sd]_�7߈n�3�Z�X�ZᎽx��q�����C-��߉V�}n�~��r�<�B�`�|ID�떽��w��
��m��� �'�y�~S�6�X*�����%��ض\Q|vR;t]����˒[o-n�����^����E.\�1��������Դ����BMU��!�NېN���Ey����a2'�*��m�����9B|v�H�p݄�e9_=c*�Ē�ŔJ��'Q8AJ��%+���YS�Å�1��ƈV�j[P�:X�rT����.�;�T�K=�X2�R�IڇH�Xǃģ Dm�K�T͘.�#��K���*}�d�"=t�j��~f�ib���9�������e���K�Y8���^l��������������&����w͹-W�=���r�b��9�Yd{ v��8�ʴ���	�]��y�ǐ$�)zF�`�9�UD������N�����$�M	ju�PLs?>��������&���Ü���n%�|�0Ͷ����Zq~�E����\�#��w�J�m��.M���(��6���o�?����Ra�Ɛf�.pV��n:T�4�um��i��Kf��i G���������ʐ.�������&~��aeQ�[�|E�����{+�e*o��5��`�Li��T؁.�vx�w��0Hla���Z���������)&-;Z�"�4��
��m���Ez���O����#�&��L�_��s�: u�W2�Y^����.G3�����؝8�,����9"s52=|צ�pv02�ҫ��%[wW�u}�<|P�qc�l&���3��Ԍ�0e�B.�M����tɴ���£^h�k����&#�a��9�~��lһB��5�p��F�D�0:���y�ׄ�%��OZ�܃`�㨝Ӵ��v9$�Φ�x�;Ȱ�ӫ7>Z�߿w��,��9z*�.��M]�FѪ��P��0^���4R�`���Q��G7�T��s�r�kg���:(z��BSƱ�=��@`P��5Y�g�����`\��Fwl�6"�ޣ�`���T+CJ�����lL�N���Nݼ�7m�^)wi�Z�Rww��]�b�8G2�b�K)�*��w٘�na�/�����K��8��8��a]���%��ُ�>n�|���=E���i\
b���
Sq��?��������8Ɵ4];4��j�*V����nΪ��Q�,�ʄ����կZ@�+hFόrMq4Ƕ<�`���H�$7ϼ>d�8��~z��I�`-ZQ��X��Aw�Fqzk��+׃�#��eD�x?�?�!�/�G��t��
�7�7�f�{�eUA�K����]�$/�1����EY�݆-�eJ�.���1P��.��������4����\ڗ;v�X#t��3ɸ�'l%��U;�:q"Ý�u�/<����>T�+�y9�$x�j�&����{�h�Y��{��U�梳��Y�o�0�k��V��Χ����x&-��i"��)�bФ�i<S��������+S�J��K[-+�d��^�� ��6�� ���3�gZ�T��+��I�0�vZ	�莉�k7τ0[���?�T��+��mX����?�1��ɀ������Aaq��W�'�B�JX�$��3u����"�/���S�ꮁ5-�*]J��}z��4e��&]k���؏Y����Kx.�o#z���u�:���`�S�o��T��V�S%���P)P�o��>3�o��5���\&RW<Kl�S̉���B��H�$F��!����ÏL}!��h���ې�����k�[���ܸ++-�&��JIL��x�1±-��@c
��V�8�)_D%�����mo�e
cHq�E���v���7Ulb�Q�#�UN��1�I�;C:p�F�F\�����=�R������������K�{��Z���s[�~�����=ᔝT0��2��h`r�,例V�!*�>C�Wl��/�k]9�Q�a�N���H���!߼b��u^��aԆ�j~_`IA+��%�OG$�̇��xP"r�b�aېbct����b���}u��*IO�q�/p��N�yD��]PS)�!�r�]1=�	����t�CM��M��"Z�,U4*݇l���'�R����?d�NX�u��ȓ�a�HPn�V#}:P��|���TԎC��w|foB���������H_w�v�((�WA��L*6��.h+m眿����T�	Ro>��C�����M�m����g�S:(8���.��1Ac^�'G�h@����}��"�v�������E���Kj�"��P�RC�(��OI�0��~�9& �!aV���d��ΧT�
]XQ��ap�{�>)2�|�8{��߿�.����%��Cf*q�t�~V<7���
��}���:s�Qʣ����}�
��َ���y��o(rȺ�hp�gv��Hw��
��O�`�)"M�yeP[���!�
���0�h�bb�!ں��E3
 e̶+/��EqhY�sF���Q�
3-<$�go܊�� � �/�i��ӵ�$�m���ϰj�b���,��97��c�͚*F&Rc��+m�i���vEE�~>G��Q�����߳�c�Ջ���ܞ�Z�9ύޟ�\���Y���g1rW��Ey�)������Q��C� ll����:{#���^�!�����������g~.j���$�b!�p�p�۟�4��s:9��X	\������P2�3�/-�q�J�g/��If�`6K<f���u{�{�DS8,��(Dy-�9ܩc3������l��A�d��)'@�Ό�y��0d��킂U�2b��~���Qd���-��Դ�g X���&G2�M��Z��׶fd�`	�Fm�OO��4�3�g:�V��>I���+���ؿ��ʘ����*C��q2�����(��k�6�N_��0�!Ҍ��o�Cl�/�=�vLEU@J+�0�fK䔅���/ײ!P[<@�8.����BU��Bd��h�"_����`H���S�)~���)6����,c���#a]L�{����%�d��Y84PE��ǈbD�6�V�
����A����N�YxF�ka	8��(�P�����5�k�t�9�o���82����J���
�G��J[]5�޴}����+-�#l����,�jc��~[������6�Wl�.�͘2��BY%h���X�T2<Lآ�q��J��Nb�i�x3Z�QsИ6��|#������W��+f��k�jQ��]HE��ߚE�EQ�|���x�������W��~G
U����1��N�*%�<sg��&gO���+A;b�KuK�T�5�/\��Qo���Ҽ�kkgۉ8�0�cL�~:?��TzU�����׌EK�䓐����k�Y�Y���U��:+ƩL[Y�f��~��-���&�
� ��x�yJ��+�1#o^�c�w"������/�ׯx�=�؊M�L�u��5q�)g/`<�[�?���k�q`^H��t�5��R��!��)�gX ���-��JSD�������.GS1Vcp�ךl�`'\�Y�G���'�͈��z���@�\FWq���w||��CJ���R�$�_W=+��|�����qa|���o��}㮹V%�ڜ:p4��o�^T)��*co=I�_Q@Ѩ�4<����ϟ/q�0~�&آtD�h���_���{�S� �=�7�nnoum���aH��Xs@p�X&����+!��Cb�a���:*r�\���pMk��Itl���nc���10�2�o�O���ˈF7��TI"�=_2��Z\�{�g�P[0�i&��cv'����/�p
[�������t�qdT�_b���̰�ƠS�=���f`��]`���Ѷ��i��:o�r�g�o[^���u]W�j$Q�W�au�``��o�;3��(<��0f���Dj��SG�z�����X�>7&�(6?Z6�{�ZҎ/����2���F���#����Q+�6>Q���L�`n��rC���v�QTI>��e��}�x腧y�Cd��
�'�o�Se���۷S���=z�G"g׏��)AHѼ?�F�b��0�P�K����u�A��<U�����*>�W����� �-e��s��l�5�c�7Ñ�"zrKY���(���4����8	�ܤczU_�B��6��aD��3�/_ޤ�h�tQX{g�؝bf��q�:�IB*�G��YY5Ez��O�Cꞇ2o�tzǮ#�5on�e����r�fe��;�q�nG�85Vp��{5
l��ܥ5�jᳲO��9��}	���q�>vҢX������G;�F�=�iHj吴��j����������U��hP*6����z���v\��fm��+R��v��g�]gw�,TO� �'[�YP >�����1	oT�e��Y{l�������XI������|<*��l>�);R2V�y�JGZ�K���3�Iv5r(N���j�
�ot�*)���ذPN��DD�p$��pz��������Yx���UX\�-H��	��r�Z�I���i]q�Qx{�bG��I�:#V�ki[l��DpU��t[:~������Sg���ٙfHf1`O��X�7p�9���1Q��5�������=��a?�r�^�|��}���V�z�kA8�;>踺[_�c�e�Z�FWw�He�=��]-�1B��y\�?��V?,���Ԩ(ΖN�C���������g38pga9��[�+N�.��>�ښ�N�C$`�P��	Y#
{/�#�fM�n-�����Z^�F}�L�:��l�R��Y(��U�4��D6����'4���4���oCꉄV:g��1Lc�ʐ:��C8�����p^���öpH_�jm��VT�����}���\�W���DO�,�͛}<\OD��q.���N��Q�{&"��^iڭ�57����|��)9���w���&�G~	��(a�ۜ�m�⢖7� ���>[U��r&����S$���/�Q��r��"t�)����÷��׿���m��c�P����!՘�o��IU��Un+��0z��W��ḏaGD��te��Ց���<���U�o�A��6�:� 9s�6�"���^�I�B��j��v*�KF��|�t��Ǐ��o%����,�d=ԨlM��=j���a�!iV���lY$'���q��3攺�A��U���3�����X��y��[e���[ɴ}. t�a��yP�7�g�)W8e����1佖�6͸�,t����C�_��m�gTy�|���=�`�Rk�cw�P�c[�%|�\9]g3m�i�vMD���lH�hc*K{���� �a�`�ݾ7���jn��vW5}�qhD/¿�0��.r�u��i��}QD�N/��m[�W�q8L��{��`Q-���f{����5"���ϑ�y�����P����hq$���.vo�pDц�| ��~���x��G\_T';�0A�M�*�}=�%y.�X^(�oF�0��_E���A�O��x���өR�V�^�.��m]a�at�~�	�l*�#g����<(�h�Z�H��@cxNV�U���u�G�A�e8.,�uP���%��yxV����Z��C;D���{�&�d�{�&��=�m���~'%�7��G��Zo��81f.���
��W��bW2���X���";6����ߢL��NB��7�����������3i3ћ����i�k�fs-�Z'�:�m�:Z��Z����K48j�B����N#x��uknq6���ڐ"�Ҍ�*���߷α:�ׯ|�]��F���kx�*5��nE�f:0���}�_ѕU˿��/�=�h�T񬓢�I"kfX���x)x~+��z��rPy�+���m��������2�q�cV��� �RD�@4���!|���aR:����´(��d���a��)���9�'��p��B��u1�����:iL��^���m��Mό.�lP�^�[
��4���V�R
����!��`�J-��B@:�7T�w��a����Q� �?F-�e���>|H��g�ɑ�SJc���,nr�f_����u�D�x�r���xv��˶�,�}��)X���5S"�� �wq�`�#��R�pQ������	����h�8>�g���|�=�B!�a��"/��tvq��YHњц�@µ�rڬ@d]�L�����)���gB�i�?��x(�*��Z��%Y\��fc�L���|��5��2W!�g�3�{���s��&Ӽ�P�z,�-�-�\`��=;�\��-;��g����&o���R�^�{�7���,����$��:̗��������t���E��\��4�ƐZ?󠢏�ۃ6�cx����Z�:��^�9�ɒc{)图�$���X�m&b6�Sd�(�5�/��- ���n#FZx��xy �:&�=�ENN�S8��tqAo���#��"�
je{υ��"���3�)IG�İ�kO�(�F4��u¸X��a;4]�$�Vi!+��<Q(�{詛@ne	'�n�)�dO���׬��|}:�dI�&�����IǊ� ��!b�2܃��I�YP�0�œD�Q��sG���xO�f���&����k�����dG��XDߊ���?���B������m�c�5���P�J=>�>���uMO��vԅ $���9`p7S���p��?������������	��)���e��(�m�ÞY8/���\ �h���C%��p&�\�fH���0j��$�n�c����U!(�����>K�"��4w�ǳ@JO��2���ߔ����n����������!��$d�P���Rw1b{�ϝR�Xh=���6*��ۛ>S!�$C�kϼ��
���i��|���Z8��d���N��O�x ��M�`��zj/\#R
�Vc���H�MC��t3ZOY�;>��_��9(}QU��ӛ����}�Q%"RPn���6j�W�� C��3�Ut6%@����%���ME�����L}nr5_4DcFw��(FFԩP�!�c�z:q��t̌w�6����혃��x/��~�X>n߱��"��1t���fd롥b�eb��F���6�*���áS]gdD��������%�����!�Nx�h�`�����ֻ�Ю��N��b�TD���]���y;�CD���}C gRz��PCFo��_�P�:T� 3�,��p ���g�PO��w<[���f<�ƠQa�H��p��9U���Y�OR��5�p�`��U{2^�"�_qJ�;�z���gOT)F��N�QD�8���=v���j�3�NȦ?���:�)�[����{���������j����ٶ0���p���!�� C���
1i�3�6G�$N)�ߥ(�(/<��0^���V���|�h8H5����,��ssӦ0����c<=�ʢ��N��/�`z.�3w��7Ґ>�τP�p�Y�7{����3��ɰ��{C�%��?��]��O��s.�=j@*�G��}��k����Qtj=�S0�Lw�(��q�MP���n����t�>c��`�ņCH�������͌��'�_��.@�� B&�M�{�R�IŦ0 7��z�����.OrJO�.ra�b$��$�����P'cZ��B.���>k
A���)�`��6�
���=�o$<h��$�{M��Ɨ`���b�zZ �jd]�G��g8x_��(�E�Q���R��#����e��nʳm��[�<��Gz�>���X�s�Q=��~_2����U�M
��+���H�F�=0 ���E�ޭ�Ě�4��%�َ�[�] �����~U����!�?����������ar�Z�H�xE_�g�ϵ��bŖ��ag�
��T�}�C���kx��������U�=�|�F*3�2^�,%�06Gͮ�!��K��Lq�,�=9��z؂O$�u����gUBe1�MnVu�uX�H�P@��E<'�/��a3�4D�p�f�7��gB���o �X=�R�������|ԍuk.7u`���#�9�"�nN)d8Jt#���|��))Y04���}�r��ī��X�(�B6�g�5���F������K�Q���6r0ñH������s��1�A�Ն/;^�O�&��8X煎紭/���11�m�� @D�1|n�����[��h�x|�s��
a�M�)�����SMad=��E����͈����hT�����a�ʎ8\.���b�I���)&�iL�����PѾ�ʺVA��{|s'�_��?�|X�@��!��[�/��+!�����a&-�
��Ws�[H��7���6��� ��!�hL���^wJ�����D� m���|�L�X�*X��6$��`QiE\��UԆ��X�*
V�؋3i��j�F=>�	�G����3##zkB�oxﮈ��H�_�c�*⻟�E*��Pf�o����{g�v�j�)���`'�:�.���ھO3)p�Q�L�4��Tz��gu��JM|Y�ԶQ�a�.�O�b�q/�쑽<GV25{`I
U]c���m���O�i��r'N2��c� Gnx_�ge �n;�̈�����눭�6ď�~��&�`r��B�i3��x�����)���HV��34�b���*��?�J����Y���?�n�n��Jg�[�W���E�ׂE���cvΠ�٦;�AsZ��0��gwR��t�̕�m��5#�H�\�(���bR��B��u���J�la�r�ºG}��W���|����«)�X4jw֑��|���!��;y�^�4�
O���:�p�^��7;��}KqW�iL��zᪧ����E°�]�`�zHgR��KVxp[u���,��%��.�zH{]��ȜE��e;1�VMTI��w��d�`a�6X�Z&��t��4�Yh�h��� �0�`��^�����oj��� k�rVЇڈq��E:x��>1��QM�F]���,Mfõn�Gv̽�r�d���`uw,�R��{�VZ�,�p�օ�3J,f�ڨ᜻�
�	8a3�!)�7��Ե\��5���L��=��+h˸�,)��$#�3�N!�����`���H�� ya!�m^��s�0/^�fʰ�jo�F.��/1U��mqyR�S|m���~�M4��]�د���8;�2�XG���eh(��k�W�Tȋ��A��>6�E)}Ua]��I�!-���.,#�N!.UϏ>#b{�*��w���Pa�ޫ���]w������$��W
�6c��ڰ����0l��M�H�������R��(�C×�T�b�&�:uyW8����*��i�T�Pp6ǠU�~��`&j�IX䋠	��{4��c��:Q|VpJ���W����HX#�U�Tald�Z�F%eb�H��<H�Cq�:���u��`���J�7��FS5�S���Aܠ��N��=�*o�{���r\��p0�i�C��#��ߦRQN�Tm>�"* �׺T�ʮk,C���:��PÜe���C�L�N�H���g�hI���t=�0�3��̈g#��6���i?�yҨ��)���g��<'��j[뢬?���e׿�}�\b���tT��v���1R�<0G���>�g�lT���
�A�_Ԥ�@��ʨ�^���p�y^����R!I��gD9��CE��D�I��Ln��Z;�" ���$���t�(�d��d1�*�}�=��:{�����,���֮��]��j��C\	�,B���o"/
�,(L��Z��56x;���� ��M��DF���r���F��Hv���Dqx�`�®������ ��r5n���SD����{n��=�Q��\�%��)�*�k�Z��ǁ����p�E.,�ݾGwu�+O��L� �z���cD��}��u��D�^ p�|
?l��Q�3����K�1��R�t�1�V���@E-*Z'�SV�mTa8�@���"���g���]*,٨�����UZ����Ru^�	�&�����O[��*�� Қ��Y��`A�Y��M0~�k>�_�b&���ohL��<v;q����ғ��d��ض��-�tr|A�E]>nZG�/g�Ԙd��),���?_G���h���eY�)n �|W��-��Ϡ4�勶�V0 ?��$�>hD8���;��Z�6�v�J����g�/Yg���g�H�q��;��_��C��������P��⁓b����a�Ԝ�q8̫�	��F� :��Z3ӰIe*P�^�Q���Φ��&I�o@[��Rj/���̒J�^�%���#�a$�h���+5�,���h�y��|��C�3��_����P�Gѵ��9���8�������u�6Ɲ��48��P�����ٹ�PS%\�s	���Y4���>�c��"4�|,����u���������� b,���B'�&'����黽����Yi��9�f uI�S�(���U4�l]�l��+��}��K2=�o���Ad1Ǘ�h��2ژ���e��0�s��>><&3��t<!�~�|e�QPTÀ[X]�`��ʲ�\�cD���,�7e��~w{.��i x�b��ߍw+���,�y�R��ciM������̕x��d
1	W\�8�Jb-R��~�i��ڧnWuz�����~�S��\IxD+�V�j�u���r�ݏ�$�wHո��,}�gʴ��0���ƮꝢ���'H��*�T6���3	4��6��ZuIE��٢�\�7�V�T��^s�$
%�y�eW��W.�"����i�5���#�7G#��Wb�h���1��܍d�h�Lvn����Ү�Y��.�l]��ਣ��g6uQ�`�[�Y�I�84B�9A��2[	����٦���#5Ӥ*&��2/�qn���:�X\�m�'�5��K@\h�(�ptF]O�4�\��(���_5��f5h�@v%)�������A��0���0˨V�)N�>pj�uW��1�Rd��y�J���}m@kP�}��;ӟ��}U��C��DJ�y@���Q#-*��e/��l�6~@N]��!.l�N-$�i�8,��]·�b���U������,"�{Epm~[��o����V�*ks>I���������D��$��е
�8����=�p,�zϵ(��)��+�ު1d1�tG�^7b�y��^��%�ܥ�9ش0v�S���*k��Y=][Ȝ鹐�y�H
�9���Qs�p_�U�R?E�?O2�����DǶ�Q���.C��,��J�M��3/�ERJ��z�^;�fUosys�,g��Eσ�7m��i�^w�`]�Ί��ϙL���9��nG�A��Q�c�%�*��ɧ�Lxl_�b����瀱͍��j&���n!o�uP�h�g���ʛ-Pfٌ��s�H�>F9eቒwt`7��� V�̵�w��ۛ�9..�lN��^Ic��7>)�sU�k�!�!����K����O��ّ~PA�?�"��*�ϣa+�Ur��4�	�q0gW�fzd)����h#��T�_��I-02�����fɂ1B��o-}��V��@9���"6�1?4
+��|�I���)������H5��H�A��掂��\�B��k���~�(�?�{�0ɪ��VM����:��E��	�LeKnzٗ��7�؈-_r�4��Af�ScHo5G�k~z��L�}#EEo3���R�� �q*��R�HэtG��!Z7a�M�����X���	dj	�s\��_�hS�d�Ds�v_w�SR�(!W1C|���D�=�>�lx�:B��n�eD�Z���O;�6�\��ρӆC3�ϭ��#���cm�Ta�l�#�V�!����-�S�g)�=%����ۚQ��>2O��=�%���,^F�x�f���nD��0
���d�D=�w��,��(�jR�i�	W#�
�,u�c��C#�}���\D^G!�F��i��h8'a�-�o����Z��{�.6���/�{�ƽ��U
A^����z�ￓ��$B���=7�j����j��L]m���Z��{�#�������헿sV�����u�u� 1����MwȔ�r`�8O���s���:~���)R�w�mh���`uޝ�}Y,hR�/�q�hO<��y��p=q��ϟ�7:M��^�1���S�(�#\c��� �w�4�5�N
�i>�$��y�gOu��ta}��f�13�H��b4��3�MЦّ�j���r`��4|%��q-��5FQ�2B�՝�
�����w��B����.��֢C�*��9}fPQ���L�o2Ev!���`O���^���x�蹡F�!c�#ڻ.�]na��N��h<>����N�t�1B/�(H.�:3�\T:���	aͭ@gչ�s��26�r%3jK��Φ�+��?�-A�g���7Q\�,���ΐ���	��!�Ñ�K2�)�4�rVG���<{�~c�DP+���O�p\�C+^K��T94ǎ���`����5��m㌯oRdG����>��{a�cα�sJ�L���Do��K[�9;���h:O���Qɸ����V�Y><�I��Na���z?O7�B���x[��U㑓_���ϙm�P�މ���1�]U��?�ӡ�cB��D��I�b(��=�����?�9.�9Ee<Z�wWb1xQ[������*X)�xb�|��f��8)�����(��l�҅�>}��&t�������$Ir$�A���!�X�{'w��E9�[��ú�IU� /�T�ܳ�g	�%P���UI"�����T;u�M^7ͧT͝��S�v6�!
W$ ��K^'�[���0��x!�ol�m�F�-����ٺ伆6�T�h���n��{WY"���Y���L��Ч]WI�	�Ĵ��S��6{�Z�z�5]��?R�n5�oGW[�f�m��e��j���?D�XW7;�m��|:s��D�f)����0��I��Y�� �����Q���t���o�U$Y�A��r�����\`����T"jU�=���uLA��ٜ�Z�StR1X���+�-V�u�����7\J�$�s�PO_��I��sv�]L����ٙ|m�)�{��%ϗk2)<R��."�[���ok�E��@�~���l��K	p���K�K(����D��Y�P���kl(�����o~0J�oA�R��Z����+I���ԓuO]�Xx'\f��;꽡�o��q9�,�m*9�I��ä����A'ԒX�1t�旬�"�?���	�����c��`s�m�5��I����Nt�%7<�ȸcp�z�Ъfr4v��tM�q"�1^W�X�0����gz�0I❂]����C�77���N^QRR������4��U������|6R�aa���Aa>��߼fSg�;��M9k�����\R�d��0������?q�(�v'�O-[�"��Ւh�x�!�a��`@�"�}��hd���}�s�t��n�����R��93H`�P����.��#3�s����r��b00ëzJp��Y�r��둄xIZ%�YT��Y�/��+qY
�fY������O(\nY<%��P���v)��|�5��E���^#kEV����[�A8�v������г\�{C ���3��������?����� �@ښ,����Q���)C��:�\9��� ����E�����B��|;��I�q@[��h��X*��;�׊�jh���)c?wÛ�T���p k=?Q��u�2�C
���]��\g�R���d4��ލ+�d�Y��
}��>Őz�F�)B�Hp���?K���/�������5����s_�h,�d�L�{{]������6#�n�0��y��=�χ�ڥk���R'>N�N�Y:�}��C<��3�Ň*(��Q�$�q;�[)���`@��H��E��N���������suX�B7����z�:-M/4z�f���NCe���.��3�Iy����{��Vٛ,��0J����"=���̒):����f�{�N�m�p4���Մ�~��0~m���ZC,-��Ž?q�>�φn�kf���,J�^�q�=L�[ēu���u� ν<�,;SeJt1�������:]���bzѸ�y` Tx')w��c�㐊��*�vez˼�i��#�O�>l�Ǯ��j8��r��38()���4~_;��>�"���{OK�[}��W9*�Qn�W?���!�U��eҳjH	{dW<O�f�1�B�z-~��Zu���������jA�[2����6{���6zv��6I-��4���������Anu��� ,q:��k�/d��dwFy�#�k�\JInT�75o�	���oj��
�Qr��f��d�[b��;��m	^6qڬnP���7d5fI����h���UO�.ac�xNf���@\E�)g�)yt/O�`�ωa�=�9{�aC�σ`bkl��c� P�ȩ�l���Ǹ� �c-܎�������j�ۍ��a�k�#N�^��{:�)8J�g�wg�$VAq�Bț��5�T�\P�c� ,��5:Jڸ"��:���3iY�JL�RE@x��u���M��T8dƳ����΍{X�JG1d"�� �m����R� ��盰�>�Hg\G���*��\\P�
1��!�l��Af���|�70]̕����p�萯Z��L��[kS�+Q¡�����g��A��p6[_���M�d*��F%h�_��z������:.�1y��t5����$��T�ә�#�7]Ҙ8I�@�gJJU%��%��u7�Et��l�e��r���@i�����p,un}Vv�n�/wH]�Ō����xA
]ɽ'���
<V8dC��OĿ���L�:�������j�_ؤQ*k��~���4�{�U�dd/k�Âl��h�? ��e��]��ͤ�P����?�6���w�^�ǟ����g?����a�R�+�l'�܀upD��>�;�#�|I�m��z�v���Ի$�� ��4����'*�y4q�T���	�����9�aiH6a�V'u��]��PL��B���M�q�΍��(����*8g�nd�����q�=}/���B&�2ؗww8(���[�^�(���~[޽}{�_��1����K��J�ВpʲL����1#��*h��bY����e�_	������������l�v��O�/sf��=}@_���m�q�s�Ѡ~J_��I��J^��^�
4�`[��y�n{2��A-r;��QP?|A������(�_�.͜�"����]RJ���vWӣlU���v�}Ԓ�A	��0џ�����8	�]��8���|-�E�L���۲P�|��>����pk��.���)H��9�k����b��@�z>���c�x��m�F�/3ue"G
��W�)�k9�h2��f�/���!3��6��	~��L� ߌA��d�YpG�� �Z][���/MSeT���2m	����7�5�eU}ӹ�s�Ʉ�F����ymtU���&�M�R�E��bu-��GPe��9-��!L뗎���-���a a�p���ļĵƇ��ۯ����q;�?]��v;�/	����y����4��8W�y�
�=�N��e��0�I㩋��T^�����y�#m��R�if��'T��3�~6��7ֵAo!VڄX�(B5~f	`���;��a��A��&d���plb���i���ٜ?��+/�^t��qZ����1S���X��c��[]@���Sm�7�^R�E�#�#5XvM���P�l�x��t"W�2m�ʷ��I}�b����~4&Λ��28BY�G)����.���36�2�'�k��,qLS���	�c�����Sl����{֤�����`Q�ȅ0��@�>K�Ž��%~Qg���y�sjW�g�n ��NB<X�$�۷�$*���g5A�����E�ƀ�q��3I��	�X��vx�"�6�˵wD�m�
��a��n�� �S�O��P�o��8�'�Lw)�X� �yY�{��p��l|Ο��T��kHEU�0fՁ���G?�0]"�;�����[�1
�O�@+Z���&\p���p{h���_�r̬��cm�O���뷱�k��O���	o0�1��x�I��@��:�q$�))3(g�.���%�e+ZGV�'Zk4�P�X�ռLE��L�d�.�L��}��[[j�MZ��7�z�8��<�k����:]?�؛����=�\�:h�� �-Ⴌ�c����X=o���
�n\8�� v�h�Z�z�I��:����9A�߭-Р��PUC6��]뫔�����@9~���9�-=*��;6--��~v�=>�PY�&	��B����c�x����F" �-Q��^��*���m�g�����O>~�����-ZKfgTII>1;�Q~v@>�q-�����>�#��:y~��������WƈL�q	x?
��#�H�O�)+.R7<���?�esp�S�Z�;�{��� �P��o�>Ӓ�ن��6��X��sR[��#��/�0C�x���e༭�M�o晘�l���ky����œ���~?;��^	#���%���N��D:��M�����#���$?1s��j����YiPḱ��A�����T�K��Ms�r� ʇweN ��y�bë��\�9�̝�6d)� ���9�����a��i�P��_��Jf��u�AT�#-K\�Էg�'��_C�� ~8شm|c~��?�{�X�,Ec�Ȼ��Fn��02��/�C��z!�����pc�Z�2���P1�-U�ą��ZW3y����ohM�Jpo�^�=>�ԦD�����!�?O��4q�$iG�P�E�	�E>P�~�����s�[ЄGE�\�e !�zRs�9yӥT�	H��B~̊M_�ږ�s��Z��� �i����$|We}��)s
gџ�/��*l�I�G��I(�3�_�(��=�`�'��蹾�ᱝ0�\*��u�XK�g�ݲ'��yk1����Wk�<:Fj�uK�Q+F��;L�p���d{����D)���C,��L��L�]���*��4��,��rM�RN�5���M��t���Ձ�<Ek��c�U`�S.n,�����P<�m/�K<�'I��C����{�bv ���(�C��Ƶs�i��M'4��;f��C�&kɿ�V]%�;w���r�y���!��/I/2�%(T*�=gtp!5}�y��O�'{ꬮ7"/���� �=n�.��)�(�E�����Fz=�#�inX��]q��>is�ڒ]p�I>���O��x �r�j�k�qU�n�8���Vý^����m�A,���ג��7���qh ��,^�ߺ�h���Xy�x�dR�a&�
�H�@�!a��j=�J{rS��K��2�:9Q5��S�Ow���Ԁ�eD8V��V{����f�-�؋��R�����������ޔ���c�Y��V���	�褍�T����
&7E��������;��2�Ð�]����/ ���@Q�6�r�J�^��Z4�2�y�ve�ؘ�d6�
��A�ƭ��+5=�n@n���79Yn��wO[J@��*J�ꉠ-e����mZ,+xIs?�s���'҄>I����G͆[k��4��������Jn�)�2�Y'�
gi��j�A�����k..,mw������Pm�ς9J eR<<���L]�eS�V	���s�69���I�E0���2�Ku}\����j��^�a`++Jq�����<�q�;H��A�b���-�:��-5�z�,��G�E�	��O���t�4֘���F&���6&�SP�EC���	����&���w?H�:mu�C� �Ȧ��c���������\8}�`ڐ���}.��q^�H�k��i/�
��k�|+_�HM�#�jM��8%���]��&�n�s�T����;Y��#h��#��߸!�6��v��i9�X���@let���^�r:�hM��=��c�����H����k)7>�.qPB!�>�bH��2^������f@#d'ZQQ6�e��b���f��/ZQ�f��G������97+~���c,�m�&��uv�F�ۙ���	Q~�Í�k�m���=�q;+�IGԎ�4�벌K|:��5�؇}l	y�M�8ȥ�K��A�Y���i�0����W���l/��C�S�-�md�� �%T���Nk��Q6���I$aW}�bS�`W������'�*�a�����~�I8|�����`�� �2M���Ym��A��������Y�1���Ӷ�y�$Tu~�ֻiG��}Z�CDVp�1v:��fhki��[�U�K��s�G��N�HW�|�0����O�BU�����O(��W��γ�uq�?4�7������I�.?��7�[m@X���3F`[2��"/���F#+l/����^��X�`*+�,�??*�np�Ť�z�n��kaY��v���xp�G�NȠ����~T.!���߳� ���kd̕����=��wmwu��#����nz\��s�ln\e��F�3?]<G��;a���Γ;��aK�к����(��(+���~f��,�k��i����H��A�E�Ym�Sq��,l�s�=�j�5����F���;��r��능&�p��t�'�f`�%vj"��D/�vo�Х�f>~)�F�{��%�SL:��nR�*���qf_�8\��E�Y��=	�x�x/5�j���(G�3FTdUS��*� O;���2�4ͦ����y��iҵ&n\����}�#��Dw$U�o����[2U�΢�d�x��`�1u+ii:,���i��U��Wo4N���4ټ��0$�6[N�i��z�`V���S��:9��Q����ʸ��$*_4�*�}A�Y��;���k�_��49ۯ��L�ভ|_��ή5��kd�|�u�?A�]\f4��msW���EVˠ]�Lq?��ӟ�J
LB�疜ݧ����7_�ow������n`\R���4~��"���*�����`����l�%�aw��y�eߣ��ꊬ�9A��a�?�����?d��2��b%��*�5յ��<�f)�Ag�I���:�~We�@R����N<�����O�5���>��[mq��e�� Z:�G�R_l��y�uf[6��W��44�N�|��Sb��uQ���9�j�x��o�f�C$Q��Z�E���(b�� ~p0Y�[-�R5��/Q#j\*���s�-�^��֌��GR{�MSW�}$�j��KJSQ*ZSR��2���$�0��y�⦫�Z�j��۳d�iɑ>r�v�ʍ�9�^�\pm��%�������m�ݝ�}�FC�y8$���7㘣��X8�?}�����`j"2�f�n$q����h`DG�0 �j�A��t$���Z܍v����|�������̼.�s��g �۲��{�j�B����|�X��Jm0��P�<�v\��;~u� 辣3�w�;�
U��y��`XI(��{(�b��R��cs��>���. c}AiE��B��3��Է��o��6>$��&Rd7eε�[ۿR����CN�=���=lCMYF\���K��A����N�T�9�-w�F@�����̮y���Ἵ��{�Za�"ۚU6���2�;�6����a�n������߾}c������BIJNu�0='��K%��^ڈ����4�c\f�Z�!~T��t6�������]O��1��Q7�7��b}b����m�zvE�S��h/���:�h���5fޖ�+m3�N୳RaQziZ��l�J�Gg<aU�u��3�M�E��ˠ�!�z���q���3�4���b*Ь��>�=����h�f��	S�������tkv�4Վ�(F뢌��c���V��!I�v�|��+d���C�zۀ(�p��
��Y�(��:�V���[Eɹ�l��۷R:s<s]�o�㡰F���W���*N~l����O���ʟ��O�@L>���ˏ���l`�`A��o��n����?�g�����EϋD��]a����
Z�L;��M��s�(�C�R��Sh�V)0���(~���/ߔ?���D:���h����{���(���ߔ���o��sP���kQ)l�C	��dӫ�ϛ�o�]���c���M���
t���t�sn-'�gu=f�h���u�x�	��nI��G�fF
g���7���s�d�!�Q���q����^ӂ}�ئ3I�!U@y��HH�l��|H;f�e�ػ�p�)x��T)U��f�]@h��?����`f�5�u.��gn�`�~�Sͦ���6�f�K\���^G�Pߑ�n�r-�,��i4��B�\j>A˙�]�p����D�6�R�����z/6�r�o�u��/�>fsq�}8v�\U��gk�F�s���vS���-���1%q���G����g�PZ�j�ӣ�AI�.���'�v7��{�ga�94:�����W�%N�`#�����YSk��=�s�zr�Ũk_\��g����l1m���!���}�����AV��-�w���5Ij�5��&D�2�D�>�N~ס��D���.����u�542ͷ��~�кW���9i�~UU�
R������{@#�p�<Z'K1Z=�S���q`�wׄͰ� 	�@j,c��Or��A�o�r���>�U��N�k�h|����NA��"-3ᚵ8\�[<\�k����i��?�jw?;�/���Y�|D�w�Kٙ�g���.�<�	����hk	��K���Lɹ�.�e}.�Pv������w� qY��9��!b���۞2>q� *`Ƚ��?>q+dZ(OQR�=#�����L���) �0�V��>���H-�L��C6�b��4���&�<��M-�Gɉ������,n�.�AM�k~N�[�eс��AX��[����o2�w*��9��?�;RX����?O��	b)Ӕs����e'�� �3d��|H�I`��k�g�����-cň�뵏�������� &��3"�>��poI@�uz>��ú9�Hfc\/�R�?s�\FzﴢSdǲى[|/��Z��[F�dv�G���Ͻm�;����0ѣ�Yj��mu��� ���=DV��'�`L�5F�b~��!����a��57��-��c��WcGZ��v#n�ц���>�J�v����+G�5D�r>����~�>�l��2�y�}���}>��|r;��x������`'��n�����J�+?�"��[0:_2�8*���Q�I�-1�_7��N�E>
����U��&f�T�*53
��k�������7qs�*`�8:�Ӕ^1�@8�v��Yw�������n���6ʼ(1��GX�`<��#�"����<�v�>�7]�쬊R��l/�9��Tqke��o��&���dS֎Ĉ����V�C�*&^�cB~_�����<6'��c�,�f2����gÑ�#Mq "���k���ꈘ5��7x��u��5�����x�H����%?dJ#^�
�l��^��T�&����_�����{���u�f�tJ"��֩��{>s������X3�p<�ն���?���M��_����_��"$ _�~7L�R̲��K���Q5z�&0�}ϳ�W>Л�V<���Q��a+��ƚ%$����c�ˠi��������ʌ��	�/3Re1+�޼���� �G��ʹ����6̋��.v�;�j�hv�=���"�q.����T���a�� ��Lʌ4������96�S��c�� �Q�]ˏł�q�&�Y��TY�"�2	�*�
��(�U�Ԅ��h�5	�;�<uu6��v@�{��ԫb�H�?c>k�����z>�OH����x!���ݼ��ز�7������M��7ހ|2�<�>L�d8`�Iӳ�a[fp挾X gAE摺��^Uz�!j����l^)�z]��؃�����u��WuQ�E���2'T��\/b�h�Y�9x�j��k�]r�^�kr��Ư�{�/5��q���g�ӻ��U����@�x�9����C�P��.�>kC���ӭhrp1#@uJ\�@z�h�c��Fh�K��dУ��׻�\/��a�P�o���⢿��s��L�z1L?H�'��4{�*)��޶�x`6�F�Hؐ��鴉�����S#�d˒[W��[X�c�Cr�$\��D�Ϝ#���c�{��i�eP[�k�4�w��@I��9ի�X�v1�0�n G(�r���=2D�6�������V�ϑƠSMW��%57�i�m�dzd|fp)ׅ�u%'����R���uU��S#�:4T�D���*�#�3����8�H��UgF&Xg��������c�?���'H�x�N�!n���U<KOVY�o�W�a\4ۆe���U�].׫pOR|����b��\��p����{pqh�p�C {������!�G+�8�\�����	׽�I�}b䰔�������xH�+9�k�6d�������Ջ�YTC��ۆ�!��B�iRv�5Yj������E��aLڛ���p���1�{�� �8pE�s/m��5����vkN��������>�����q9�_�D6��&��N�P�1���d�HKwu�o�2\��qS���#x����x���!�`��"���Pv��WY�J��	׹����Ό3rUI���c/����T��@P�ˋ�P/��faA�`���j���m�� x�B�x�)�R`�y^�~��xKIƁt'�ؼ���y��k{Ǜ��CCg[�8ݖ�,������*�%���F*-S��%䶵�~�BƗ�)��yJ�Gݫ�cjZ�.�bUX��MNE��h7,hxh���_n�Sq��a=��h�l�"ή�yt�ٽ�(�u��b�&�b�K6��<�zцFӇ�R�����tֺ�ڧ�h�G�]]3�N���������}po�`���yr�EE��/_��τu�Aՙ���� 62pV%?��	%�xI{i�b_�ps��=m�X�`����=py�.�Dvf"�����6�����/����eоi&�4�\�'���Ɩy����e������3����	��5}߹��1N*�>6OGM�SJi0�ύ�0��`��� �<ƇbMS\�7=�O��9�0v+1�ikF��s�E��zŠ�Ec��=;�X��	-������ ?Ԓ���I�7�z�ʉ��q;<7��%�I姽��-E
�wY6b�b�yءf�
���`w���6˟�N�:Q��DQ'�BS�r~\�Ai�l�`��n�2�����x���(��7:�f��c����M�<�*����%��Q|�R�c����_���B}����דw�{A:3m��A|`@F�N�䇃n�>��1H�gF�r4�G/au_�Բ���/�jw �~�P�S3�5},�u�������׿��|���X��	��ٔ�t���HF�'.���ze2�%�(�/3R�[
߻�@����HnY5�2���C��A��l�ob܋���&S�Yr�Z��$YWnd�ܥnK��r�򔖳���]�%/ ��8���R'�}���Ɖ���tKzo��Β����	ߍ),~\<S&�Md�5��� ��]��<[l�^�L�,���Y�q�A�LA�,NLt�-�RD���'��(Oo�i=Yt�����y:�~��͔]Y4����"2�٢ȝU�x����&�p_.�Qt�dA�ZYW�/ǉ��H��\6�]�:����R� ΌG�����+!&�ڳSnT$@�>ꐆ��fN���]����3~��~��c�D��l$�:b�u���ڋ\0���P����$$�~�s����u�[�Ã�t��cjMe5��NN�U�'��C��	SL�'�\Ϣ�~�V:�Y���e�P�Np�1�L\�בW�`j_�����}�)?+�y]��O�Z^C��)X���{q��ÿ)������柚s�$�7Wүb����5���V�p� ������-M�����B	1��(iwj�Ĭx �E��P���Q�a��A�9�j1�Sjs������s_4������I����5�<r,��Vc�BΚ��$�u�$���f�;³��ÐT%c1x��y�h<ܱ逮7ԗ��Oo^��:>��Z,�C�J���6\[u�=E�Qؖ6�Ӗ�m�&�Il�:�s.�96�/�e|>l�!���,�}��=��0⼇��3$�n�]nJc�$�ӛi�F����VOs�^�+�s�R6�F|t�B؍;�2�D^�Ce����Lա�qNe�����s�9sPe���k��]	>�+ye����ӳ��!�;��1�.n�ik7=�C����G��x'���h/�)8�Ac����dp�*2য়.珧��Y�߶�N�)�,���;�bϵ:��χL�)D¹�#a!c�A�92{�m�������Gb��Uk�d��\�z��K�����(K6�;dl���."U|�� ��$����"� 	0wZG��q�x*���ޚ��Sȟ���� p���y,�bj���D�M5{�#d(ۄ?_j�M�
������8D�)�	��Z�uɓ�vΚ7���Oi������	�P`?Y�^M�F��c��90�[���w�@����.|d#[�.�IS�~Φ����!5��%q	�,'W��} �,)��w�����z���aga[�0�k�M��Q눙]!�bf��Vk�#o+K�x�l�V�����x���k	��-�D[B�>FDe4hoyg����j�1hw�����_
XL���&�r\{�In-�"�!T��"��0�v$#���31 ��m����Op>���uܮpT\L~q]�@�^s?[�1��V��+)iN�8\��9��q��Q��ىM��H�>��<"S��gs�j䶬o)PM ����T��h��oڈ��@�]i<�-/�	�t�����b6N�FT�i�F���b��XHn�8����M%nS���T�4k.S."��^�:PR�R��=�t�E*;�e�5�1��TWͲ۱F3�������('tP�c���&H���:gVϑ�����P����J�d�v'}G|h��چF�/(����U�6�����}��D�*1v9���s��T�5&��q�uu��~��q���k��#�3q�W~f�́���\�����
�@���8 �ɓ��hU�:�g�3Y.ѴقFW�y�)���:��U���d#x���eR��m�p�ʵt�#��ԔM�k��AC*�
�:�!�S~�W���y��_��^���M���+I����� �/�"�$*["^z��n e��gm��Ҿ��Ϧ�Ң~sQ�/�:�>��Y~�YR���^+��E��UcVervus�.��u~�⢴nm�_�lWo�^��|C��Fv���N"��̓���XMP�ix*ܭ��}�Lc�)d�4��F����=�>��"������^���Y��8��:U�n�[0=�̒&�"	|ɃA3,������UK��=�l\�9߫�N�5k>��}x��Wu����ὤn�����pΒ��}蚆� %��MV���Q�wQ.>QzM��J�MG� e*�?�ZQ������'N�����E	U�2J���k��6�~�M2�,Bَ���Ʃ��'���J|��Zs|{������ ۬ؖǪe-t�φ�����5�8C��c��E&Y�-�Oۑi�K����F�X�������3s|\B���]|��F��h eW�p�<��d��їA�������	��<�M�?�,2��{FrfX�F<귈�̕�^@�q��Y�mDy�:0<��C'p�|c���=[O��t��l��a׍�PY|@�E�2D��Q;���̞����ݾ�����	��ĸ��V���\<��DX�����WF���CbL"�� 8DP��
[��C-%e�]���/'
��cv�c�|�%�z�y̯�b�����1M�)a3D����7qt�yk���rY{�U�g��[�xz�p�,�}������Ɵ-L��F)1궲������Y4� {,{9�j&��[�E�.�Ӓ|H��}ec��V!S���ύ��/���Q���t@n4L�Fa�6�+���.��;}�x��ľ��J�!����'wy8:!۫R!���ʪ�=UC�Ӈmu�+֭�5U�v���� N�rH?7*�2v�-����s���H+ �m�ܴs3D�y�?J��WY�X�0�N)�!Ԓ9�o)@���!�4F�IBO��Q����r�����o���D������-6���P��`�\��͡�T���f��U>������-���)���A��'r��
28� ��d���b�c{Ƭ����
"C�kFF
ag�{e����� �U�$��츒括.��J�l�a��C��e%&���`s�T1��}_K�c�%���/�����q*�ݷq�m��9��������f���v�x�X��.�F��g�qO��q]^�E8�D�7lF����e�`0��5�7݉-A��Լ�O�a�T*��5��3�[麪�w�l��֚�ޯ�[p�B�O�&䚛ܒ}H�p����З����������@s';�g"k�Dۛ�nJ{g��3�8�G��KV��ңu�)��������z��?Ta�'�ط��s��6]K�qm�>g����oJ���oI�QY��T�r~���v�$�|ǡ��v�ÅGm>J�yN� �i�,I������Z:S �Lb�J�/�~Q[����8bY�+��tC]������g9�,yr"�5D�R{�I����0��:��ZzF��j��R�,�����4�U��}_;��=�Y��kEO"��)�mQ���)�{7D��)���N����]t�,����ce�j�F��>�=3@l�*�a^�ks�" K��n�Dè����e�7�!9�Kfz� g�/>��s[g�q�.��XJg5����R��qW%��vl�Z�x]�̓|����K�a�������Ɔ�xcS�$�|H�_r �<�-�gc���=V5*�	���!3	���Ȁc0�'�#����m+u-v�5G4՗�}�k>i$�=�~n�(����Cl,7|P��eɪ��oB�ON �ጴ	���9�t��������� ڈ=�-dp�7]/��������ù�1J#|��c�V��'��7��� �l�̅��}�	�߉��12�h߸3v��t�92Hi��('G50��Is�9����m�2#�gƵ����oLq]*(��Ye��}����e�9v`�G3�)�l����:��&G�QHƙ�*e���=%��K)���-t�03�13Ho��da��%����pM�?1x^�3p��(T���gW�4��M��5 RY�E�Bf��[?�X.���0��X�p��w��sZ#�����
���LєS���,�?Nὢ��ݕ�Bcj!�]]����c�'MM���5N�=;T>x�f��Te��5���,���I�в��&���o�q�s,�=�^jh�Z{%�U��^�jk�duT���h�L8���up���]M��o�z���YN��-�Q~"��.�f֐+�������H����G�0�>�I�0�g�h��72�*GDY�y$��{*��"�؜#��>���ByV�e���p�a����F�<熻���O��b��t��L��]L¨�Z� ��� ~�%<���g�Gb�����ӹڞ\�ªkӍ�,Kynbb�?�u��'���_~��	6��6N���Gl�e��2/y�[W`=
ЗسG��W�?�9��ӧ��#7^Ã55&�ƒ��%Y�ED���(��XC��gMU6C)]67|��<9~���&�����ǽgY�^�q�<��	�i�q�	�)�����~����L��mu�wǼ��*w%=�^�y�?T�g�+E~P�\^	��aa��D:S`�#S��Y_7�P�y��0g��HMs��oh��� ���;9���y#��6zd�����4�O�An���2Qn�kvν���n�".��C���u��"+M��gzT��/՟��8����݅�6&S�2s@#�(<Y���3�����(���(�n2Ŋ��F�X'YڇŔiJ6��(�z7%��P�萴|�k,�-���e��w�WQM�=s(�p��>��,��yROqY�Q���;�qb�`|nd-ԫ �x�����\Ж��Wx����ʴ���Y��0=�
*�ƴ�V�������Bة��/���$�hA@�P���z/)I�R}���U��q�R�Y�)j�4��Xi�q�|�%zW�lx�1���r���^��5Gfs3r�C�r,	{�o���`��[6��:����:�w;�� ��VV{�ά]<�:����k�t֧-�yg���X�3 �]�L��(P���-�]Gd]�$Ωr��J4��IB�!��L�yg4K(Y.k��6�m_��o/,�S���Wc��W-���������}��Mv�q�(�z*�co<��'9D�3�c7��I�����y����J�-�S᤬��JH�WLQڅ1���9q��YĻ�*�j�&r���^z�~]�7U#����9����6�3\�E��Ӊ�.<Hc����?������}Pq �Cٓ	��ϧoy�uх=�X�21by,���u�:S��_Z2fb1;�ߛ�o�LS�(�qݮ?�� �˝�Z;�suq�l����0�29�<5͆�b���%u��lv�3�w!J���{/�����1�Wxϯ�Y���L���h\��y��e)�!���HJ���|�
7m�'}o�2r��b3P��T�K:��g�Z���2 ���C���� ��Z]��0���1�Y=�(����a@�D�'Lr+���FQ@z�S�G}����kPX��G�����!�m�b�'�]m�l���)Ɖ�\nIퟎk�: �Y��'V���}�Oi頛��X�gP�f�N¡Y ��]0�2Ͳ��?,Ynn�tь��}����{宒�����%�{qR�B}��K*�������^�cnZ�eC���%���T�]�M���#0�lg�Z�vIA`��xo_~�e�0���N*N�Y��?�7bӂ���Oc`��J`�y̿K����~����'�IԀ-��t����:={.������17�`_�$�>��ǟ" >Kَx�n������k�Uy��?�xt�*���!9��
�	��4Js�F�Ǩ-U�������4��-��C�_Y�^I��c���!8�C��:�&_�<p;4������x���g鿺*�[���Ycd6�\�lH��ĩ�nq8���&��ϵR܍
�����yω:*[���!�c~,t%�[}��H�2��Q�0�b����Z�F�ߊqMm��LӞ�6��F�)c�ZR�Y�z���D��u�î�}��cbòwMѸsH�g�(nx��=}\NV��K^���u���8��r�#Tm�x�f�$u�era��n(x}� �)�P�FwU�'7��j���Np���^�{[�WK�d�����Z����W�aPf�&�gz�����im�1�`ab�<>�iDpD0@���ߗ�[��y���L�#������� �,L<�{*���Ȫ�EF�k��As�������]%�_�?Y�ib4қo���Ȧ�}I��00�ޔ(��̄2��G`�_ƿ�I����w�[%p����#�`Z@�@%�ydb9�R�LL�����ԫ��w?���ى�@Jؒs�\��3-:����H֚E+���W��b�V��X�p��D�3�C�Q���{��o �~/3;KL���
�l�AL?���o}�E�]����P�4��G`[~���S�%��/W�;�llkb�M m��~���ڷ���UFu���l�f���=�ۧ�7	���~(
h�JիK�ε�]g��F8ES%]W,����7?w�i�k�N��IO
Q������
�.���0�+�k���"�# �Fb�Qd�<E�,Y����6�_��_�d�2M��,q͆A��Y0ÚЀ�yv�Ǫ]���cp:�����l��������%w�,�������lrR�9d�y�ƋKq$^��ƃ���y���m�a��B����]�kn�p�a�Ԁr[�����!�k�*���W6�D>/��z���U���ۉB���<LT��@v���J[���w��c���<�F��2�d��y'��n�=5�]a.k)i)~�X�i�W�L�;�����e؎�"�1"^������X��QP&�k ��U��Ϝ$�l[l\V/{%Ss��z%�^����ے�s�_�&�&�?����x��ET��FvW�����I�8�A*N)�*a���$�
���Y���8cf-o�e�U���&��Ӣ~Z2kI�ځ#�E�I�a�f ]Ǫ��Eq���,\���%x�ʥ��l�V�:�q2�ê��O�ɱ��<�-��������i�x�z5���J�4�s��Vx�;ǊF�!��
,���>�MOʯ�1=(��`zT��mF��)w瓟��u�\~�J���C�R�$�KIj�%)l�	t��Nc�2�R2���D�id����vݤ���?��+'��Cx�X{b�kH�R��u�ܰ������N�a�2�����U�U�,���5�~�S�'�oШ��e�r̖��b~tW�(�"�N}���(���d�7��� �����O�̴���V.4��N�.������:Nlyr�h�a�C���'ao��5�ԥ���U7�ڊǐ&/_�s'�&W+#m�������T�{�)���C�������]j��p�H�9�t<��XMI?�sR3f�@6�l]�8��"��HW�|��]ROܶb�G�Y]Q��J�sjA���p���JN_Df	|�
>ۿ���.m4������qXH��P����b"�ڡP�|V�aHVC\c�xS��Ј(�l��)J���#7���?��C�*fe�U�k�@jb��-wh�D ��@j��e�9��tv���s��#��p��>>ׇ����)߇�}��G���S�I��]׶��Yk1Gr�~�N^�I�#]]�!��Q]�bQ�s8���U8C���{��>�]eM^���8���"7�AR��.p�<�`����B�<̍}�5ͺ.�d�j��E�����'���YҘ��zb�M��X�
����_�V�ŔKqԳ��8��\������ό+������~���?�w��R,�ٰK�5��7�g����t�M�w�./�o~�'mY���8K\�d���
�z*�:�bP��'��s-��U^X��K#b�`�ճ���t[��M�x1>�fO�l1��i�`������/)A�yʉ�T��1����u�����i[����*/����Z#�봮O�a"����gH�w)u�5�x*�eN�HӸ������8��pw?��t(��UA��L�����d�k ����j�����lӿPj���ee3�
\2h1O	?P��,C�|'w��M��J��R�#Pm��t~.�xnܿ9h�8}��q�)�m��]�K�������f���xm47'N{��!���jXԱXWNn`�k��b�e��FW��:�˲}��&ovi�*��U��&�sQ*,牧ć�Q�ha�o��&���	�D��7Yc�,��tlD�fF������S�j+R�jE��-$S=TsĹ����Z��"46��Z����)�����k����0dh����h�ΐ�)V�oEO�Cc/�t���j�y��]r4:bzC[����TR�ԇ���dg�A��UV�t&R��(a�{��̲ٛ��>{�*�ߋ�*��Z��/���E}�Nr<���m�X�&q �(��:��X�Sx��D����쬥�\�ɽ\D�fFG��1�8k'6�>��cs���(0jX	>�! ��ĕ;�}~�T���C���}X�D�T�q��@�A��ns������|���^�/�4PP���Ú�&2<�ږu�W`���^Z�.?�f�������� ��]��-�rW�g`�θ���w%2�k>h��2�a�`�l$����`��qC��2Q1E�WF{e_^}�*��u88���Xo�{۔"�m.)u��)YJt8�v'N�9лX���������Y�Mwc��}��X쇏O��e�y�Uq��t$9��o;���EE����Eж)`4���ܳt#��%�y��Z!���5WAN�v�xe3��E�R���hU��ߥJ�nO�V����Y�M5pƢ�^��1�c��ʢ�()�HǓ��5��>��H��Y:��s�~z��3(���(D�Z��}��q�����ݗ[�$k�!:�8�&�`U���LW���9�����e�Oz^��k<�O�q�ef��S�!ba��9i������ԫ�;��4��x-v�<���&��@:���� ��r��ޗ������z�5��$�'���0#E�����/�����:�0!<n�퍦�������qz�e�8&lT{5�h#�����5�Lt�T�������Q�ӝ���CE�A�\`po�P�!��Ə��!-L�`-��t�ꉍ>�E8>ዧ8���D����7��OMD0މ������`X�`������ډ�=%o�R3�z����[�j#Jr�Hh@�����`^V1�ԅ��Q"q��`�m�߷���x�1����}�}��۷��{X픊sR��^m�d�е���O�ʙ-5u��R�\���l|�^�oRӵ�V쵴��~�|V�	�V+�꥾�71���')�#�a�C��Ol�ڢ�7B��ISLL�O�Q������� ��)�mh����G� 5  ��IDAT	^Sd���F�M �Y\He��6��I���-'��1!�R_�\��S<���R�r��ט��A��+NHϥ�4�Eg�*�k|����:�4G�e�1��L�ϊlP�AI'�5,�JB��M9F�́�q;�t`=wqm�����z����- �������=J=dJ���C�,6���H�(�	�\Dy+HCa�0�L�x����d�>3��f߱y�M���-y����]/���`p
=�s_���~��.�i����G��Vb�Zi� ��1��A$24��b+�*����?��m|a�ʥ)����Ǟ��ڴi ���E�A\'��Q;a����i�m>�����ѕ?s ��ڼ�ɫ�Hp	2��I*\?��KE]��V_��?Pa�aKt���m��Sy����*Û�<j�ǌ��
��ګ�޿��s�>m^��m���x�-�F�����s6��:�Ns�0�����e_GILi����H�h��_�[�?����@c�I�-ʗO����٢	R;]#��/��fJ����^�	���+�G�+�%�Q:~�q�[��ĉ����xi_5%�6���Y�N�˙����]], �;��o��6��(�K�i�>	��2��D�x���d:F&�H�Sb��-��2���TEo�p>q�N�!1Y�g�)�14������0�l�t���(o8�8M�j�p��%��.�|�F��Lq�LL>S���X��|��>%��<k��Xօ����I��E;��ê`@����.��9����E��^�����DzT6$����t����Lb$wj�-�Mۢ��++%�J�/����d�;a/r%e��^�mr�l��������L8��E��F��:����`HЩD�d�5G[����T���qLq��p/=�E��������q�Gx|ٱ�oŴ��r)^�m�/p�_�ڋ)p�P�jl��%��R�� ��R8���j�Zd�7H`w�����JH<<_k=Ã�΍{����iG��Y�����h����$,u��u�����\Q>7�`���HM�5�M��N/��>�M�����:��3�[���>?���C�IZrz��0率Es����.ͨecu��Hl�����3�{�,]zL��K�MJ�kSw���a���CvAd�;
N�Y#K�i��r�DO� �l����(--Z_����q��*��~�1X�+�e���HOaZؘ��o�5Ґ ��4�C&�;I_A::&�XL<q��<�GE���U��k�O�W/�
kV�R�$�"!���k��<o���"XU��Ś����R�=��,����T<8�Pa%
O�J����޽$)/a.�XJ#x�^�l��\�X��ٶo^w��_DÊp��g0]�;�M�+���)s�Y\����*�A���BV$jtDC�H�	�(j �͜���%j'n��頎	s���dZ⦂f�O�)G�tc��}N?�A����^�/ys���7���Ep��7��[sY�=�F�Z��s�|�m����])=�s'g�5pa����g�">#-"�7��%�\��>��=��J6Ѱ�������'�"�}���کn)[��4�]Uq���E�-6c�ٿ&��A��C6(Hў�H1��C�!��agmh
2s�u{ߏ�����A,���S'`Vއg���]��G ��gk�Ȇ�t�v�fmd���[�9 lf�ގ�֬�Q��!�9#��l�K�ci����&&��� u��Ab�(zē�y�C/}�k� �~�,~)�St�������`Gׇ��q�����'T�W������ �F6��t�i��=s�ڪ�NZ���՚0v�lB�mH}��'�O�P_k��]y��S0AO¤�v�M��RC�y��.��$�������u�q�`S��g�X5I�'x>W�x<�Si|��'[sAr���#�*�ʖC�Z�f��cs<.�����)�!]Nu���|O}�m�W9���l��z���7ӕܵ�'�j�.�7a�K(�LoGs/�0"(7��"3��1_#��m��,�ρ�⑬�ރU�>(AӮ�ǋ��a�Z�k=���2�t�j��@<���m1	���;&�]y���XZ�YC"� �*{@�k�k�3�7�x�q�f�*�f�U=]VD�F��	�??���[������`K��霊����ݼa����7T�f]r�ɴQ�Y�` W1���9j�H\����0�ڳ�y�V�Z�L����{!����57�+�����ӛG�A\�_�(�������`j�%P-�'���aS�!�o����]k�� ެ\ܖֳ琝��k�g!t{�w�qp�eR-s��|J��6��u��J@��sww���Tw��pUL����.9��r��4������ڭ�"���V!���i������U�RZX���р��m��K�MO����,���SZ������&��d�¡<��kX�����	6V��8^/wJ��Q���q�M�_�
��ŋ�j%=�"���)pT��=]Yj_��C�"�F�GRK��Jd��ķty�gt�CZ9Q��9�����
g�]���˿j��[s_}��$�������Q��#@]��7�HI�qow����5�X�`�$���I�������:S.�/_�G�ş�n�'ۉ~[B����p���?7��.4#qmrXik�y�����&`:1��m~���u�p���6�������]�J6wv��w*]�A�oE��+	���fVZ�fv��T`b�B�o�<�Z�-��ɥQ�m��>�ΰ7	��^gެ�����luLӺ���%��?�`�T�J)�����i��*л�,(��+Ŗ)z�u�nndZ��l�V��Y';a����(Hm<3�~��g����{�oF0ؾ��tv
��X�ȱ��'��F~�Lai��p�D_+(�
��yӣVm���X+�<��G�[յ�'_ه]`�=7`��t	 ��p�D��*Y�'�a�N �7�0Q	����I��R15�G7�܀�RW�1�0h�cА�S)��s�YbIݣy�k�uy|k>?���T�5��1ڄQ�
�#K��XFYu�9���$��ꃲq7&��ڍ٠�m��1�/���t�F��ʪ�z����xc�x%�5���ᜐ�ݘ\����9���r��$�ȣ������TF��v�l�V1.�,���*94��te�74���J��������^��s9w��t����W'��A����z>��6�|7�P��(3����P;��1o.��8�!��Y���^�*�d6���N�}yj%���BG@�ٷ��	������m
������'q��]��sQ�Y[ܼ2���`�eł�<[a��swS��
���*9b{w(�Hw��>�
R�}�;�g�w�}�J�v�p�9⹦���	�u9�ɘT������-uD��U\�yݾ\�.iHǁ?Uy|����#�R�.�a8�IUת�׈�,�Y�S�@�k-��jXثѺ�yz�3���Um��;��!�?w��w4�f��yNۏǇ���|E��ӾIF.�}SԦSt
]�=�}�;Á.F����)!�Q�~c��X^{�S(�km}�H^�y=i DM����H}M��q�`ɉ
N��~�m$�amgt^� �K�D��P I���-Z+��Sץ[�������Q�������/�pnbg�}�6��QJ)!�i� e�xMa��d5�>_dB�[V��U'���(KZ[��V���f�Vu�yqm��]䎚���Ȓ,�#��]�{M�8�a�3Ŷ�m��n��=qPA� ��"� ƍ�[Ux�)[)J�
����c1gXI�Wf��[�y�"�^�o�A�
������u��׊�z�; B3����%��/[Y��?��C�x ��d���*rb?����'���A�G�B2�p_��[ ,�5�F������Wb�%�X�b$���Q� ��b7��z?d�Up�J�{W�d���O�R�/\W�w0�u�8�� {`�>�i���,?��Lj�]��D�l
[ʜ��I;د`>��Vގ�_���н�#/��}:�q ۵�������0P<)�}&a�!�rܒ��>�~�]~�q���?,E��.�;��D�"u��0�e�*Y9I���p��r4������>�e�M�]�6�fl-c��_���&Z�hJx>w�)�f�)𬡿��A�`Q�+�j0���Z�Ɲ��͙�婸�'�ɹ}a�n����9u*�i6����N����������st�n�.�\�x�x�j+k+[XN��!i&�5�:ϵ̟ĵ���7uU0^8���ڭ�nO �}����6�o˻�]V�p�8Y�J�Rljt�@�Q9�|���-0�\���T�m���O?FF���p���^X������s����&!�B�P��k�D_����O�7�f����b�Ŝ�MHn���� z>�����JC�mnl�Xo��s����b�n�1i��
�P��S�Ӌt
�')�6��a�Ǜ�M��%�?����㚮N8@�y��6�Sd��>~J?,�����
E~�ݧV/1 �/QN��Z��}���~/���EAu�W�����'�8FK��,J!~�z��.�Տ�fS�W.&�T)�hjO�����
�u��Y�ˌ�-z��Xe�~>-*�FM}36��{��fZ].�1��>yr��k�	,��E �\Hӫ��݈����>ˎᄾ�&�z`O�4uEϘ�Խ�<�&�sc�,23�̀l6Tp�`E�<��]������M���{�m��u?cwK;����i���	QU��x�)�����u�^bSQ5�$��.&@�x�{��n�O�yx��<d_#��o��~��~_|~���!s�����M�Ʉv*^�I��*��ľ�����35��b`|�5���o��\�&͊����@�,>!���n<�����3���#&{`���2U\˷o����TXz��Y�k��ÞSZ��m��)(;8�4�瓦Ӱ��7XcȲP�L0G���n�0�lf�����a��E���D6y2�������a�,�|Tew�:�Q��@1����i�K�®�ʎ�h$>߳rz�5q�fAO�%��z̓��.5s/��И�\�jm�����6��ܟn1uM�%|���������GПn"q)�/��V�hF-�B�tSd�^*��x� �T_{=�ʟu���S�x�{\,f�]_��3���m��e�,_���#�)�3�":�/�RO`�E�!'�,K	7�,J[�ܐ����@�B� �cO�)��Ź}R�P:���L1Ϣ�U�I�ua�g%ot��a�w?�9����/[v�6:��;'���ӗ��Fr����*���ڟ5]��<1����ǂ�츯JE��K	6&�N�n?1����{���"5�"j�7iR��]4��"7C������H�Z����
ig�O���z�������J̞�7d7<��������'�E;�����[~$��]6ȴO;7<�z�h(�ؠ^���?�i��a=��0��-��J�.�����"\9'��p=�	`�׊UcPв��ġ'!��f1z%�o!�u�>�F���ե�]���3��&�2��^Mm6uk�d닧k���,j2�f_�/��N�d*nTi�ɦ��=e��P'�i8�+�����^䦌1C�����@
��G
Q�Q�#nW-̢�g?����\2��-���3&7�,eJަ'JL�vy�bR�|�����uRC�J�r����fѥH'����)'��^p�~�2Od����lY�w�G�hm�^b6����"�� ��π����ӖA��e���a���6�����%�^)��Xcl&|6yQ�f����s�����ރ����n��.�q{����fc�iCB<��u�:Y�<s��lBxw���	�p�wm3��f�+�%�5�O�/xN��}��`-,U����E�pW�x��	����x/�X�����~��Q�@�b�7ؠ5�t��r�l.}�w��Ĕv({�[���������l����{�j^>�]���R9n�#�{�`��U!�]�MתlFiF�����|�Yέ��YX]���/�ￌz7�$�B�ڶ�?۵ߩ[�ܯϩ�khG�T'Tz���Hh�p�[E��m��O[��_`$
�]g�P�]��R�Z+	7��,w9�rUV�At���q�o��J1��e̐Ap�q����n��(����,�8���U��Ͳ�16�Z���lnL���\No��0�B�m��+c`˜��i'R`���}���{L�(K
`{���ͷ�_~�;��?�xf&�X/vJB������@*�
oW(�qw�4틦�0�P�W�!h��-d�߼�ύ��Γ���Aim�*���`�]�>�uұ,Z�/��U��Ն�>x
�*a���*�����?�@���x���Qe)uvEÁ���92�����w���=����tR�.�sL���������Il���	���[��C"5w�믾�����Qڢ#�E��V3�[O�S܀q�|�z��ob?5j�^?��C�,�	;�׋�dM79բ3v�2Z����ٻ܍m��_���z�W�F��qõ�t}Ѯ*�	�E��Q�^2W������c���0�2f�j��^��K�ِ.�J/�z����Ew�d`���U�X�OR����.,8��l����	��5��No_�,d,��"��̪H�#J��(�հ�8�7�F;�-���U5��q�<Q�x��
6�n��)��.T�a_�^���?�#.�k=����o[����_q���[��t�9@�~�6۫mc�wU�8J��:�����|�!����|�Y`��j1���M�nZ4�ο�Md�x��<�(O�E
��]b6��.�A�{��ꫯc#c�;$��8�������zl���b]�?�R��_�5��-����)2((ɿ�2�����L�5��k��w����ۧ�I��z�a��!A��t.�8(��:2q��ή��)��&�(Q�q{��"[�5�z�H�N���]V�=�P[l���5�kb�j��"�w����aOS!��OмA�mQ��̙,�E�=hdMw��XsQÉ@��v_�i4��Ϧ{wP_ƾ��* Lsf�)р�����Í闻�]ߗJ���ӑu�j�n`���;a%�P=qH�K��dR�-�N�xl��a|-R��_E@�3e�3�V�1%�ジ�����X��C?gwݣ��i�baFᙶ�-�#���U\�*(;7�c`�w�T�!efMz�$�<Oq_�B�e �Q�W<�Ο߿���6���xV����#2����|z��#}��J���x~Fऊ=՗Ne�5B@C)�k�$K
NBu�^���Np��k���t)_lb�Mɹ��E�W�/)}]�d����j���(��c��d�i3�h`^N�\����|���=l)+�g�HMX�S#��z��^���}�h'��vYk��pN�`#�pܫx�ۡx�2ЀKcWf���7����L���}a��C��ￋ���UQ/��k	�z��7�07=!���}� S�I�S;�p��Ly����VIڟ�����[vѱ)�����d�	r�L0���6��4�Y��_wg���x�~����� ̆JrY^T!h������R
���b3��e���Sj=�\\D�GK��b�=E	q���~'�5�p���<�<�1�Z6A�@���Ӯx��oP�N� �62Y({��נx3N�sNjy.�ﰫ�D��u�A�Rg��w,/m(f���l&��>||��ݲ#v�?
���|M�"6��A"���2X¿�Cv��{U��&.8O[6����p|f`��`�~ձ����3�ٳ�:�p�m�L�@�����Dbp.UbF�NtW;ĤwA��m��u]��X�r��"h6@���B�Tk�A�*=�):�o�w[�AV�a5|�; ��Hm�v���h���!��������Y�a�^�D[��{�0̼�z�a5���D Fј�� "@聆�Y�^q�~��|��)��Coù)��A�l�3���>M�q�p݂
6ŶP�>�R������ �� .k5����1�`۶SA-�?���1�k	��OR���w*N�����ڑ=g��X*���P8����ӣ�蚓�4��r�j_.RohX���)��Q�`�6
6��\(�_F���������2#e&cJw��)�X=i��2�cv�俍��",��C]�mV;
|.�aR�n�˭�3ϝ�Jc=}p|.��i�;DV�L	e��ۿ���r	e��X���:�����E��.=�)�Q���D߲�k|�����T��LB@�1�Y]PT)����<����	��.
�,	^��$|��7�o����r��n/�Fb�'��N��|X�zT�x�*�N��wB�8�8W�Ԁ�&����������m�\�k�(%��c��~�z��m������` %���5<���c`�j[�d�����x0�0�n�s��8 0O�*�q=�1�yA	��{{>H㿷l4���U���N��%F}��p��Ʒd`�վ���E�9�l��lR���RӕU{$x��$N������Ju���}��|[/M��30�����f���㒳WL�#��X]��Km�1T���rYʈ1��:ҕ�������Uc�&"⢮jRQ�T7W���Y�F�j|`q,���]0��sGv2HA���k&Y)ksP�e�.���]�T[�Uԑn�%S���?���ߛ/�����+���ۻ��R�%�_\[�v�8�vsF06Nk�P��+�2p����r�2�̗@G�ཱhd>�n��K��Zm-'��)�WB�����<<�.�ؠ47zh?lPuy�өD�Ͷ(+�	{A������,�ל�_T��`����١�I��ڮ�!�V��t�Yz,_H�k� ���w�Q�f��z�_"��p�9{�MơK�cP���؜��2�iIkp��i���h"p��X�n�����iX�s6ׅ+��x��:����g�J+�e͉HŢ�T�\�2���jx�Zm6��M�|���"֟��V�cMN�^�-U�,��q�q��L���h�{��j�sN7���ܔ(�/�8�x�g��6���5&ya�nj���|�%�{u��n��tΟ娤����[L���@5�벋K"8a��I�]�����#����e�k!X� �ed��6=�6��^vc�F%����5t�����K���6�,͝��]�cC�(+ab�U"�bN�@}ZUle������'2�!�����\� /��&���(�l�5��k�X�/���Ы�#�f,l�����#1�=�{O>dۋ��Ş�C���E�2r���Z��l�H�S\h�E��}j�_�f�E���6ꟺ�]��X�rL���^:���Ս�OŴY�ly�B�K*�]�`���S���љ��D6�6�qJ�>�*qx�(�r�حu6������r�솲��T��p�(�X�nn_�٬nGu=�W���5K����7׼��������u�n:B�{X��xϨC8!� '*� �`���A�V�0��ӧ���Y�2�_0���s�i��(b��Aa�=�씁Ya!<iƅ�7�K~cCbZQ���4��Ih����7ю$9�E#3k�{O���CJ��wλ��9W�<Q��z�7 ������<�0=$������%3�����L߱ #�>�w<�B�S����d����NDK�ÀGv�d7ު[��(dX��P�Xhr �C&����$�c�Nоk����W4�۳��谡�� 8��9\O��ht�6�X �J���C�KN�PN�<�1�.w돇��b��ذZ���8Y~�����EƎO
�5�3��Ø���|�1����|��؉����z��vbw����T��	��:��DUB]Tf[��K����f�����iy�h�����8hl�eiOtV��!�@�=u�sm��$�q`R�gO�ym�j
+�C5�;�
�n����3��r6�v#�6G�T�fuФ��&�⋲Y7�fą{2nv��MU(n�!"WY�?�L1��ǛH��@����`�����E|Avϐ�?�P�?j�����.8k�M���P_ҁt�>̱h�z䍴C���a��
]vR�A�:���o��?|ҬnH��[*��6�b��R/�es��ڶ�F �ȭ�f�{s8~҄�j'�M�x^Q�Dt2�Gd�UB�R�5\�)����ԛ�k��Y�����?��%9�QHZ4�����p8V)V�>�+�oKd�;�.tW��ͫ�Ff�(�� �h8İ16y�1��㬌%~�y�M"d&G���Ģ�<�#��>��͇���q�{T��CJ�J��ðո�a]���\B�*��!(2��Ngf�񾩠u,��H���^M�C[���A��Fad�de��۞����o�C.|b���v��Mu�C2�Rk`g�j�w8�=��ڧmTV1ew)w9���5�N���:^3���Q����Qb�$�A��7�6�.5#�Vq��gU��=j�ڕχ�_��o���Ɏ�J�Ƙ4�|=n$2P�a�	!z�Vb��4Y���XbQ���=�8�R�l.*$��.F��领������������&ZB_�4��l՚b�����gYJXޫ�l-�R�c�AM'c���u��5��>�B!0�y�V����:lrlp�����X]<������R��G�td馋��X4��f��(.���#��`"F^�)���]?�Sp'�/���u��j̹���M��eנZ��w4Sb�(���QNs�F�
���fW����F�7ŭ-s(K���������c�gk ��g-�{�/r/�(9�;k]��6}/qg��r���%9���X�?��l�c\ҜKVg⃚�2�\�ݸ	Z��%�h��kZ��'�s�	�j<z_�t�����Ic�]�WafM�7�pC������^������ߖ�7��9��nU�z,�r�V0d��Hz(/�gW��M#s4©q�Ձ4n�^&���c�8���T����}��c�F'�P.k/�m�rմ=߷�X��L�7[(�x�0 ��6��w�'�:�J3)s�C�$����U���S����F��]�ߛ���c��G�C8C���*��3� �C��oR�d+p��9v��60o\�,c��R��ﾥ�݇��s�c��� �g6�� ��$��M(�S�h�/��uw/\s��Z��*�ۊ�wS�z�%�~���r�4��'��>����ȵ��-J�p��47��S-�"��@�m`n��=��cm��������H�5B��-��.��)�*��~�<e\�,I�lhv9gm8���xT�h��(���w_S欁Wh�e�z�s� ��oO_�}�&1�V�~=2Ƒ���e�L-�~���2?[�ڨ��\�w;5w�`N�B6	o���|������ÒSCn������9E�e��{H�Wd(t�
��}��x˦�w\����h()�6����_H7a����Y_Y*��iX�B�K9K��Q6�e���'��;�usOLg+������	�M�&�Κ�~�,�e��*�X1� ����ÚA�Sey�'�1�>R�!}Ĳ�'kX�X��Y��s����h !As��_]˹�{��)>[��O?��֌�6p�;M��WJY�V�tN�/2t\L��$�U%0���"3��AH���[`�a6�@�d�O�<*Ϟ>-���M��������3�A���~����π��F��&�s�w��|�}h&X.��/��%��@%��>>��{��A�+X�杂���q�b��vǻnІ\�!�Ɖ���X�Ҕ�U=�،,:ܢ����m\[�W_��������睆���3���@������YD����yZ��2g�N	%`�Ą����p�sɕ��7K�����A�SO�4��ݡ�<#�\o��g��˽Q�E��n��Y�y)3��B�����,�Stq0Y��*l����&|>�C�!���`j������?i����(�R��ϧ�X"�Z	_��Џ��y�.�Dʹn�,���xe����Fą|�_/@)h4�ɡ�XĿ����{)��<��v�et�n���>%�9��l*.X'���7���?V�aY��`��b��2��Y�H�G����	���C6ъl���FZ)��B�&1�N��^B��ll-q?}�{ALmmD}	O����l��gO���E�$�6�IuX޽�	� �k6<n�a�!NǊX�Zij�E�7�1��͖<�	�������/��v8D���(�Ŀ'����c�y�IC?����Ա	u�g�|&��)�m��K���t<7��`:)W�I��7���>]�׫�_�#hg�z麰h"K�S����*~I����Rg������ù�?��[�3�+�cվ �����~���"�B�J�]�hJT1Ux��R����H♋���%�D�K-��n��E��Yg>U�����b�F�m$�HU],�p�u��d)�v���z�u� �����>��V���qf�2O���b�*���F��g,��E᱐��-�E|�-躼�g� �H&-e�$<A��{[;l�Re�Ɉ��{���}p��$Tsv���)өx�')t=o��=�Y��k��G�m���ML
�6���	%=�(�G��麰��v��-�����v׌�~�O�3��[v�����>ǎ/Sm�13�K�4���}����1$W*��X�g���a��1;~��gF�����Ԯ�+�ހ�4Z�lf�Z?K�n��(��Z�;$���u��&�mjq�.%Thd�|�Y8�r4佮����V����B1J��vw%���8���?����L��hr!���a��3������;��y���w�{M{Q)i�E��s�g�"`�:�t� ��a�����b���J�䶻ٕP�?P\z�v�Kw��g=��?���!D�R��b�@��7�Tļ�QĦ�hsd֎؟��N������p���kz���G� 3���HUM����d`��m�D^ه%�\��Py�.$�̙�R�w/1b��\8sb�f����8!��Ky.�������i�����I4v_�ad}�p�ߒc��	ܰ�G�BMPY^ pK�h<�shd����HѵݪQ������D���e2�=�HnEa�/��,�}���0Y�vn�D��Z%>#^Rp�n�BG�:s�JA��=��~���0�=-�vni��N|�L�:��B��Ӈhsؽ�4���\0Zږ�KO�9]�s�Sv��=w>�PD���;+(I���n����piX��k��k��'v�q���5l�6���B��Z[��n�Q!���/2r��b�������_��G�����e(�c�^��������!~_�v�i��s��Md�����P�f<M�Wؕ���S̷wwj����ǠL	�G;�)�c�;��\�pЙ�=(���Um�����:5c����<�0l�Tk�>ۨ�[ԅ�8��N���*T����}�4`�Ue�ӹ��I'h���:9L�wY�.�F��`����/^����g0%�l��:j9��k��MR<�u�,�JݻP�	%`�&��>���l��{�WY��և]��Ԭt�RŀxP����}��-��	����������&��M_���YVx��M(0 ��<)>"{�$�9�_�SlX����wi͸33`Sd�MW��������zp�9:e��	Zo��p}�P�qg�Nt����!xS ��.5
̷�1�m�m�|���tW���1�d6�%�6I�Sf������GXM�< '��x��,��s���K=O��R#�K�5S���g�d渎��?�@�=9�g)���i�Ǡ��x���)�^�l�^���+: �b�ؕ6&���%�����g6c�	B��uo8v}�f���'��7q�=�)��"x� ��W������/^�(1hpu��.�MQ���*^Nh�Q�c����6!ei���HC?�c�]�}o9�~��� �g�45rI��W�:6f����,�ur�� ���&5+���(�X��(w�47����3���/_ds+�����R�+��Rxc4�i��E7~�QjQ]�T(�ww,c�\�ww���U*�7�Xh\�`&��6G,����꤉[�x�	��g��[�5g|��^�%�]c���L�b���W���^W�om9d7Urx���H����3��k�t���h{��F>赳���HP�ر�?!SY���J{��c�n&��]�hVp8a<�ɸ�\��$b��]V+�0o3 �����f�4-�:�*�+Wpz'�Ų�F�m}B��Pz2�g&֏&�u(�o�xS���-n<+Q���|�*`Ff��^6�P����J!3�����`d�\�}�O�eC~��s��k���̻�Ae��rKxL�o�344�!���C�5����R��*̎V��Ϝ���:`�~���z]줳0H��s�6�.�qU�jB8`Uéݯ��{!�ll%~�y���(�q$�l�&g?�JZd����|BA���L���d+9@:�� B��(����8k�T���Rl_�vspc�_9��t4���|�HR~�9Wou��Ʋ}u��.��.}32WR�$:�S�~o�a =K	����Pa��.�MOR8���4�(p�f΀\,���G7������QY@�w�[7Y6/uY A�~�f�xc�d��,�4�	b��c<�f]���#˾��d9�Zt U�z���^��%���a9�VSI^g�7�s;Kt���(��ʔֳ(�(�}�9d������pד�QyD�����NA�_�i�u�
hx<y�a���<[��ω1�9gґ�W��T<2"�F�ac���	`'컠Z�M�����JW�NT����۸߸�'�y�n+��C��D���b��Rg��\q,j��M�Pe�*4�Խ�,5;]�b�a>���T���Hu��(܋��S�vRL	��:5Mw�%�N�ࢮB�Į��(�������1.^�yB���M�v�,�=B���=����5M�����l���C���M�2�� ۊ����ڜ��ח��X���!�Z%f1HGI��}�m(N����*��o�r�� ��%e}�w��#@�x�Ic��3);C"�H�BQR�y���^fv�1~x�y��h����������85��[Q�(���݊wh�9y���p��}��]����e��C% ��jpѼ]dn�y �� l/��
�F��V/\�̈́M���FMf�&�/<��n#�RO��c`7z��u���U�c����
�	K����C��7ڡEם�ߓƅ�?���i�_8짳�n�����r���^��� L��G�5D��Z�8XE5 �>��{��)��5�͈�+�n���t#��Ŭ�gQ���H�g�L���A@��R��|��Wc�u�Ր*�g��t�����z�Χ|5��}��r
qW<6�4�P�C�bbsb �v��nI�ߙ2��꨹�����K�rf���S�(�6�)ox{�`!ͱ�lK˃B��i�ԣ.w_����M��h3ITy�3M�þ��,_O	�6�w`H��ρ&'y�!�V&�/\i���G&#{����'�ի��A��p���m���P^፦�n]��ۻ�Qڨm<�T BWl/�U���3��!>�b�Ae#&0�u3�����m���9N�,ߙ��I]�K2�.��rWt]�8ƽ�^���N�D����*�Z��Z����m�g�� *!�!=��Z�R@�k�M�e�,/����6�9���%6XS�g77�ym��9�]��68�>4��OЮ6�R�~b��2��S@v��E��^C1�2���@X�K%�{u9�{}���"�hL�-D�Ў�me�
�AF���.�b����ܴ�3]���YĪO�yh���YЕ%��(K�H�3�C��f�U�ߔS��%�����NQ��Xv��jJa}Se��ϐZ�.�p9c��,V�mCa9=�}�$��ӔN�'3��/���)��d�E��bj�T2���\S��Y{L
K6/VâL�����Ds�]�wG鞁�/v�?����͵tfO�u5���j݈��Az}}�g�I��)-����������w4æ�"'�M�&�څ�!�f_~��m�@7��:o�f�����6�:;5\c�a�6g��:H�8�K�7�ᖓ\}4~>���qL��>⳾y�[��qu5bb|r#�{�8��?�:l4���r���J�����B�O����X��>|���I���As�7�ٓ�Gu��F�-�	c�8��䣧4�]�7�r*`�����^�&����C�'��/g�Kf���))KV|@�^��/T��R�9��� <���.#�΢-���2��w0�	�E`�Qf�S�R��{�]~<B]���?-
�]��@��j�f���S��n����e��L�0��'<Sq������fϕ�˰>�#��S�����`����HK5�S��2��A�%-'��M	8Z���r��R ���Gj��8Mvs��'�n���7�������tNz���;��Ca���{c����"��j�K��%�L`ӝkL�B����\��֌�w=�/�����b,����̒ڸ����[�LJ4B'�x��,�*Q�;���~TOذ}��9�^�~!�?��/囿�����i�ɣ���p������t߃���Ǖ@������{��2t =���Jg��8�9Q%/3�ޟ[�qg;p䰏��F�9V]�O&�\�dD��h޵��o��v�`Y.��5(w�/���b]�+ي)=�H{(1�βL��M5��bx��y��nZ�K.Y��U�,`�]LS�"8-��j>U0vٸ���٨9��n��є�Y�o�UF�;
���}��7�^u��9�Ug��-P�}8\��V�y����5pg�hbB�g�{�)}�%���5W�ì��f����aϧ-���1�v�̀�,��O��M|��q��W�^�R�����Ϋ&Y��D���Y�؅���b�e�*��s�Tj���%p녝�+}�����e����_�9��u;��?7��Z�8�`z�_+�6���*�_g�
�#�#�Ӓ������`�}h<���~�e���_�Z��7�Y������'�'���cܛKV>�$��4G|؈�Bh��u�����|x���Pw�k4,�܌�S��9`2$���j�S$1c2]�خƲUV�m�͗N0��i�6����T�.�e����^}X�����]{���\�I�n�@��]�Ml�5� ���4�"�&y�Ys��[�s�k{v�%48l.�-j����i07�qHuO>8�59�z���T!���%��=y���"�kP�%q��4��<Ņ�Qhӫ�b�,�>�|b��C�$W�<���ܙ���!7��Ce��I�T��C*�Ҿx����sgM�HՈ�����8*�o��#)R�&E�!�ls�!4*����8�1�J3�T�yiǏ��Qz��� 泇L�w�]�p^Nw���J֕��D�r_��뻒S}ь�T��G�ݒ��xF�{'�Q������7>:
�e�i+^i�R��'�t'd|�ʗ	���o��a�~�͟yݠ��� ���͎A)o�(��sG5r�.�Ȉ8�ޡ�Ϻ.0m���O�hl6�3�������pfR�u��aY4�s]�>�u�kI %Ľ������� ���ڔ`���U_<;ۢ��P�3�濐���P�YQ��n����\����]�t�$.�L2p�%��2��O��mb}!��w���m%�jb9����y�/������&��R�?gg��O(=�|Hl22B`R]�8��a�?��}��;�����D}�$1S��Rms��1s]�q�\ͪ��m+̲D�U�T���f����Ec�t%�M/5�א��o� ��a8�S�^\_�0*�]���hT�rR�'�{`��:S�:�m�+iX$"(4��I���n�θ��c�9�.�;�6s ups��o$�k��h�o|F����ld���`,��5�h$%�ˈ�3�E���C�~������R����@L8t�˗_~������4�"��S}-٢��ؔ��@zT���� ������勗���/ʣ�O��n���gR9\�/��V�����p?��B����ϼ�e�����錴�-�PT����k0������h����l�T�J�D��_f��T̨�����0A�_�Li��XpΜ�X/"���挟 x߬������{����Qx�=ţI�x�q�)T�?�z�)$3��]t�,PHǅ��qf��lsdh5#��jg:���9("�.��B
�׆Ї�.?�9�uJ%*o�!̬b"]<��b?�>KEV�'�'%�Ɨ���j�&��h�񉮘��F�S�L)�7.^i2�R����3�E�n��5r�������
b'�BLnͲȰ��6�.J>褶�67��f(El�
+x�K�W����{PE��&K�m3����ʢ�7Y�t	1x��H/��f��1�m/x��<z8͡&O���P��! e��/w�i?^�5Ƥ���'y���g���c�Vm��lF�t�����,�ǆ 
� �[`'J��%{�}n2�h/~]��P!������}R�l4����Tw���3�_d�bL�*i�m����_Iȯj��6`9:�����.}�g�L��X��Ew���B��
��$K�,�{l�&��T� 	��&�z�,���(��qM�
��_]O�Ti�K�MDl���y�q��~��.n[�����xN�V�G��t.�۝/Ev lWQ��!k*��M.�>t:���\��fS�l�z��(Ê�#38��^�Ao����'��Ԭ��˭��B��FUY����m�p��~�����̞��f	8HP�6j)�>�x��Vh,u��rP�������1����M�^/���)�C%�k���`�^��gyo-*�Q��,�a��yԤ����~��|l�nc.� TS�d����
Hh~���������U��@=���:��]i�����'0���~���Q�;��k�U��Cl�����Q����:�1�RM6��Y����jΚ���o�l�(�k	կ���s#a�c�Kf�=�[�@���qb[?�;�5SSi$���$^a2<-;�c�c�D���S��x7j/��9 �qG�������<�8'�r2t�D���J��R�!�ʲ������E�ϒ�<ϒ����� i̗__��q�N')�ܒ�b��ˣ�kBl +��u��e X�|��*<�y�tp;�)CQ�3�����Z����R�f� �����i��Q��	���1�6E��(9��Q��H|�[3�]	a�"c�M4�'�RJ�Q���j��Is��&�*h� ��v�2q�7R�u>���������Y��ZAs���J��)/���M�z���ܿ�aJ�'���d|�K�0��~]��g�V��φz��5@�f�	���۷l.=���m�Co�	 X�-��ޱ�艳��YM�PI�C�4�[�D�$̀b!W�S���Y�Փ�����<(y���ѵ_D;��`��"�L<\	FFKZ����<L�q����_����@j|����T��T����6�H�Klf�6�x�n#۬�(��Xﺰ>�$�'N�Md	x};g��,�M�}��������f���5*Q�8#�8��Sן��d����k��ݐ���@Q�Ǳ=5g��ܐT�J�n�g+��ؤa{A³(K�_�eI�mp�c��׽����A:��o^_�#MM����W�����:�GRrpo���.����<߀4��$[3&� [Z3�kQc�<]���f���#�>"+��ב����$JZ,0)?%n�N��%� ��*��Ǵ�U��9�m����?� ��__��ZȲ��p# F�P�<��w�/�:�vq8�b_o��t�v�
����(�C���k���Uy��>�A�'R��C�o=t�ѥ@��_��_tpt��4��i���1�T�`P�hZsQiG8k�	I3�R-�&;��7�n�e����^���)|bӾY<⒳���o<����������w`�%�HFj��I�/K^$/�(�TڍuF��7�X�U�y�sT.�������(��	�c/�Q]͘ư���Mg0� ���G����o�q�@��m�������0P�� #��(cn�򴩴���Ƹ�8p���,�����v����g����,�<__2�f X*��aX��O�١	�1M�I�s8-2�̶G���������W_1���p�!��`0�\��e��t�����!d���b��fE�A�ޢA6'��bfe���P{�$�Tt6!�Q�IYL��NT��TN��'J|+�Vq�O�	 tT�g�a�yz��B��J�Ð
[`\��H��:����n��:e� �P���De���~����Nl�]�DŅ���ߕ�?�T��O*_|�"�t��@/���˗Ϲ�p���:ʜ�Xd������퀣J��&kV��uV0���nӇ�~稵6K�jIVG!4H1��0x1l���cV�K�5�jcƾ���RfM��3��y,��?g�;[��f�Os]vG�@]r�i'���f�40��M�(:��&̚��@'u*��e`�cJ�cHs���$<��{G'������I�f�m5�H�v�B
��S��=d�J4�I��1��!����u��t��zV �]4AS:dF
[i��w�ҕ�9�eZjCd����t� \�=݊���!v#M���f���<�I�G������P����=�s�_��k���oZ����`���$��Y�aר"uY���+�sw�F9���k����L���6�"��Y�.��Vܶ&I�G��F�a��;��.��:J~�Zv�E���KG�g��{�dR|VV<WU��U ��!�f�9��Gj��,�ϲs�d�Z��ͷY~���Dd'�:���������?�R�3X�����%���&�B�<l҃���� ��m}�Q���?SO�_pN%i�Y�0��J��д(�B��ov��P�v$��J]^��hV/�s�e{�->�m?�&��T���<RO5Y�jR���S�e�ZՄ�/x�I�fq�3��1
�%8k#
�#�qc���$o��I�&Q�ȒX'���P�����/n�Q�ˢiJ�"F3�oe����	@� 4 Z�!T����Ff�����$�X��H2>_��ߤm2���w
b�އ*�)�c�@Z�l��Z��N�4��ʦ>���q�`�o�����x�u�d��������� ��s�ϟ>�pP>�cY��u�Q%��J�a܋���sS�;>��'���C7C���ǖ��!��������~���uX�\��->�` �E�7�$
jʋ��lN�Q!ߡh�Tr|������1(v	���0C�`{�w���tF1�I���I�	�k�Y4��CI��������������tWEtD� ��jGK嫫�`���9t(��=����CWԤ��q�&��N���D(�Ue:> �b�J���d�P\��+vl`9?��PɊ��yeD��V��B�^��ح榳x�x�����Z\,��&`lٷy��M��\Pu�����\-��.�ۛH�!�o��聉h����]�n�˼������4����,;c1u�ZQ��Z����I�nd m3����G��P4��)'|���Of����lP���O�D9�Qٹ��9="ˆ�?�ݬ����=�D'�{Xb�k{n�/�|�a�zٗ�5��=���r<?�I 6��o��A����ޔ��U9����3��_�_�.���o�����J��=����|ï������v#�dx��l1��Ϋ�H�`z����c��0d���7�	�K�/is�A�,`�{x�A[*�!��{��P�l�z���r 6ɽ��)J��NCW</[)���������7�P�z5a!FB�,$h=)��?��
��x)���5���t����C��S�O��w�>�#	��X��|�H��ʺ?�Y���2�'7Ot�~��E��ށ����9�to����E`^��}���3$?�ٟF��M�i�]�4���:WJe �J��=���]w�����׃��������j��GK8�#q���b%M��q\P��4�T[f�^u2�2�+K�j#�,���fLS\pf\�$S��+��D���mLa�
D2ҫ�7k�P��_U���ØD��R#�s��yR2��Jz� 9Dw�n��4iќs�۷(J;)ȫyR28��o�Y�2�4�ayK-��$�>�'M�B�ew��3���)��g1#q�?_�|��!�"��V����C�QH��SŸ�/�B�8���Gтf9����e��<�����������A�i��y;�[ȕ���TKF7n!�#z����[e�O!n����uMK6��>{��\��g����r����t�����0M�qm;�S�H&nu�U^�C����wT[S�;��V��� ��ɗ�LH�8)�L*�,p}ʺ:'�:�,�r*'�}���(3>3,6J�r?u�[|>�e)A벹�ț�kd�����g~�hI���RZn����@)"�s6�aA�w���)�0���t�Eb%|^�d7ӯW�ϕ�K����SY|DOAY���"�OPvVS��%������c�я�V��3�1��RQ�W��a�fB�瘩�I\�(u�=�XJ*f�6eՒM���w:�B�eZ��̼Wa������6����v�F�aޯχ���OW�AaS�^nmX?�<:��%m.�ޔEE)���a���c���o˟��g\{cdop(e�43�b�p9&yw��^[sv�B�Y����Xr�qHz҈�,�I�{�ξ����!�ክ�U1T0�䔇�R2����!z��7��`��af����k��#��j|�/߼���r�&W@(�?X	j?��`p���T߿���^{������~&�OX�G����>0@���æ��g8"v�+�����7Mn�" ;k��T������	���!�M����Yzo�3h��O���P�p�k��ek����H��y��@�e�����eWU��[��rN�x�¶��
$��!A�N�At��<�NJ��0F��7��]���r�w�N�*VbB��VW�� :  6*S,'��H8��x/�s�;�ŧ�ʣ��ga��fD=�+���pF-��茔��"��	xв	�����B���!�\jq���I˧����~\�u��k��I��پ���*P�@
��}@+��(��V%�Z)� ���/2��t�}��b�GyFկ��:�W���s���u�~L���ambew7�|]e�^{^��{pyq��)~3�}Vu��O
@��Ï?��u3�6a���l��q�j/�?���_����/��PڋS��Iv�v'Nx�	�u� �Ǒ���߽�P޽��̖��~��[VT�r�=	(A�&����(���/��=�]tg�!�4�d�Ӑ2S"F���&\Z?~ИiF���m3���8�A)�h���3��ϣbl.��ϕH[�\M)��y0�a8&�h<�. n�xn�U�2u ��֨&O�Y�Vt�hQKB	MgϘ��V�lr��f�/ޠ)nR��2�M�:�T2�&�ˉ����W4�{,o&X���X��ns�PrZ��mJxqrJ�Up��
��f�8�Z7Պ\W�{m�SC���y@SD9~>�O�^=7g��4�����!/+�R�>CC��D�ppM~z�;�������7���9R�Z��E�Spc�ɀFi�f@R�?Kڍ�Me�M�;�s�˸^J��Y�E22z.	{g�z�0�;��hR=�5֟���46w�����˥=)P�^�0Ĵ��P��l�*����~����y� ��	�q>��G�l�n�6�sQ��`�m�F�fӁ����}y��ܬ�2�?��M��c�m���w��r4�pս�B�K�*��{-]	�H�����s'�)CE	�{)��,T:���GL�&��}E������l�潥�x�,�=6�`���]�v�Z��v$�oG��>����s:�Gk@FB��>��V�g����ѯk�3U�?4'�!ʇ�2��F��rҁ���3��s��`�6�|8�F`g�ZAR߆ �Vvִ�ݳ�83�]C�1⃚v�sa�E��T�`D��4n��4�2?s%����Y*��e7��M*|f���Wh�K? �7���z��xԟʻ��qB�Sn���fC��^e9�q�h:blL4CAhR�ӚA���*���-Az��sO*�l�X����|ٿ'���Q�̂���0�3�i"��pswσ܊dW�Q���$j�'\��g��j*����@O���v���c��_�����y����^�� p��~�l���ՔjY�Y��v���Bb<4��1g��z�k-��x.҂m�h\�f���JVV��[����Y���Ɵ���j{6+ι;D�:�Bd���i�X�g��#��.13���aSO�x%���n��3�4N��m�B�CU��p���=eY�ʒ~�������$6�%�X���`���Y)�l�o;�nrK��i����Ũh6T�nˋ�K��P������}��ά��E�/R�@Vfp���G�geYH/����\B�c���ۋ���3��'>�tT�3J��)���~�6 ��J�_hW:�e�v<��Jz��(?���~i��8:�e�ؐ��t�H�~-c�3�ނ	��#�Hdk����UFw�̚�oY��f\X�ō#/�6��f�9�*B(����Ca��S �	�����)T������UzC���|�����GZ�N�Zsz뱂gX�Z:�;>�s�:���W����G^�o��.D�!Q�r,��j��{������q�xآ�@Ѹ<��Lٷ��C'}a$	M �M���P��:��ڥj��8Y�eChї1�t��3��m���|������ ]��ˈ�e���5_��r҇e��y�97�D�{�ʯS7+�R�8$n����6�'&�gG���K�»e	�)���^Ä���Q� �LE��1�h��Q6;�>�AT���0���Tp9�MxQ�D3�+�[ݶ/���N�2RRg�K,8�b����K����#�C��?��rd�ܯ�l�G�����'�4wv}A�B)�{��N1Jo�N��KS�5��KJ�d5��՟Ε����J���1�����'��a��.h=��@
�&J/i�rsc�b���h� Zj�ou�#���Lg�y���4�7wA�ꎙ����}��Wr� �y���~��O|߸N���(]�h!��y�|��oH��-�8�gP�w��b(����jO$�㾜8�o������	6x�q�q(aR��_�z���ua�04U�S��	"��,�.-�yr ՐSf�O� jrWҝ!����b���]���z���P/;�\>�8�6M5��l��q��<�џ���X�,~�c������Fi<�[�	(3��ɀz>�o?_���N"��\~6�Ɉx�	C�*z#��Z!���/��3Wـ��Aؽ� �B�9��6e;n�C�I�u�x�l�M���\��=�)hҕ�w������X�L,w�m����^S���[�ku8�����.�-[#�LϦ� �\�,�`o��V�-x����`��X���H/�˞�։8��t[n��<Շ�~�ݔk��K�O#)>$���__����%r� ���gϢ�\��ׯ�O}��%;��}t�1G��� ��<���5`��gӴS��T5�Ƶ��\\�usuK�`�9��c%2��u��ր�ۋ���ʂ���6F^7�������"p��U�2=�8����u7��I��zŠ#��j���K�L0{�B+8iy���d�ڝ����0pB�*T�b�$F�}}�taL���ĥS�a��Yk�l��j�ۍ;���}7�6K[�W���� �M����\%�;��җ�ҳ�fP9}��!U�b���	���C���%��3�����vI�r4$��گʌv{!�&��9�Ϸ�8G���w���^�} އG`(��}�����R��#}���9t<n�"���mG��"P��ȱ�<!�DOz��	q�f��<<T�P��*i��N|O�D B����q�~��SD�F�#�5~n䆞����Ԥ��nI}��	�e�4K��V�]�뿣�͉�CYM��@:޲\����=�;�#�]�<���؀�&�s�ݩ|Z_���X�{�#�+Ϟ<-�4+��!#�QI_���01�����oI��D��F�i�M�Ӓ�sm�<p���Ȱc$pf� �#����V�B�<At��3��뿠��
�T37G�e�a�Wql�����J���;8�	��X�t"8X������O�Z�@��Νx������(�}���6{v!�m��^xNf�࣮k�4&�s�G�֞<eՀ�;�`�Y8�LD@�n��נ���S�,0_g�JTO���{
]� �Q����;��t#G�C��{��%;�K�l���+�ge�m���=�v�Ӎ���H���p,�T��p� ��N����~� z�9ԬL�7�#q�le�j	�Y�)n��S�eT��RO$�"\H��9:��C���n)�#��F�3H��x:��x�Y<cÃtN���X�?��%f��{�7��Ԣ"r���fp,�:tB�o�� N|p�DVq8�r�i+�[����T1c�$��;Jm�y�.k37�e���=�C�����rW(��?���h>h:�Tfb }���~Q���"����>��Ȳ�ZK������bW�"����!��DB�}?���|�-E��e� '*�J�i^��� ��ei���x���Dk�
�Ŭ�k �/�t8��C���Kwpc��Ox����.�"��$䝃0K�&}`�}[��)f�'�g��0x���D���d)<�9>��l
�W#!��m��^3dH�a1f~�=���h,:���?d@���+R�zjZD3��k��#��m@^�>�!��p}���>/FbI$��Vs4��,�9���w�>���t��e�Ϊ%͎V�!?���:Mj�Z�hɲ��?>�Vܨ��*:�#g��'��{#���8{��(�v+��#�x镲3ɧ���r{Y��ip(˯�}��өb���[�iU&/�w�$���\�%�P��q1�U��c	������=?3��NQ�ز���|.�1�w��@��J~��\\��33�ȼ7Y��;>3��t#��")��V�_��0]�Y�a��@�,<��0Y������eѧu1�%?J{7�n0B
�e���(�w�-��p� � ��Z7�T�}��3 ��Wgk���8ޭ���7ߕGk;��ײp=8���z�M��Ĭ�Ns���������m(d��'i�6'���s��g�5)�����3��ʏ󫈣+]�2t���p c�ܮ��6�`���2�����e�����q���N�u�~�D��Y��=���I������~=01��E���3 �Pv�(�Az&}ӏo��ϧ����X=i��-��W̊��ɫ5��t�~��qu/0�J�_N�����0{�+�8W��vX��fu�ج��2��5��|��N
�e�}�h�Vg�_�lʥt�Wq#��+E)���.���X���+��ԑV��x�&��'H��$�)��8�-��<k����_Z�')<��7Ew22�>1K,� ���OE0D����3�!�V���?��,W��9�d�\�N�x��K{����\ҶX�+���r>+�-���P��W�*O�~���R�ϺRx8p�j�M9���Y&"P�Hh 0K]����r�0?���+L6�P
b� ��)��8�0��a�1���<D&���r�JE)M���FJ�x�!�"�"���Db�߱	�Te�p��ʺ>J]46�m��%_�M/�/��V�. =�����,?%����:��|��N�l5e�E��,
Cpx�~z[���ӣ��E�N~L*�
�ڇ�2���X�L?S�l�W0ޢ�����J�X�ptC�l���D�k�5��!��
	��&�jk�j5�_��f*Ta��v��kU��5�$�K�� ���ա����#��AZƅ4�Ds:�嶛b!rO��> ��P�@�����xJ�_�fx�F��F �Nx������t��@(?�0�t&��)��L�"l���L#x����>2��w9^	�x��/��2ũ[Q�X����`6��%)b]���� �@�TF�Ξif��:uM�I��u	��K�ސNl��ح4�(�A��Ե� YbV=Z;(s��ofI�s}�����͗l,2���!�l<Ċ$%=�h��?}�Ƃ��q�76�	�pw]4A5��Tf��?�85/z�F.~z�jW?K�v/8@�O��!r�C��o8��Ӷ��4S&n�.)W2xW�"�0�/�X��/(y�5��;>�ӷ��cX�@�p*� ޯ��ǈ����>��]�%s.�c^� �J���J����� ��M�9���.�UL"5�9Y,��[���sò)L���M:���S
�<r�Ջ@*��3� �����%���R�����X�������%˩v���#��4m,��.R��_�ݥ�0́D)%tx�<_X���(ZL���HV6��`��ӧO�b�OI�
1<W��V�@Z}*���|;N��j� i﫡�b%�Ab�k�i��{Q����5T do����g3�jܟs�?7D�<s�U�WD�/X�"'uS�75]߰����
��J��/�L�`�C�h�|�O�E]�z`��֠:-�3 Y��`��ki���e� 2u]隣���ƳJF����^`�Iߑ*�F"�nsM��.�%��-}����j�,�G5�+�IW�L
ƈ���R��~��5�SWt��W��Ϟ���7���X����L�v�]VbY��ەTTG�̤f�C4g���^Jp!������|J�̼�ρό�@e����Xf���W��}0���ۘ�:It�M)�J���ҽjY>�-xY��7�����T�п��\~��bs*��Ɍ�t?3�ӇQV��ܥ�T�G��w�������rt뱩ݍ[�8�"�*�i����io��\�%R4����Yw�W�(b�l<_@hb�/2�F��ZZ��Ȣ�č�f]ko���c����F6��[��XJ�����dKwy���s}S��=��\6�����.�.,���~/'H8!�t⼣���s͒ݑ]e0�肩�k.�a d�o|Ko!d�����Zֿ
*������`G���OL+>e����~l����{7j����
�,�ݷ�G����)�9��%�%6��ᥤ.����2�^�1L� A9l9|��Ff'�"�����L���v��)��(eia�SU���)R}���J���K��VL��!�J����8)��H��j��f�7Q�	��iwAO���m��ƭ�:}��6���{�s1���7x\l<ov��!�g�ߛl�;g`��1���K�Y/N�ǛG�|��jR�u�b�1Es]��M_���������m��dƅχ��5*NXX^��LX4�fA�6Ȕ�*dY҆���ڮ�U��e�N�KK��Ǔd�,ivY|$*�(R��N?嵰�@�.F���@�[GP�� ��rs�D��Y���ƞ�����g���t'x�� {���[Q�~�Gf0����}��0*{�Vo�n��8h�%�U��Uɼ���d��\�n�o�s���a=�&�S��2��ϩ���lb8�&ɩ�]�v��x�o`�!Z)L��- T���3�%�|�09�/k�R~��P,H�頳�_�f:`�T�m�2�x����rv�����Ϻ��E4���,80�H(>~����NR��y�sB�7}$N��#�ָ���@�X=�R4����v��ei�����E�0�F���_�	o�܁#1�i̩'җv
\%��"�Rr7�*����[7֤�NI��8�Yj�<J���/a2��bx7F�$�[�i�vV������ä˛�]J����/y�T�:�<7@7���k@'�1"Ld����pee��l߁�N�L� MkR]4g�oAi3O~Y	+X��%:��LF��pB�U���L����c��)~��pPM� `��E�㚁�;�;�Q����pH7�MDt/h^�s⥋^��%��z�a���f.��"���|`�]m0i,4���`�HmG������>Xsh�aW��*�;l������}��S@��tnR ��+�J�X�H%�#)�A)~}+�kh�b����������'1�]&=�ׁ�"�i��My���#�}V�����-a*Q��Y�89�b8��A6Ⱦ�	��'�H���KC��Q�
X��h*����s��/E�ei#q��=�r��m�ƛ�%�˺:ƣ
�7W�\w��鐚�xFs�\o�\0NR��Y���i�ޝ�:fS-��l��X��^��V�y�0s<6"тZ�ϖ��p��A��8%��
V�W�,��rf����5������U��R�@��SH,��.���sN�.%H�$���/�@�� �/h5�f��XXeL[4)f5�B�w#H%���9�N�#~�?�� ���v��0C	�����FV�����?���Ebm|�y��xFjtL��vM	����½�Gy�r��_-,0��Ti��K���?�JŽ�3ŊG��I�.��<��mGضD5�go$��~���19�Gf��{a��������zj�j���>����ә�k�j�n���@�ဓ�6[�����Wt�#��sy�KWߚA�{k��zԡ�
��:���T�pQ�"��uwY�7Yͻ�w���q��?�ڷ�����C���ҽi2�������� 9/�������^�uQy�R<	��%&b斋�+��){��м/2�e��½�W�]=����'~L%�9ic���=��),R�I�Z6㳗R�	}]� �@���b��q��7:րK��3�C|����j�@G��7���Z ���8����:ʢ#ӈ�0D,�~����FY��E��x��������C���x�,��G�n�������o&y��`s+#`���9�q�T�ɚ����_|Ů�N|0[�����y�����j�2���#�8T랛u����ǝ���Yf�%.`̡����c^��9�_?HD���N�pә�!���U���L� (&A����6|���<�f^o[��/1�Y1�3�l��.����;0��fh?4��*���}#ڵ��B]���\,����ӟ���i�I����}�iz�����G/)S�y���:�`N"�k,�"1q`��>��^����w{t�'��)ˇ�t���υL�,<\o��Y�0FC�n�����Ɇ�'���6��|xS��¬c��Xi��ʂ��v�� �ˇݧ2cl�ѩ�FP�Z*�����A����Ä�Ⱦ����+�1���,�Q���gg��ٽ��������i��x:V�� {lP��FA���d(�ݶ�Y�ǉ�41��������ݭ�ҹ9�fw�V�uo��뺚�}%ㇿ�Pǃ6�(��o�a<��բf��T�|w�'��ѐ���(�%�|ntؑ�o�����t4�qa�:�{�q�`�	er�7�CY9�qAl6&����i�{�P*�kzT%F�|%vF6l�'Ա�)�}H��m(��:���ji�rM]�\�P��|w��n�dW�m��0����݌t�L�(���&pȋ���)fW�{H��!����(E1��(�Gԃ��˅�����ٺ^/T��Am�~F�zv�Ǹ�8y��g��N�C(�/��:e����e �����j:�s� w�(��H�E��f|A��z,��٢������׻�x�3���]W��J��`9��:G4ů"�I�������ẩG��_K��u��Z	�Ӂ��m���ch��psh�˃�">-�cn�v�xx��nF�����h=]i�K{}��k�]Rg|�JH\k&���ذndCI5#]�ac��3��z���#)��A���*^;�붼-�^.1���D(��R0�{�B�\W�!U�<���2�SN٘��:�P	t@��>���x�����"�NM �X�H�(�:35��"�Ɋ������H/������g}�K�@0&�u�oxv�7IY�9Z/�^Y�U}����E��73��-)�r�^��'�RqQ����o_�����).�qӒ�>�"�R�wu�jiJ1e��-)XL�
����,�l�&Y6d0�$e6M�������L��q��z����b,M&����Y�#�+�J`\s�ŚL�A�ڮ(-&ޑ>��b�$"{��!�s"�'�a��sp1nz��Ō��S[�"]������]]tf���Q!�G��oK��?c���R�`'��qH8@�����VD�w]�Z��
%��p���0���	f:��H��h(�)��<th�&fH˕�63�C>��@�~�$T	��+�S@��xh�U�Y�RG�ƙ8�<�����I�nQ�����3���x��-��h׃��)o�gM~�J��T�JR��[��'�m�!?p[�%F)L)�e��(0��}�]�	��D&�Ũ|��P�S'm?�^�W'lƜ�>�V&l|]-����˧�F�� Z��(�2%�/��أAv[/�)����4v)R�?�2�s{T{��M�Z��F��W��q�ċ{P����e��!�����m�[m�ϽdV�4�*��3�"�7��e*4W�ጃ�or�D|�f���x�@�MpD��q�0|s���pY�}��^_�	&齎����� �z��������J�pă�Y�r~�+�w*��|�Ek�辎]�߼���Myj���FW��)i(��4]b�5����$�������Iy��%����p��նߡ��ʲ�*U��O(����P����x����͢M&B�P��CǮ�SRZ����A������t�M�K��G��.*'hc�@�Sj�,�$c*\s�"���f�S����X��Z�+�)]s���%S�o&�/�.�G܂�4&���L��V�q��FsF�`�ٷ���R"�s�b\?7�6��i͋s���@�f�,�&x·;�x//��d �葴��xt|ޥ�ƌ�� ��x�8I+�5�-�ğiC!��<�ys.��dш�4�F6�]-9�βvA��.3>��R3�6�a$�s�g�u�������,?��M���D�~�i6b�U���0.�������x;Ѿd܅HI,�6���"��<�$p��Hn6����N��7E��z�u�j�.�1��0�w�dY�8n2@���z%@h\K�Շ���
���I匠5P�e��g/J�"Ll���a���7,�}a��C�r��n�B� ����Z�Y���x�]������^������aF�5ծ/<�ߣC��ɼ&�f쏎�jO�I�����:Y�r�L�"��soO�) �-
��
�E�>��cC��C�����ư��,u�8�Z�'<<��Y{P{VՑξ�r��E�7k՛ ���vsw��u �`H�yM7���Bo�>W>$<O.��Hh&�z8���{�~}��F �vD2�(M(�񳽰�R4�����w�����l�l��/�L����\E-�ک��㸡��E&�s)�SK��C!OЬ�����?�KQs�	��`��K����v�y�K����d����g�k9�o�Ȣ����A����l�\�Ϛ��s�9	8׊�9З��Ǵ�����l��i�U��X��'C���,�zǤ:���}�>�I|��x}Oi����O�r�?k�!
���)X��d��d�_������?��P�k�4�"�/ƿ�e����f����InvL�xw1�)��]t�z���̇d�s����S�=�0��=�� ��P�W���t�i�V���@0 o��cq�wblT�֙b���s��o�Z��� ��=�������E?�( M7�m?R�U{���f���bi�������F��$��0�{��e)"�sl����^�/�q�� kl*��μ��6Z�1�Y+6�I�O^�,����7�'��%�gF�$��T��'�ܪ�i�
e(�s-e�e�?߈�WЫ�i�#����Rjf
�^-T�ϩS�E��6�k3c7?�)�C�)�" k����[B,{n&s�	8��-�)X�2��s -��-.�ES�Ą�"�js���գ1���G��C����QQ/4x�K�B7(�[�s�:��d��`˩�7�g�l��=��4q���kɿ+�I#�����
�G�|6����/� ����e��<�e��[/�A`OQ�ܮ��xw�cҦ=�Qچ�׎�����f�T}����l�1�K���_���tNH��;��eG|;]��W�t+ ����	��l�Gp	#@�z���R�Ė�\�-ϳ������8Z��g���7�b�?�����_S��/�s��?�'3�5��=��T�<r��?�*����� ��Ȉ ���+OETn�I�͇�~�ČX�(�pT�M�2�9G'���r3�+�Ģ=�LTY�V��6�K@H}4@bp���W���﻽ֱF��['*�A�R�֯�1����Xa�Ҏ$�O��D�l\M���(�⳺�aU�5;ż�1�,?�k��ס��>����Fj�"��Pt���ף�����ۗ�O�gO����H����81r�Ղ,���I�g�6��Hy�Ͽd�P-Ӄ"	U�asHƌ;��oERC#J�턹ڊ[�B$�(�Ej��c?t�6��3��Ҁ->(�z��TJ�ҙ+h��|�b![6���R�ڃ`o�A�%F0��r =q�m��%�f�w^ڋ������;��}�(����X�q�#��9>)C|��� �a����2��t7ۮ��{O6C( Ŵҍ�E���|���,��d��o^��Pb!�~���E��̌6���4�����i�C'�R�$_.2㺾�fe��䭙3�ߎ�[����ķ�׃�2�a�Pc��l�y�~[|u��mr�l� o#�*>�fJ���ǡ&���+��H��7sӐy�SU?���� ��_�Z��\ͥ]J��]r��lW�'���3CW��a���Θg���~��L~��fR���G�Ž��2v������e-�R| �{���x�r=��,��x��}LHTRk�hw��׌t�r�v�b1����A�U�7@��A�C��]��R����e��ץ���X��e@m����=������fiTq������9���6j�8����8L�"#���6:`U�3:���Qdx�?*����JL�|�K%BPY3B3��oN����	����u"f����5]��`pާ����[�����-�X<��kg��n�w%@���Mr�
�P����o��M
ŘF�A�'q�.�b�O�ţW��ͬ�̹U2�ŧ�?�RN�(�f"���	H u�J�0���2נ�X��&MVw� yE�Kh��x���d6���W�Rh�y�[@k��$H&�AP�RY�e�"S���e�.�� sB��y��n�Kh��f���6L�K.��RrM����hvjn-uM��.�����P��Jw�j�Ce���i�WS��Qq����}v��ɭQw%TK��RU������{⊪r�}M6����<���a�dm�?X���6����}�G�����Mr�RSr��_����Գ�0k�%�����W�����1��p� �7E��MC�Y"N=�*�$�"�P�A��S���]�c��TJb^��K��$p�w ��w�6Մ�"��5�V���rgxި"��2GwH�n@!���g��W�)d�=E��ГlDy��C�N4�J��!Y$��Q�iߧf=uj�z�e�ػ(`G	W�����PޜQs�k��z�� 
˗Ǵ#~Q^�q_{����3�QӅ���Kh��&�藥�q6�$aL���=���=z�-�&+Ö.jTk��zY�(�LjH��KXc)9�P�e��>�+u��v�'�,����%��0	�5s静�U��o��_q�庾�s���|��XeR��(?^�Pi��]I�a�1IB�;)������xy[vc]�1K�y~x�jI_~$�� �f��/�{<��/�9�Wf1'�K�j�y�1��肋d[��t�B�{/1�#����YZ	:X�3����44��#��	C��w���H��_�L5�j�}�Q�$uC �&'�.=g<Z�i��PY����m�M���iOb�3GެMx�[��/�iRFj��z"��� h�p�r��)�$���G��S`���*�&��KB��jHuu���~$o2��R5�.�B��k��ur��FLh[�W�1��/<�|�g����^4�����T��QK�_A�����\@������?wW�Ǽ�;I�����n��5�O��� +^�%��&�ٝs=�4�P�GC�o�~��t�:����.�ڰe�_�Di"�	��㭇T�H�Z���� ����֦b���L����چ��[qoG��א�a�������H|�,i�y�%05�����P� Z�}�������������=��5�zE�R����.j��W�	r���Sv+�,,ؾ�K�0�)J�6�Y1�g��s�U�N\\L</�7 7'�p�/�do�z"�J�{�F�bX�M��m!��B�,��+�*2��!R۴y�ʑ��!�	(��\2��Z��7�7y��[��t����.��u��zu���e����Y�5���t���}P�z����E!���q�^KIg�x��ۆ����R��qΛ�͗�&_藯������">�
4>��`լ6�֑Uʫ�k?ls,�B ��a5!�����B`=��j ��E�OҼl���bZlϧ\�Y�u:ͱG&Z�Q�_�fVe@���/������0	(�pX�\�7M�b$��>WȍY���x���������7��U'w�P������ԜS6�����I�G��� :�������ǯj6��d�X��s���;�"�ؿ�4��r��E��1�� 	*�;�T:?��xHC�z�#8��˂&�/����٠���|�#ٞ�91�^5Q�EI�Ʃ��O���X0�v��.*���\ov���^�$>?0+����q�z�\���kb���F�K	6��ȠBQ��Y���i�1����"��Y!���ZT��_ڲ��;��ݠ�i��X�ᘪ��ә�����{U�s�싗�_@�	�>O������5����Q�.�0���{�Jpo!2�3����]bddඓA��$hhn���
�M�*5�-� ��{͈[����.�<���{���vQ��jX�K�6!��\{�q����K���z �y�1Qd���XkN<ܔ��o�-.��c��o5�o�v����-���d�qȇ��?�^jV�}0n�pof�d�SV$�v�5�֘�K���Jk�?�2����r/�����C
{0���EeH��_zG�Mz�lR�"�Cp�B�'���u3w53�����������@�]�ӟ�ěg�FS�p��ͼ���ہ�^���P>�|�){f��7%Et��}����чz�V��6�zA���)�3Kah=?��EB!
B6��QXw�f &M,��{ ��1�c��ٓNMT�h�k��YN�%�Q�P0�\���.��MQ����I�J����UvG�]bh��L�R����]��_k �������D��`�j�m�-󒽯R>oq�
l���������	�o��V��9���=HHĺ
�F��Y:���?��8P	Xʰb~�Y�wK�����9v��F����߮���+��l����'z����O�\~�O�Ĭԙj\���� ��ӄ۝���%��	���I����D �3�듧����ʱ�@���EV�2>i�OQ}���򾹖�&k�R?H�k�+՟��T$a��p!�l�l�s��7
KK=/�a�x	��c�<�Ouk�UOl��YNn'K�'�Px- ���@����[�w����������Hy�:T�)ӵ^|���A��A��׍_s~fbŚ��k�S��N٭G[Ķ�w̎�9��w�����@u^<�k���a#%�ི�<��`2�6早A��.U�1�o��7>g��C�W�'�(3�P��YN�`S�����ט�u]�}���rkQ:�[�������w�����|�W�Z)^�y;}x�1f�u?����:��}��+>�RO����x����r������n���E�"�7)��l�\�E�#P�yI����Qohc�}������HKv��%˾T2;$�������S�������������Ì����;�/���۲Y��ڳ�1$݄�O� ���R����O�~���8��εT��+�p��~���w�0uR���������Qyk�.��F�M[&�=w��bJD��8^�Cה<��.�����W� ��b��cu�n߀�>�k���a���f�s!h@n �8

/%O?�@��E�h��g�4{
N�{�pm��(62��FR��P�x��C�'�$�.U�,[4�{k&No�O�dĥI����M����9QvִJ�c��`�ts�Z��`�K�.���_f��X,yYJ��K��u�bė��E���׿�*��.6���L	8� �CO����oT�\b��v��5�89Ŵ@c�b�	2d��F��)�T�G�h遒�N��>��PL�La{b��V�.:�`JXw�SESfO.㗸�pNW#�	�o��Ω]�ϥ��,V!лHܓ���̏W`=����U�н� ��P�0>������I�Cd]��������+M��������'i�-�\WX�#���O��j/!�3K!���n���ϺJ���6���F��|Ef'%��$7Cq?�{��F�6� A���iez�8(}NJ�'��gvIw�G�]�L�&%�.2�?mo�I���/� ���z!�x��_5<w�4�]��b�e\TD�,�ȪjNTG	"�mQSE�O�T�7�`;��ـR��7j������j���A[�|��&�y9ǆ�[h#8��
�u�r"W�+�ԃĽ2�2U���>ȳ����}=�jü0)h���61�&,�8e����O0$'��8!*3�'3�[�Uv��
�]s���b�EriyHu#=��^'!�ԝy��8��Gg����UD���m����Q�D2��*��Z��;�zx�⨮��=�h�(��Ś���1���$V*}��û{����}���R~ݼ(����yph����\�>����zKM�YE��<P�^�Z�6�I-7G�SH��7)
�Ա���zA�0g�?���q@@k7�_�(OR�?<��#�2|N$���6��o�K�=-���>��3)e�(�����"��a�`�!�������z��E���jD�(v]׬�z���q-啷z͈�ħ���3D�/�5��A�yZ\c���E;�M�8��K�8mH��`b(��z�K��ZkVY�OC���!�mum�+�M�/�e��dԞ,aH�ȷ�O�֚e�ˠ_=��������B�|��ݷLp����'E�(���eG ,"CSt��?�Ʌ4�1��T�&}�6879C��.���.��n���g���(Ȑ�ȁ�X���&i,���	Z���E2��	{�Hx�ۿ�[<߽}�̑ɳ�S�ȱ�7X�v��oƴ��n����q��B[�P9���%BWxP�x@2�!*x�ž 0�0�����]# %����Uf����\�������{������\�����=p�?�h �ID�����ޮ�5���,�	Ӌ�/�	�N8�xў���lQs��	#ڍL�Xs�0K��%����#Hk	�e6��@�g��++l�HF�"7,�v9�R!���c�s|�@�k&O�Ѫ���c���W뫏<9�7�����=���6��8�&���
RE*�i�zu��.�#VG���kz��ì]B	��?`V.�[�kҌ`TVe��w���|=�������F��)���*��c"�"��혛�L/�7JgjR����W��(@�0<3�󪊐�j��	'<0&ͯ�3T�橘i%�nn�����O[��G�'}$Ԧ�(Qon�QA,����>=��������?G_{�e�p��x�7n���R��3e���m��;o����n�-Op�(zb?*�-��QP���ܟB�@Q3�z�Qڹ����iQbL|��4�!I����m����B���<�dތ��cDp0:��i@��yWx���"��^d�̍`��ߚ�[k�<�1=�N��sx�OOSޝ3��ws�1��A�Ar��*jO$9��'�fTW��	�*����K\9�b�-��}���f���mQW��sܸ1����i��ά��NL�*|�
xL�xe���(�߮���iG^����E�<������m����Z�xɅ������"af�K�i?̙�k��"˫�G�5�{+�!�#I�=KD�e��'z9��R�A�~���#*���=�^9���E/p�pR�A��v���"t�BP~�6��Y>��"w�ǁ�]$�@������OT�T�2dYfx�-�x|Ц9���C�J�7�Զ�~�r
�&�}ǚu�+G�7x?:� 9�#
�1�u!l�^��BB"n�R~���x�����TQ54���RP�� O�O�K`��p]���h?D��rS��&�8�^ρ���>�1\/n�MVɵ�Re�'�׹��p}d���k�\�z�����+L���%��ѮG���E	w����!j�Ѭ{�]i#��<.���n�P�${:d�����9(�"�W���>̎h�?j,��R��A�ˊ2�ڨ�JL��!��C5�1�>�z��o!*j�1�E���t�rÆX,�����o��S����=���c�c�ӠT������y���d8���yֆ���Au�%9��m�f��e�E�U��D�p���˯gb��?�����-�g55õ�UPۢ<���4����}
�)�N�]�C~n�Q`\?eS�gqlkE1�h*��S��')WK�k()&�A��;��'�C�����N�K�C�7�Q�U�ȵ	�5CR��L�7����ً}�1��:�ⓖ��xf���6�Y/��x�?{X�\4wKz�ħ�0��������$�d����/��ϒ�[��>U�iP��)�����!��B���z.��k���,�0	�a���׷�ފ��69�xZE?`6Q�Q��q��t�!����:3u1֏�\
Έ��H�bͣ"h�h	I�4k9��5�ǔΐ���I/{�x�gS]�y���I�J�i����kR��;X��h!;tl��Oo��FI�R11��6 NR�k�7��>�}�M���ℵz�>4?O9�'-��Zz�le�0N�M�m&g����mdʿ��`�B9�׊m-�gQk_�Ǜ��.iSx�өSGMʶ��-�#�Kf9�NN`�����R�[l2�T���>tJ�c$h����aO�X��-�=6�?B��g��R��s0�d2 �d}�� �7�)���a}/o��UΐF��ǨLB5������0���X���f2&�XŴ��;2�
Akr��H��Xn�JHd�����T~�	��{7����K��
FQH��x���ah%�����������_��M��s�߮�*��"]���z�&W����\�;�Cy �x��R����ٌ��oj��	�[F(ƔMK3��a��ʮ��#�>);%���£�OQK��k�vI��(\�C���EB�d)×��/��և폺�ѫY�{S�-#J�emz5uiYjwŖ���n��b:Q�%�G)�܋�'aP��\��H[9TUt��Xk�wc%�/�Q��{�!� �:���2�� XA�������x�E��}����e��͢jc�|gZK���׽���u�l��~���%�C͎z\�T��e;vm����:��Ld�! �=O�?�qaCpw��?n)�Z�e�����k���|���w�m�w�ަ�v$8�
-��<5:����.�bPo�11HB*��%'�/.뜧{q�Nso?��?�R��(c���^���5����
,�������q9*��������"�,Dh�2��L�\���� �bb@ۼ��F��1�pG񮭐�ŵ."�E���"ٷ�s��-�6���v����jq�)Y;�<���Y*�����(�Bh
{�*�e��l+y��\r�ԫ�k�I��E�[��� �?)+�eD}aj����T�N!]�B��M/E=\ƅ��#���.A�M ��ĺ�Z|�1m�R
���P�{��O"�d�;%"��a���q���:�NX\%<����JQ�#z�bِ^�ɴښ9���Qn,3�~?�=���6����W�'�ɈgQFކ�uah$��{������%�~�)��_?�Z>��!<�i������˧���:�sM�Z��*y�=G��hG�����W�ӄr����\e��$"��혌�LT�	@�M�����4j��wX7q���7t���Ȥ�.�S!1c��k~�h�����<( >!�yē��G�)qx't��l�Qಚ��zd5>��c���mXp����a�<*��Ȭz�l��몽��=���6�N����~`�0x�F��	�d��q�Nb	$���W-*3���Ȑj�&������ژ:�o1ӱ}۴���AB2i��B0<.)3="��qdI��=�m.���$E�/�Ԗ&�[�����ROB�ά�T��e�&�
(�
��8��v���I� ���̶�-])�{��!������W�S��]����Rn��E�7L���U��'6'4Bipugz�V��\t�(��,b�d"��IN"�$���&5� ]����~���X|��������Lr���,2�d����+5S��fm�;�D)�(E���G�g�Ͷ�{ml��3J����M��Ya�uY�y����"���?o����#m�*���Ak3G%��t8t�}�jg�����Ϗ�Tߤw�;2;N�#��QG/Z�lS���17��0�!D������D�E1n���E�#���`�y 
�S	F}Ɲ��&s�d>/<v�H�[�zR6�aC�
2�LC
.��(����k���@X�7�a|����j�����,-�l"�I'�����t����T����"~6u��D��DAG��N�}�E_M˼#�@b�O��kL�k�[j��|Ԓ�)X���S�ӧ�"�xd�`�э�Ԙ��[)�W���ј)NL,��ԉ�
k������	^V�
��VI�^Vh��>�J�P5�������%==�'$|f�<��&�a��&����Cy���HX�d��E�r��&�k����!��I�����fyP�A��W,^<²ޗG�a2�f�6Dv��v{�җJU�|��.Z������]����'|ӜԮ�֡�v&��aJ�C���4J��]���w�b~�Ys�7ôa�>s�+B�r�C�!!#B	��K���Ab�8�^��| 邎���^�����a�I`��Ebz��VFs�Q���q�

�~���e끺'� ���{>�/�&Ы!���[i�Z^�9�������7)�+����9L��d��og�M=��i������Sm�O�������cf
1!� �{�p��ކ���}̺�,��$o�0o]3Q�G��[z8Q�&�ױW\Ų��@��Ȇ>�G����Z�c�^��Q�Br��&1�5�4�
V4&Ɯ�y��G,�Q^&�i5�2���_��~�	�Z=��ez��oi��ab����[�X�6�	���WxE(I�m���Q�����*{, h�F�	����`��gb뚘�a�[���Qdь8Xg����)ֆ#+^[�&�Z��b^��h��3��"�JzIg�圴�p��91֪�d!?<��nY�`i�vngUka���ݻĝ	��
����ib���v�k#S�Q"v`>Je?q��jW-�}�|4��`�����n9�X���o��/<�W�,,�W��ݞ�_ϒ���â���D� ������8�Ǘ�U�]χms'���������:�+<&���u�L�EYHf��#%�o��|��e�u5���*81�R��;c�Zf�:�9�JtL�F��^ҧ�G��(��<�j���ť�"��X�_r��{���� `,wҋ����ʹ��JV��!�j�;x��5�L�!�������:���5�C-�ͬ�e��n��<Ϭp��da 3�!�?�yb����o��p�5���)����=m�(�-)���:����wU�5x��II�d���V'eҫ�^?���b,:�E�2�W[~�~ %ѫ=���^���z��yU~zMH�1�O�(<�������/ϟ�>���z�G�Le�Em�.<WT0R*s�<öם�c>⒙y*�Y�tI��[�
�^����~ȉÊ��뻵g����y����ᑚG����;�4~"�Ag�c�l�����y&��v�E���0���Pi�֎��w�YH��7I���x���X�P�1HnB~W�!`�^�R��ݫ���i��K3�u��׈]"����ۤ�Pݦġ2b�a5�����BW��N<p�?3��x��)��)2�Ƴ�Ӧ��k��ш��k�!Y����4έ�=��KG����@�˗�Klfױc��H�2�e8�̂��
в�G�1P� ��p�X"�ޏ!��!y|�)Y#��^ۺأ�G4gb
���x�/�x�F��ſ�3��>�䫲�N6Y�&���ʎ�|E���ݺ0Չ�h���x�Q��ڮ/����9A^�x�j[���}FyW)-9w�������,J��m07ܱ�{�^�.� �p�w�6I��i F|fW�*�>�Z\��O�B�-=�i��@�cmC���o%ӿ2{�-c��C���_v/��{�*�)����H��O�R��������]:M*�޼mS����&�N~���>>�W��)y��5�����{���+����x���k�12(o���Km����i�cc�ZLY��(Q�Z�$t'y<>�=Fؿ��q�삃$�+2�rk3W�dc�	�~��<���]�γSɡK����G2 ���j[��8����'b��Z��aO��&e�̆L<x�9	�̼aDoS*&�*��z|���;���s�n��Ѕ��T!������5�BO������W֛M�0��U��r\�`�Dx8%�va"�Љ�mZ5*hD�rƶߒ�wz�<]�)����c��<�'�K�+F��G� >Q`��R��Wӯ愼�w��n�c9eY+�(k�On��\#Q����č�R崔�kjN?��̥1t��j�Ք�������UV��ǩN�=�j�ǈ���}-Z��IQ��jT��D(2�w�G�{�����>0jبT�~L`�2iQ�x�ݝҝN�I�R����83_�+��s�$�/���d�"�Q/�6Lh�k���&x;Ӈ0ː�ENچz�������]y�=��a��nw.��R�dR��:W�}n�k
Y����~�B��ɼ^��Qs��
�8�)�,�գ�]z�yq8�E�u75�x����I��14lM��M��݇d���%Ń��#%x�R�][���)����׻z���@C������ol�Ñ"`t>|�D����A�l�Y�rK��9��0u�@0Tz����֬��k�S��e`��\\��^��|,mG;�CĤ#�s�,�n�E����d��Q�
�cL�1����YQ̤��l:R�w����eqB��3Y*m�;�K����珄����k�h2�%tׇ����n��m������G����G_y���Y��G��)�f_�6TN]/�?K��[����bj��nZd���|�}�T��΋j�q=Q��t8�b�!��}'�;C�P0��L'��Τ�X�I8S�}X��I l
2�*xTT��Z��S����Fx�P
�u�����/�h8Yf�;g�G�VowƟ�2C�e�,�Zz�����r
��":KW�R�v��92#���J�L�g̗���zT�kd��,����+��	0n
{p� )�Z��WjѪ��&���0�X�(�W��Ȥ�47���S}�u揊T:�B��{2xs����k�Eob�و��Sf�}P1fv�!��N�C��Ug���t���l�kWⳉ�>dN!<�K��I{+�-�ٶ/�����dkp���f(J���c8<x�u�褻͕އ��{�������O�&	�k������潞���-]~�Y0�w�n��NL����s�аZo��G����x���Uǵ���N<��Fԛ�,pВ� c��ߑ�9[1�Z�1^6.��7����Z�o����N�9�Bwr���,w�I�i֋��8�o6�s)fR��5��9x1�K��U���:���hh�Q���w��d�t��Р,)t�W���%m�ȕsx��L���1��{4'�Z�^ -\����
k�h/��;oLE��\v{e�;U�]Û��=���<�s�.��
��K�H6��@2n�W���ȺB�z!��8��$���s��Z�\��T�Jq	F�J�5&�u��*f�CiJ4�ue��2UF	���q}XnM�J��o���F���>j�qS���P��=��'�֩�hO�u�]�(Gđ['�7{����O}�����*�Y�@�w]3�A��C<�2��Q�0��N'
��`���E��볔��z�u�+[ZR����{��k��H���wlh�I��z���MS
��w		aYϏ�\���%�#��ɚe�˦�[����"#7q�\�����n����xK��$��&��1^z�6q�ߤi9��n�ߡ�������]Vz�;���|����"n����_��c�a4q +Ku)��V�R��^_����	xl�� �Ql�P��fa��-����u��DVR����7�%��󙸠[������}�Sg��`�өꑶP��Hz�Xl�OO���Cr>�dG���\c��w���~|�>K�C��O��AD�%�+�z^g�w�!�$���n����p��Ѕ��xf���� N ��d�n��\0��̈��ez���)��L�^h��M)����.�#�r�!>)��}�U=�5Ƕ�Qц����^��R4��L�fٰp�P��B�
� �ްn'^7����5��ZArܩ;��[t'��{��B�t?�~4Y{z��i��?�遼I�8�Z�*]�D��(�v�l��L>��3�|���H*U���F�7N~�7v�q�S��-r]��I$n���]/�u�Ԉ>�8�b�z��ZQ�����u�ſ���،e%1��OT�Y���o2�F��(� `����,���+��fu�k������$r�B��-4+�l�U����m���)X�1>�l���Ñt6��L2t29�p�5ؤ�`��:�C��+"�|WR�r���Y0�Oj��+��^�gׁ��5��G�:����/�5	mg܅��nB���k�	BW�'[;�Z�%���aT)8�%���CtDާ�zSrK�b��cqM}`�9�u-�*MM|&�:�1�"������d���f�5��ض�r�ї+���[kFGZ�1Bx�B�l�1�ƴ}��e�?�+�ݰ^ؕ��1x�Hy�i������O� wK^ߡ�D_�/"4�!��s�r2��ٕ7I=N���d���R,8z��KI;��=4]�B%��9���H�J�~~��?�!56灲�C9cw�*4�!�N�%¬��Ha<@�\�g�_�Z����O���}�q��q��-��T�Z�*�<��ŐE`v{�nݕ���d��GW����oW��*хaǵ�N�;�p�\�f3��s5��!���q�7�cˉ!����>��ck�DhB�K��w�
�FDr|J��j���8D�od�Q6����	�$_D-=-R(X=���w22���=R�=��k��Z_�*O����G���6��L��	 ����ct:��:�iCp���dI��������\�f�3�c�l��>VA|�W�6<�V��PF8M��8�NVwǲq�6��v�g�M�[+VK���U���3��׼�H�{џ��5������l������X�d���2���h
ňutQW�_�X���B{~�'�9�m����QM�0�nl7���*�	͞x�s��=Y���Wx��=��F�+3Z�����3�T̼�u�!��13c�	o�F-]������bv{ge�c������s:�j٩7�M�:���p+��5 xh���X5 �^;���3Zqǫ�#
9{ܢ
Q���
R�<F�da��,��:��b�c����y@�w�z�a�&�6$�B���1 $pm�&_�Z��x��L���T� o��來zXW+�$�R+��Ą�����Ze��v]��rqǬr[��YK�3���"�7�`��Ե�5�u��B�a$M{�M�<��ͷ�5�w�h��:)�4]�D���ee��	�r�q3lsa�+>��d;a�.��:aGx����ڿn�~��F��hL͡=]��ucm�Rn"r �r�]�'N�u͌�=��8�bK2��@�{s5�"���,*[]���`ׅ�r�4`«m�Ko"1C=[�2�.��[r6��{�x<.�K�U�LЖ�J�̍��Rd��z��#3�cq)Z��\1�/�X�7���b�vB8&6�^��>�Fӱ�9Wя|`P������PnaL� *�0o��o�m���c���툟�����(�m<��&L�	þ���w\c��V�����K�y:�<�m5�1���+���A���Xc�i�eС�u�҃���%�ǣ��$�*�`��~�f(�#�C�/�^�D1���S�0�3� �}� m�����@�f�^����A0��SJh4�iY:&�n�9���
/퇤�Y�e���%��tT�2�svy`�.��c�дb$��>_w	��tb'�7��h^#�EzB���|�-�r����1�֘�ޣ�OR�n�D���)��K�"B'�v!ls�ݓ�u4���d�)V�V�ǣB:z��/c	�5+)���g��x��V�@�f�>K�܀m+�֐��[I=T鄁T����ϟ�|��
��\ϻ�މ^�&��Ã=�v1N�uw�*LbB�k�/�E^S'��2@�q��1(07��%=�ݰ�:��>X��.�8�U-�C��s�AJ"�{�X�p�6��� m�|����K-gb��a��m&t�J��)m�W�\��8%���zz��r����nRo��q�"*עT�ˈ馌9z�S�y;8�8<�Y�йr)�{�[n|̽�#�ab�b�8�M��eU�A�M�'\�����ņ���2�w��U�آ�9+��aD�.EP�X	��:;	�~�1�/���)<��k0_'���}�2�Z�������K�����)�������kCK��C��c�U+��ޥ>�׆��7Fj#J���M����f6t���"�T�t�˭�tux/�t���	Ց�_�������λ��&MBySuc�y]kے�:q��m �E��6=^��d������τ�j<�nL�bh��H�
�����<�����}C�G2�)�L�|����đ���9t���.�"I8�C����&���I�ɋ�`�X�=�RJ2�5��3�a�>�;0�e��U>���p�mS�	5�1���XZ.�4�ʈ�pO��1��d+���^s�m�'�&y�ز���H����Ty�Jp1�C�����)��� zܱ��P����t&�3�>��֔XeD|:|ݔ���J�RP��8V&D3�##�z�mX�rUm9�Ϝ��1-EI�1�C����X���%yG.H�� ���{�nWn���e��/����ׇ�A���Q��S�{����;�tr[��+�NYԨX�H��>�M?��o{��	�P���� ���ڠЋA]�4���g0�_[¿E+z颶C7jb�7���*'��� �������٥�������Y�#B�i��'O�|��M�V3�i���*(3!�2k}�)\m�K�lk[�G�!)�M}S��(5Nc��i]lC2�������&��W�^���;����&�	<E>��:��T��A�*����l5b�B�l�:�W7�1��"3A๥�u����l<�O2���І����+7����Ĉ�u���5�-�=-�A:��.!��u�(�cn��.�\1mؤq�F�q���Rfr�6AE��-��t*Y�iМ��l�+l6�v2\��[�q� iNzԗ-�{_�u~���Z*>[]�5a�4i�5n�Q�\~e�hWjh��¿xdh_�/Z����P	��/Ɖ�#���R�w��Ӓ��b�1Ɉ��a�
�p�l��8����9!�9��>�:�c��C1ׯ]���`gʚ��"��;0��x�;$W�tR�y�4�Q$w���t9}�@���ٕ�߰jf�k�g�a��#���^��_>[��F���lx����`��2��g�ۇ�U��*����c=Y�0=�^	9�.=ĈPJU������®�w)�։��怄ln!\�)3�V-r2��\+N�:��P$�;AY�JFg�M��S��x�����18�ı�$�����ɪ d�8 eD�0|gaB��yT�I��e{?��_�����=�"6a��\���+����}|0���t,'�S�~�/Qe�m���]�۪[sבa�~dr���O��<r߽�Ȳ�>�� �`����}��2�mDkh���~I7}�B�Q�ԯ���ͣԤXM�6j�M�i� r1f�p�hL��!C�IŃ�����
�����V{p����
��3ؔGi�><̹��� ����IB��x�I�o��#X����0Jx�7����'�:K?�B;�j��A�g;�)�F��������ϰ�'Iz3����}@�4�����׿�t�{I��񟳫Q�y��,�䂱J����Ԙ�RwT�f�rOob��QX�N%�U{@�`����<`�]I��2�N><nj��|ΤM�cF�'k�5�[;q;fRe��f{|��I ����n����������*���ڳc��q�h5}b馻Q��6G,a��p6�Pu�������ݓ^�Ο����t0XCI�q�=��1+��:M*{�2~���F1_��tU��]��x -�3�B������/�#ǁ�1���_��/�E ��B�z[���P� }��4�M0��M� �k� 3ac#˥E�P*]Ĉ�2��y����+-�fw�9����KՆ��*^�K}"8�!�P�l��
��K��06�7��TA]��|�kÑ ����	��)�[��}��l���76�ZR������ܘl��x-�����#C�6<Ѩ�>oF�֫gn�A)�zCu�r&�����ӛ0�Q�-�_�{�~�4�c���leQ�}M�~���f���������)@�}��]�b�s�Zb����	�� ��'��v]WѲ�� .ˎ��T�2De�t�W��KO�-Y�%�%�j)�䌌Nd��u�吷����~�g� \�ظ6Z��)jï��rȕ>�\Mڙ��Yk�	����D�K_�a�b��s��	�j�'��A��^����`Ōs�Cj��5E�� ��±t��5���Z�vq��������c�Om+
{\�,�Nt���in��\.���Z_�5��ɼ�h����!�}�����MUs@�옢N� E�u?5<�^4)�	a{C���r�fۆ�'=:�`���P��g����&L�gB^L��U:�zW!v����'�C}�?���A��J��	��]jY�T��m���d�܌)������2��E��H��$�'2�a�{���S�n��ύ��>U�R��0�;5�s�������߼}Ì�9� ��3�}Z,��6$Ȉ��|��s�>@4xo�F1&3�0_op�bl���ZUI��p<����3:��Ɗ
���lP�D�D�q��^�uSHi��Wo��;F�A��sx���<��_xGxB��k��v�Ǚ��=�E35�X�ޕ����z�XP�LA�k}�V�O�{J���=̨rJ��gl��*��t�(P���nA�qP��0�CUW��9ƌ���{��R9G}=a�q���unFH���98�����w}�d��4�_=]=�2����<@SB���E/�ڷx�ɵ�[]R���ېv]v����L�q���0&+1���A[\��'��p��iN
O�o����r��zĂ!SNJK$���H���`�W���[�k��)��=D頽���H^�2�-�s�ު,��ֶ,�o��t��{(R���d8�y���Ƶ|@�Ǐ�B"F�k~�W>/a�ά�R�dV��8�(]�e��Ǩ+_������/o���U!�b�\��f,1k�
nJ BR9<ҧ�mil���X瞆�s�>�W���0���_%�Ъ�r�����3��")�m��KI��;�2�"���'G(.A��#��.
C/�քܥ�t<w��������P5M�A�6�zo'��}3^0Z_��1_GDk8�e�GtN��if�t]i��}�'ʩ�����/�}��6r{䥛p���u%{��Ӱ��UY-+NB`۝����UQ+/Y5�Z���Z��2�ݮ*xq�5#�y�^hت���X���2��W�&�Z�y�ox�!��v����5���׮��]K�^�h'lT�6��Bķ�i��T�")����M�H�S��Yaz�_놮KU����B�l}0�bd����B�	�f���V�-��'^b5�qwI!襙X��Ε�g=s�k�,{�S��z�[���rͽ�gU	���\����~��^��{@��Z�=���*Y��+L!�T؃��c��Y�{�����cVW-�f�qnd�Xco�&���'i��jM�.���n��j�ǡ�,��yq�ޮ6r�(H��h�&�ލ�G�_�i�b�����H�ݙ�EԪ]�5��"����%T2�q�M���z������
m��eÃ9ӓZv�8�t����&���usy��঄�����F�I���Sp�f�����V1x�8|P݅�)\Ւ6��w�[��{#Z~�漾�z*%j��.�v�[���񵤭���35ú�ق�R���Jq�7-}3`�t�ځ�\�t��i�QWM�P��a� �K�����s����P���?%��I�/��j)�-;X�cg���� nF�ͥ�^D��U�jI�t��X@���z�k��!@,ρ^�Quף4��^��w�Z��q�,O7߱��2�z�58�zc��`c5�S����6��c���V���y�K�֣�'��!JJ{a�X3��3�+JR�Q���`�RtY��JWxQ��N��+�%�0`�BA!�j����4#aHܰ׺t&|M��Mm6�9���o�{eK8�����H�#k���U��g6���� m����Y�`dT Ѡ�Ɖ��r��N�Hv	+�.�0DC�cm�G����K&���_u(̍��	���VZa���s�����i���F��;������&d�']��z'�jK\S��Rգ�2�J� w�b���u����l����1�E�4�qw��Zy��%]���	6v
%,,LP�@EjY ��10�I�!��=K���GKf�a#7�%Swݧ�HQ-�����mǬ�=Q���I#�n�����"z��qx�2���e'Ԥ�<Q	�tS�i�6[FveEO+�ioϏcn?~t�����d��D�A�B%ЧO_��a�M�K9��aR�)�|*|q>��ؒc��OѶ�ɒX��s9/l+m!od{�n�B�v�������#0�jm�Jhg�㮅��+ªM�"��$1gR����K:V�?��ڍ����\�BW.5-�-^nm��OQ�X�������n.R�=q&?��э��Hh�穵mOڜcF���xNvົ�����ۿ�����R����3����M�fBhP9�XC?'G���`D�Λ���rK5�C��W�H%�Na�=1��x���q��\�}�}��.��)�9<����q�?��S�IT�I����8�����nz2ؒ�?��*�g�ø�뷭�dc
��P�l����i�]��^�tRbǳBi�3W�νvA��3�Gj���+�?f���A�,�|�*�L��+6���o��Ǐqfн��@�rwX��O�o����B�>9��Ww��W<XBy͊%jpM�D��2i��j!fl�i�])�ҎA�B9n#�l~OO?��#a7V��F0��羼��h���)\3��{�q�o�0� ��̒�g5����{<�G���H#_p`}=��	�/aC�[%�1M�l;��)޲��/���{��rhڂ9I�b?/1PwK8$v\ԗlҚ!��&�i��ԏY���(
�KY���{`��봷��a���d����Mîʖ�\��V�l	y���W���:u�n[�ƞ�'�,,,���X�}�)�Uq8Ǉ�,s��
�r(�:�u��i�N�!"�>����k��s���-��C�ҕ�0���,oz�}-�3Q�E��Cū��nA��p�{��XCR��b����F5z������?V�|�󼮢8�#��My�В�T�o*9�qh�%wD%����5'i�S�szd��(YSB����EF�Ɋ`D(�8��}��ڋ�����s�D�<�Z�x�Y�䵊��u8*�஧ւ�aSe
X��OY�N&C/��R~�i�gYKE��i3��ν3��I�~��A��N#+�`�Ia��&P,���M����q�������GF�"̶Z#+���VTQ���G�Y
H���^�y���F�60��x]iB��׻Ĕ߻��5
Cʪ�D�j��!�Y�#�l�~'JVI�7��1�KP[���<#W���������o��ŉ/+hI��XL�t��6b�\�4t����c��׊�cnG�1�ɦh�ֱ��P�3���gY��kI��KiZư��O�Pr=t��w��`/�\b*u���#���ߑ����czh��6弸�I�����ׅ0Zz<��v�m����g�ٞ�����r����%qm>�Z�,>2��0Ɠ��q� ��Ac�:��=�;c<�*TI@�?�m߬�~�M�f��^�v��^�`�8�5ε���9���Y{/��Ү�w5b�sY�z���<*�b���[�ǟ��z�"�zͪh<@�8�=�S�e�ě�N;�"������?��a���a�;�aD_M{e��
�6Q߆�f���4W/K�'8yA�xf�H֝�vwxj)��T|��kˋ�Cdx�x��I�#�h=-����$ �~]���6چ�LT.y��s.>7Pki��D�q��_��jh��Rq��1����ky`�6�{I�ys���N���hq[mztWC#��	�j1�ֶR1���.��3CE���ġAQ��y���S��	�sa�9=Rc�>(qOOo��L�f?~�P �4���~G�-G��t�+� �])"���a�$��K�1�f��.R0�����2��tY-�]kҭn�>����f�ΰ�/�=e�=YC���Vw���Cd���,�eVCG%�b��ʲ�5��xhqb.�V����T�;(I|U��5�����5�H��}����+C�_m�7���k`�;"x�V�|�XF9Gw�)�,->$�,�f�o�G	�����9b�¡��c	�|U��S���^-���˼�K��c(����x8�oq�6	WG�dH��q��=O���z��z||�/�C@�����J�Ǝ�]7$�� i<�z�T�6!��f길����4�Xt��=��z6Y� O­����00��Pinު����^PP�0'�]B��oY�%3̤���E�n�B&����c���k,�^�Z��Y�$����Qk�6�#�,�<��3�2�IB��[���0Zg�p��B���+Ӧ�^���Շ]j�b\����g� T���k�S����A�|2��nJQ�ʸ����n��QJkJ@g�g����O?�P־��E��>3�Y��fJm�^pM-х'@�~N��	�^�>�d����)�	�Ɍk1Y~�	�Mb��Ҽ=-?����l ��d2���ރ���}n�Y׌�-v��r��ƈ���3�*�1&��F�^[�m2��	û£��.����V�?HإS�,�����L�����wޖ����:o�!����}���"�y��di�Ξ��Vb�U��a޻���r��`�@�� ���?G�{h�>1�zd���]�Z ��^��x�n��4}_uT�	;����E���)^�s��ㇻ��%�xT�G)s��Y���E}Oc��s���9�'Kԡ1�?���%�ЁHZخ
IH&$�{�p�N�����M��FB�㇏����0ce��RV;_�
�:NͿ���t����ߑ'�*�5��/(O�&.��p�o�9ޭݗ�����=���ZA�r�:��Ґ��o��rVޜ/�Z�s��EW,�\�	�c�ƒ:�Mh�ɕ�6����f6�{o�#TG���03���X��F�1���(��
�5�f�ZȞ
��v����Ε	���:T1c&�&��`L�AHla�۷s��πt?8ٝ`�&��%`��;ER��/��; \G�4���e��.�\{N䜺� =cy4���=�]z�+�9�i�S��m���N�y��킔Dl�%�Lȷ� �ê��;hY��@Fq���Y�c|�E�����0�c��6�3�Bz������X�S%V:���2��}��{6�#<�{ó�?�|�P"|�Cl<񙕵r-��4⡷�2��}��B��{iq��:�SjtP���5�o��j[_����rN�l��z�ޕ1[�#l�r.��������Ŕ��=���~wwx�q��'����x���#�P��z�2�M�BQpQ�hL'�Ug��<�B��i;Ԭ�zZcA�"c��}kw�[hBbB߽}��»��t��Cie({y��ǣ��Sb���M�	w&��V 'W�	�VVRʧ$�hۮ�ɐu��=6��G�D�19�!�+�Hʥ&=�Ge�Y6����Â���f�u%�<[Cʰq�|���U���v0�ȑ�=+߃�8�E��=Rx�y��{�A8Xo�W����ujwR!�{}���L����O����8�g��X��V?l�q�H�zdP�?���Q�����k�?��ShD�f~>��ꔴkڱ4�b(��~O��	`]l�H sqVc?����a蠫@���{ƨ�}�+��V�E�����/hW���q^����/���8�ZUB^8X�YFv���ܭ��!�dB���P~QW�x�t�ꙺ��y��e���!m�y�Ү���7w�BQ��]qQ�L�{�C�]w����>($:����\�.)/��z�  ��&O1cR�B~O^DܠXx��9{�Ж��*�r�
w�l� {]�����5�7�?!6F
�kٳ1Ó�Y��d�	H�Q�*���9������ڬ$�E���b����ř���¨[����`%v&y�6��J���UnpV{Q�$8���'ݲ	�)��~�k�
q9�)8w��2�N����~K��v��g��a���t�t�L���_g_xR�N� �����v��W9�N�{���{`n(�3nF�O��؝��� fIcڧ��0��,�(��+�`�Zv�#�e����X��?��f�����q�f�3�3ߑ%>������i�f
��?Ǿ��}"�D�lkuY�5��)����dT,bL6�nü��ߩd12����m��Օ�[\���F��:��v5�7$sg�^5��E�VZS))����Ә��-KK�r��+U@=#!�W���z-�c���z9�"�4h�PIὒ��4���B��؋naMD�#�Z��͜���d�����8�k��3�Φ�PH!VHY;�b�m1S�T)7O�h�ߛ����~�����4dy��/$����������Z[���(kiQY����R�����megWDȤcЛ"����4S#��@K��d�v�c:�sf;(d�g���l�'��2��g�y���-���xP��%��ı�������}�hG�Yx�U��^;�Z�h����k�����u%ik�P|���9X���~c���C�Q�a�/�0O"9�8�{�0��c.�9�H�e�d�����d
��1�NBkk�A�Ib;�CVu�*M^�0"�����݂�Z$(ݴ_��Uc�ڿ���L>w�W�'�/6���G��1�*FzgL�2��Ċ^ik�7�'a#!b�Oc-~fCi��O�4:7	��zQ�x��GvwׅІnƉ�T/�'�mVqǞ[xl!�<%^8ٵJ��#��m��@U8Zء�_Xs��.�$��9���P���T-˫y�5D��N9!��8�B��x<R!�� 9��@-�Q��St}_���ɿ��\��E�6eR�J�؜0��F������K�N�nqϵY�����5/|������x�sj�f���u|��5���e�D�w����i4�v����@���b��q��j���Oq_��M��C��4X���Eoj��uQ��U�*�8�����G��c��۞h(�ȉ���:>�:�w�Hɝ��#e�Ae��E�@�f(����c�DϹ?������f�2�j��5�
1/8T����w��S�Y���-��u����-����K��-Vi�=:~��ih��W�������Л���p�&���y%7[;�J����%��a��n���X|3� ��R4�d�����~|QS�Z�����91TׯW����s�1To��l�[f4ݣ��VٛqF�z�z���p�w��>�o]�\p���ȴN������K'�w�a�Z@�0�d���VE�k��(e<s�P��-	���͋�x���V����)�ww:�oJF�:֖	2�"���}�;��_�4������}z!��9	郕ɠ!KIɘ�@�n�K��8V\S�<��ZFp�m�y (P���a}�0�
P���%�޼y���ے���WәT*^E/��-�W�R���v5�
����}��뫅� �W�z����tN�c��Sf;��3�%�����n$�;�C������k�k�{���&��L�c.������pеrBY:��D;�C�V��&D��eD�m��W���_/A�����ʖ�`Z��*��*�6#�eUHKYdD�@C��>Mm���u�+�Iok؝H -�|~Sا~��I̺;\�����`�X�r�����&��zbe�[��I$n���}�~Nqwv�!���On����=�G�����8(�_���5��p�a]c����B:�*i��>�n}]��B>܍%+��\�y�4l�M�n\7��}�š�7��־"��2�5'���>�T\7�h�zt]I�Ͻ�|`����V��k�Z�,|6��'��M�$�Q'<�i'{	�6,����T��S�7���L�?D�Ǹ>�u>I��mЭ��OuŰם��a�Ē�6��Sm5�i�N8R��se�-H6�.�J\��~��F�4�/��U>�A�����Se֗�T/��.Uq|����-��M��Э�����j跮��qI��I^.�`D�ŜU��y(�2�\@Y�+׵��86\��
���w��w%���Q3�;�٬6.T_:��}Є�H��
z<��y�5Y(Ā{m*74+|_C+�!>�X��K&�w��,��?���\9c>�%n�Rf��sS��F�s��~T��u�pSGY������7�a��
D��|��h6�S�%^k�Ja���a����P~ؑ3�T_yF2��n���t�TU"4rR�x�twJ�-:lN��D,.8��Op38��4����*%Y�\����!��P�ߌ:�F�Q�#x������nL�SVS��û�ιޣU�U�����5
�
����[�}��4͆���s�퓟�g�|��_�� :*�(�0ts����_�Ҷ}�{ۻ��{�Ta��i�ڤ6���H=�mx�F&��щ���Qr�}X2W�]���
��#��+�z����2t)e-�::���E9/�f���9*4�gɎ�>��<%}B��A�L��75�,����YF��
guA��iO�A�Y�W�|*']�h�ؚ%`~jmsa������� ��;�+T�����9�g��V>m�|��b��8�aw�ʻ]�ۇ1��D����Z�Y��+���d{�~�^�|�q&����z�`!XFO�2�W�����6�{��-��ޅB?��9ڌ�Ӽ�(��B�������Ͽ�g�S����/�$�L��m"��ʪ�#hs���<������!5����4�U���������}����Qd�Iz�.p���汣ȷ��MZaH?~�{�>J�$���iG�:Q$�1��V˛�"j"�fM�n�l�"�)"��2eL����B��|*)������*���~3�b~�/]��@�62��o�Q��j@�ƃ$� cl2��%������	�i��IE���Eڈg�;��_�Jya��u���H���ޙ�y�5s$ZmQ�ՙT�w�QH��,u�m�UNp�0���txd�ґ$�X��G^,�"��Ncf��<��]��q������޾��)��8�y�#bv��1Fn[���"]$�ύ
Z7^k$���z�j*ma�p��:1Yϯ���/��j���F�I�R���nWF��~�1ĵt��*��=��c���YMԜ�v��5I�4RuC� ��/�	���6�a��7�F��)��b1����.��<[7�ks5GQ=%\h��}>O1O%u���P�����䔢��:-�;p��3���K�\{Q,��]��p�p���sx欻'��xg�VE3��X�6���6ڃ�L�]왧��,�=YJ�ɳ�����e�[��_/=U%�Zl���������x��/�&�d�GS���eҐJ��d|]Yq\�Rp����ʆWC�r����9�U�i�Tl�q�ֈ=�=�E��M��e�Kqݱ�'�+2�R[,dz��X���6��Ќ�$��Օ������y��uvJ����|���u4њ����Bi��<�`�5`�O\64A�w�}�k���hU=� F߮�e|R�MB���N�as`C��Q����HQ�]���]�&�p���ZU�`�1��?�&>�g��n�HCJ��S���zZG]�L`�a̟�(��nYy��T{3XcWxW'�Ipw���e����k�5�n�-4
6/��~,n׌�@[8��n0���Ѽ���
�u����
�ob>�*@	~;F%%�Z�+��9Ao5q���U?�i��H
�!���_%�qv�v6:pa=�W�D��^��0�7��M��F��>[���mkj�t�7���~�N��R/,7QgP]������2(��7�^i�&*=`�dH��Vf֭�]u�T����q-իY��^	��!i{�0�e�eRU�3�V�"f��>���'n�����!� 媝�	�:";YJB^x{)���1Ύ�P2l�1Tf��rC?�g!���^����ㅺit*}P�!9�s�5���}���w�v�T(p�:Ӭ����!�\.9���p��]s�q� ��7�i�g7o��!V��e��@0���t�>�)<��\���K��2m6.�==�VV������������%��8\�;y�(�dRjJ��Y��$�Ǻ���6�t<�dY�rH�կ)L��9(Y�5��͎B���X�=Z&2�B[2/,�\f̛!�%�NM�n��v���:��!��1�tJn*0 U�Θa{�X?�K}=�!7�X�O���Q8l����Ï�~{�~�}O������6�x�6��e�m`�#�?J#)����1����5��Ef0����'&ssm��x�F�='V3�^�	hэh�!/NrQI��Z��=/�f��Ъ��|P���^����F}��,��v��E��Z��}�vЬ�����[骖:lZ�R\�D�b$7����l���a^��Ù\�TP�{O"���Fԡ,<J��v�XpF��}��z��E`U���9[K���q���6'������1Ϣ�e��k���ȋl�#2W����ʹ��ʫ��BS��=zm�u�J#�����h��wKd7�9���v�xG���� ��͊"Q�:Q�XT��i�$���Ö�JY���eJA���1
�M�7�{o�YW!?�_ÈU����H6������oe���bL_��	����	�R1˯�Ε}�!ǂ��<����~�/.�Ph�Ev�"�-m'�x����R�^`�f�Ș����W���b��b=ٵ�3:3Ί�.�
��y�+%�$=�^ߑ=U�/�kp.gr-qW���*���7����}z̬1^�%f�p��-��3�M"�K�8�"�S<=j޹p\7���%��L���2����a{�����6�Wz��ֆ��k��:���i5<�Q�SЋU߫�Ԓ�|�W�i+�3A�E��������`�c�9�l�����>����O�&[,��gH!��̹IĦ�*�=Lqb�F�! ��	K����\�U�y�~��8.+u,Z/k`�I'�1��j����:8�cDyd��.�]qk&X���AM���\���쟖R����H1�����u�*�I4/�k��}��E�h����O[��!M�S	�>��6A�fX\���В�T���A�{S�c���w����MD�2��.�!I���(�L�أ�Ѳq������Xlͨ�.��B]S|����&o[؁Ę�Zt6�+�7����4�P��֌}��8��3gy� |�O���U0���!!C΁)1Q��_����5��ֵ��ŵ���j^�n ���TBh�؇i$1p�$��ưW�=���������d�kR�o���ZֱT&���nu:�UZO��7��."R��a,�#7-+�xHY��B�!�lr�#u��k�#P��ō��na셭[L�;Dh���Io�(�eY%k���a���vgH]�ϊ�Je��r�(
~H�&J;�vn�\9ن�nҫuG�1+j/�9j�`��ʁac�.�q���:d��G�H8_�fĝU��(~�}A��M�ԏ��H��K'>�K��4��[�%B%4Jzy�[U讐���6�
�*#nc\�F|_z-��Gͤ��15�w�����9�=��ѳ��5 �����5U4�4�$�fk�i�):!�$����r����7���:�U�*�1I�դ�X��1V����z�V(p���.H�Ŧ ������� ��a��AI
�(!�L���߃[D����̈́QU�9�ŐsU֬�6�nӖ������OJJE��kp�,�����IWܚ�Ʃ���ېP��@N��7{�[��x�������1�dp��þ
�8afm�0���0�4���:��'�4>5�7�^c�歹�Z#�i�v�ɚ��岦����mM�U�*�p�%Yh���-chЊ"�����P92��f��b��a�a�zkc����G8$��MO�X���{;q�\Uv}kJ��eۄ�k�˿iqӑ4ٞ�^s~�+�*K��06آ��yΌ��q(/R�������r��'3�>�������-����ʼ����b
���O9.�Y���3!o̵��� ���
[g��4��>�((���S�9������=�榲�$6�6��ņ�uͦ����M�
k�}�f����B�����ӳ����ن�&U��XYm��5��x��(7��m����e�{��1z�*.L-z_^�S�=�c,a�>�����-�uG^��G���a��Y����s��5e��_4M�5�/�#0Wu�}�Z�]D�Y�� ��a ����܊p��&�F�w�2!��U��Kx����"��K��Ѐ�r�H%C~n��-�w��.��G/�G���_�iM`k?��xm����I��O�8��!��poT;[������t�1�k-��r��Z��u��H�)��<���Q^@�1�q$dd�ƴZ[C*kFT<Hg����Zр�C���L�t�iڶ	���{@>.Ul�Y�L2lF|R��' �>�}�v�����Ơ���:�	pOI�B�ȫ0�����/�!�y��D_�� �qz��c<1ASQ���f�U_�et�Ч!�c�Ә��ء k�G&����>��q).�/K���,�c���5�QV�ZPG�:����F~b�?(+����6q=(���x��5u�2M'w�rҡ��+��vUC@γC�6YaX��Y�Х�5g*ս���Gi4{��	QYkRS��Z!8O�FF�]
�<ilUq���"��g�O쪬<���p��p?��
�~��pwR��wi0�,��3�C���ݜ{w�Ad�u�4t���w�0�|>}�|���I!�ݒ��}�P�/����C����QZ�\�47<`�?�jx��麉�(�����ZY8��>[)ª�!E2��lN�Wzk��4�ɬa�W�lW3�IN
��v��;��:1Z��=.c1�O�*7�2  ��IDAT�I	gݗ&𧁧R���0z��L�n�~�F&b�~�y��Lq�7�(#<��J|n&�_o�����2г��2c�
�8:�p1������#m���"w�4$�o;n�/#q\��W�6��7r#���7����a��&��s��N*��0�A�G�c�q>��g*he�ɍ=l���H��F��gaC*�bR`<�)�FU����K��u��ڷ�خ�l�:al�q�Y1�'������"�E�_�h������8�k@n��8�	�>fn�bCj���N�Q��"T�t����z��d�x�u�0����f3������%�l���Wp'[�=R�s��W�%�^��v�	7#���;��0>s@5�+����J��9h�]�����'�9�,d��x�7�\ϔ�<ǜv�}%���5Hc[�̚��^:���Yp\�U��;e����p�_+,z!�׺�嫇��L���X�<A����6 ��X�>�{�T��ǲ.�Di������.�ME��±�]vv�U��f�!嵆�����k5#NVc�7�r$���z|��)�����a
��XP��˓�b�E�^K�n1c�{��u� ��}u��3�]���<x�=�%����9�Ð���K�EU�̚��l<W��a�����Gf���aW�&Ɂ��i_�2ޘ����
^c�P!#{������Z���e��ƺ���1.wgRUz�{͙�Ƕ��,JN�of&��e�U�+ܕ��>���`����W����/�Z�<'��Φ..a��cp�:��p�d��N�b!e]skޏ�.������y��5+�&��!�,��4�:]]	y�r�i\�ɶ{>���Kn�=���u �e����x��揼��y-Z4K�ć�Ȋ���XkGE���ll��P&yRu�>��R��MM�&P�@-����%�� n��4�P��N�g5����"CX����)*�>�)л�6ɘY,�fL|���M"߁�x-tL�t���=�	o�M��Ħ���r�� �c�>�+�cx!.4zD7��\H�E�Y�(ocH�wFh4\�Rd�!L��.Խ�!�1��u�z�����ڷ�f�JқQ��\;Үkӎ�\U��v��2�ֶ� b��#�U�9z�	�(������g�����Â;�b3�@�5
\�f��$Ù��N�<6/��_Iȿ�nMB�cЋR%��	}?���2�Ӎ5���n'c7G�g])�7��KZY��4K�j�8�����XP�nUVњ���k��K�+��4���G���T�m]ˋ94+�V��=�$n&�����i�7~����V�Bm��\�m�c%21&E��wڤ�u(�X0>��p����<-�O$��J��p�0�.�>���`$��͒<| ���0�3U����3Uo0�j���-Z�N�\!�z���=x(/��<��>M��Cφ��m�>;�Ƴ��e���	u�}���t�/�ӀP��m�^���;k>y��Exw��`�v	�
�@&x>ǁ�1��^<
�| �T�㏯.D�zS[�0S��!�#������r�z����x�aLN�=喓�.�6�-eω�93��>I]ҫ�I�s��:xzO��|Pl��qx~�ؖ�Nʜ� �����:R��>��ub�>�(�8b�+�A]�1���cn����`�� Zܺ�D��8��p����n�7H�Z���C�2�uBX=�Z?/�j[o5#Gf��ݼ0��}��i���ڝ׉>�kC��.�I���t�e8ZCϵz�2�7Y�w������6�]z��q<����xNh+�P�D���M����sYB����~��w��N�H]�ۄAkQ��T�����$�"x�t��BW���g�� F��At���5�'�+�*x�#1��Mw�Tl�E^��ۉ�8,��f`lHC�3B�k�#0�녛���ND�c�$R���������5�cN�z�u���em<R&؍ɭ*8��HgM�B^�m'究�9D���1a���K�}QYbTN]��5W�o'�J(E�h��CtR����voHO1>-��:���u�"#�v��0ϠȆ�n�m��h��S��r�H��y�t]�'��J>;�p�s�*��-miCc��c=l�Ԩ��AX �]���M�T�6�V�F�=�Z�z��l�/��1}Ͱ�qgH�xC���^�0T~YU�	x�+y�_xy�:]]:��`]t��[Wr���d�dR���݉��?��p��JaF6h� B��s<%�p�x�G��'�YQj�!���Ώ�=��bL&a��5)~�^O�kU��#���Lp��V�N���C�8.FM��X2��w�׮zC�*f�F%]�V�1�!�7Dh�1�<ᥘ���v�hAa� ŵYQs8P��^na\�q`�3(��!�mܹϱ�V�à�n&.W�G�p����+�t�5�dmн�.��ޠ]_!�K꘰@c��\;'����Q�a���{q�8b�gŽ��(�̍{c�*qV�.�F�� X��Q"���+�;�$��f!�g/^%�=)�O�],�`��%J�[Ke�zTe�3�%�ۅ�~,�El���2��~{َ�1�BEX�E�gz��7X�_�<yįc���wn�0g��^�����%C�I����fVk&2�m;%ld�l� ��î���h<�������d5����$Gf{*�bC���",,������Z3��K����N����@G_�.n��|;���I��Jщ����F�je�L-�{E9����̯y����N�sgo�{���8�1����Y��e�����m��������>��>�����f]��gQM��^X�i_7@���j�m�U��Q*_�;�Z���z�!܋�7j�{�������"y����!g ګ�?)b}�U��UF�*/��!ͧ��ck�� ��wf�}�M��A /xʪ;+h�Lp�2܍�NcF
<���{W��۝Gk�7�eu+.��x�A�ג�9�@J7@�A3%�u�X�jX'[��c:E+6XZ�;Q�����i������a��g/�S/���H��:��S$�񸸙Ų�UF�AThg�����!�1,ǝ�k�>�D�.�%V�������$}�&�r���1AEC���^��mO�>�BC�������	RQBi���~�^���󅽚�e:T����)G���p�gV���h�02z�H�ﬤ彲
��ۭ�9�][�z��S���1����b<�+����G)���0�����3��팷�v�XA��Y����H��kF�U������|�����5��7�N��󚞰&�d�z�e�� �ˀ7!#����Z�G�o���yV�����A����+���pv�vM<�J��s�"��n1��@-��CN��t�#�9�!�58��Om0����)^I^x}������m�c��W��k�E9ؗkI�"OLV�=��������q�5���E�+�N�r'�p]�L_&m�M�מ���gx}�F�5�j��޴&���F����r����h=�fa�f2�aj�)D{�(�鶫� �Y�2UK?��^$~���e_�y�3܉eu5i��Xj�ƀ^N�u�>j5R���f�apCo��W�!g�ƀa"�}-w��mԻ�|�ӆB�deא���0���J�Y�����>/��tfy���G���8�ː� �'׻M5����}'�g%�9��Y��dF��65v1~�ޝ5�g9(�F)��{|��⌹�*Χ�$�u�<_v7p�x��y��� .wې�\���.�M�������0%v�V"kt*��s����	�(*p	�.����F3v�-:p+�0'�4��ܘD#�f�w�I��p3���d���J��Z������wԦR1<��lz푘����v�f^�$i���6��]1��#_Dљ�]����׼{W]`�P<��t�y��j-�"|Bx�zZ�/R,�K$b�:�4�ȋ<lx]WT��P2ۧ�9�Y�5u^�]�Xb[#MO�a�3�.S�z�3��� s�h��0 W�T-�#*�z_�W�9��Ė��]�A) �אF�L�ة��+\zivdf<!l��K8$B��s��Q�rc����A�O0����=1d��4�y{[��Q�6��F���O�Aw���k�S�����!t?��9C�Zq����R\�V�⫲Q7&�y�{��ʻx?�k5:��8�&�zTƿ��aF)��.����fCq3|��R}*r�Wş��M�Uӗ=�=>��A��<��	R�p�����U;I�y7��1�FQ�M<�.��E�o��#)L�[h�_Vvf���>t���/b�����x����TŚ��{�i�(��x�t��k/�s<�jц��%�A5�ә�w ��CX�*e&>� ^1W��7������>�cx�g��(]և���]%vL,D"T�cOh�TR�t��5BI&ov*S�%[��V��T6�G��e�ƭ�gΖ�4f�6F�=s����'�Y�/C-���2�偶~��t5z�����Pp�F��d�I�u��������t�U8��4(�nM���C6Y�L�9_��;�UO;������z䇳�I���p�7)�Tl��:�7+�SwQ���膕�]ʽ��S?a_��F���Y$���2]r��_�`տ�RMU�����(o�G����/,j���?iБO�l@^K���Z �;�N}M:����rH1P��xw�]���:�M֞��LIȹ��$���|��Yd9E��b�">�����,~d}�G1;B45]ݜkR��G[Dȕ���x>V�)７���b��=�n I�'͑5�"���`ڸ��Ŧ����M-����Ur�I��pL[��q�;�r�b�4qc�ߌ��1Rg6$��b�����SP ��p��=ZT`���N0�z:�	n�h��y>�R�O�t1�	ͦ��q��i�O���	/,�u.(Mb��C��!|2C�/��:i�f<�pΞ��f�]>)���N)�6r��F�z}h���+@��n6�2�h�=�;l�dwu�N9��e�[MB����f� q݄�R"؆�S��tn��?����ʃ����Q����i�����RHL��ӓ�C��;�	K�	�!۪��"I�w�G1��~�'�CD.�h��B�gPO�X-4R�����G	����	����"���v����e��������w�^)u��/G��x`��@� A^H��\a����L��6�n�D1q*�F�D�X�O?�l��47w�|'�?˦����W�1�O����<���c���D�"}�g�w��߉�0FT�	�J3�}��〷�G8��M�
�:��r�`�	L[33�����o�H�$l*]XP��Uįm������E�f�	��L�u�L���M;�L]�N ~�nM0��DA#b���u�p�G�������R;��AL��b��s�M����=xpk� ?j�#��@�g�0I;�v-1٦��'(M����8>������5���h��;��MP�Ă�����l�E�xB��T8@�1�t�1ȭ��� ������'�{Nx�x�>FӡF�����-BUE�#� )�V�|��`����X�f�8O�p/��E�v��E�?��Q����f�s���#�[6�ys�6�A[��zX誅�^$l������q�@)9����^��t�	��ɪ�h$�j�u�
�.EE�(��9Qm��kD(���$ޟ�fd&��y�}�q4Л- {��#���-Ռ*mP���Ml詡�OX���wj�*�Ǔ�}�7�hgޡ��!�z`�Vd��j�lE)��p���~�K��(�5��d_σOcJ�ٌ����L9?�{^+J{�@�Տ������bh R�!ve�1N��D�>H�V�fS'�a��@������{Vq��$e2]�q~�|@����ц��XDĔ�Af%;Zy��y�͹��S����0����Vv9_���٨�|���S�.vh%〳�h��X��ٜD������kRĢ�����*�1���_Ս���K�qz?٦"6<�y�6A�҃��$��ya ��/�]V�6��y�@̴��}Lc�������S=��ؘ��f�US���& e@�h�w��>]"2A�-ǑTC��;�T�HkN��nȉ���R�C�3�� u�徺�:9@P�� q_,�.��{M̸�&��5PKjw{T8��M��t��m3WǻEڂY�nL!�*�������4��l� Iќy��7T5��ڥB�ۃ!�Jb��!׀e�o��l+�ӎ���v��0
e�����͈�`b�&�s��m�vtϝK�3?�|��s���3	��I��#:��B�a������Ĕ��Jz��ɢt���"���1�M(��!�,�/<��c^��b��ĒyBk�t�dβ���Aw6v;��	������`��:Y�S�ObJӋ]�����&�d�K��ן�����S���ژ���)V+=�D�����?g�F/jk�dtb���"M������a��@*l��b��T�����^���$��"��Q}gI�����N)%���Κ8�I@�Y��p8�w�M�az�Q�խQt�c��p� RدJ���r�$63RM���?ޛ��^��?p��5v�EWn����j�. TgP�	 Nϴr�����{��G����L��v�Y͢�d�N�Y�`���\U�{��-L�nOL�H/�	�l�&R 3]WTD�C5����c!��9�4IHDW`���_d�P���v��+��F��+�p`b�p��o ��N���θ�"�r�NG��Y6w{ӟ.MDӽ�������1���ʖ���tϻ{�,�m>�bL+�7چ��Kz[�to�]���3�<��NW�%�!:����@#o��{t|âzѝ�b�fEυ��#5I��y����K����M�`�#�Ct,M#��#��^��f@2yb��\h�����>������ҭ�Rc��c;*���ӥ� �3�#�JOz�?H$ulHr�rI=/�*89��;�����K6�i&
;����N+���`b.յ&�6���$����c�V[�lni�F��U�3��ȇ�F�����{#R�>�J l�x����ղ��0�����>��0C%L�M���ت,���'A��xx��h�$�Ig2Khl�`��K[�\�`�X��b��;�H����`�)���yp~o�=�Nr���N�<A++)@�M�(N���lܠ�*u�:�K	?�QQ}�6�4i�dg�邩����q�1c�������DE�y襠_H��C�7xR�@�i��w�Nt�y�+<�q�l�OQO�{آO���N~���>��Ϭ�|O;��! d/,5�B������;�Ko�ҟ,,���p3bl0]s� r�úA���1��@,-���p�uK��Q�H��'"+�5�C�~����x! �� �TPp�Db7j�w��e2�ƙDŗ������͝�X��� &h�ϒ�v�f������4̃�3�w�.��Y�d���S��	�q416|ﶽln��dL�� ��rPR�x�ܝ'��
�̨�ci�10��mf�us�R�N��Dj��9	��n�!�rѵ�7�+L7��@�̷� ��3j\�$�#�ﶕf��$Q�g�Y�����A���&��<Y'"�#X�d�1���S#i脰D�Y=p�g�S�$�o��N����g��B�Ung;�@DW�_k�_��6�σ���Q��_�<?Γ����.�Ё�nK���+���-���L=BUEH�[��g�\���LR"!^%��.'����'`�`%K��l��< (DH1E{p���l���Z���C������Cc�m]�{�>�v>~���0b���y��㉁���^��~�r~��f�%���6ez��ٳ�a�OM��%ĒH&�*Q�?�gQ��ھ����q��^��&+�_ڕ�9 ۜ�4�-Ggc�Ϥ�BV����q�_$!���+Uԟt"�!�M�jQ.����%�#���!a�1]��qF5�6�z3��v`�k�:B��"po�6H��D�%��2.�δ�FOv�Z���Ү��a5�OD�)u�dJa�pg����A��ۻ�	~CWD�@�3V`]��i$�Q���mW^Bql�����cq>})��L�-bZ����m����\���30��&�,�H
S�[����Z��Z����a"��8�0��>K���,�9��I��"�6��_k��k`R�\6;k���_�RH����:U�c|PՅL|i�%�$Q	��3JC��E���ee�G���'�a���4 >�c ���]S����߲��������Ԣ;���CK�������G��>��PE�;�\b����}1��5�buJ;�̼��8�T3˞M��Nc淢Q��P[��BR��0�VJ�6U=v��{���;�U�sN
�����q�fR��@�����NU#�/p�ֶ4�I3�T�R3R��܏�90y�1l��"~_�B}�Y�ҍJu�>� ��������2Qz8��t�V<X����v�/�׿�e,�oe���������yM&�^�L�d�M�F�xc�s���ǐ��a�&~����?�aP}�m|�H��o��D���d��iLP�>2?Z��cvP�&z>�s×f�ȱ���j�1Y��)�4��J���8y�y)�'��09U��7@*�z�Ӿ��!��h���U-2��g_�g�᱓�|�ޚ��6�|r�q�vы6��v�,a���J9i�ĔΙ��+E��bzc���@�9(��E��e�̆�I�4��S|�_����,d-��s�4��)���7��6�w�X�o3r�xJ㛞��|ǌ�I�K��{�4p M Ou�8�1�飴����u��>������$�r�s���i^1���:���U���4�_S.�JҸĴ����Y'$x:<�%YDD��RP��C�LE�l��B�>�x����N�d�A�ؚbo�}���x&*P�����Ɠ~�4E�v;��0G�jV�Ad52�r�2	��0c����Ǌ�s����75�@.����}y2�h�@�6x�/�`��B���~����&��d�ai ��d���F��w�Q/]���i>ۀ��hFX��G��!`�ý->ӗLnx���b� ��C�`�8Ur��,��E���Vك�D�r� ���P��{�夻ޑ9��ޓ��BY�jͳD;��6�{C�v� G�D\���`�>!�g;�p`�ub�:�>��;�ۀ����?���,�,	��!�8��Tل Ф +tC���N��DTz6����Y��&S/D��
��#�ț&7&�V��}tqA��c���Kx���b9b<�=�;�s��2�����������+������7��������n
�����kRk�����:�m@s��g��2w�̂Xk,�lR1��X���4�.�C���k�8&������@�i@N�46�ݒIUadv�jT�>	Ŧ���[ R�)�l�=4΃��Wa]��h@�oTi2��|�C_b%���?�������d�fH�HR`
�~ro�$Y����N�{�@��&R��wTkzr�(�ɂ\P���Dk����f�sҡ�ƚ�q�?��lOY3�5��g\�}�ϗt��"%
�0.Ztx�8p2���m$Ŵ�DV�d����|�_��W������/�
:c�g�2֤n��nK�����E��%�Q���8�|0���Xǌwv6�x�00	^0��?g�|:�o���_�w�������˿��f%4[{����H:�kp~V7J�E�T��a�;a��t]�����������Xw7��v.%�Cx�g�G���D�a��˓��f�qi�>�c�'��c��_L���?D6~f��œ�������lS��ꙟ~�����?)�	��Ӏ�����d��!�5Ʈ؁N����{j=����L����%?�\w��RV$�������;Ğ��G ��)�^l� 
�جʕ"̏>!���s�8K�jb)�dS9�d#�'6|8�؎��`�,����G۔`�H��;3�O���v6ٸ� ���_��+�/<0�!t�GlQ�����~Q�Q_\xG��Iz0U��+�@Sv�=�D�运I�4r$�u:��|]Rt�d��Q�-��QWu ���z�=�m��U5Ei��k"�t�  Qw|1p�Y���NH�6�1�A�|�f\b&4��f;@
#y��Y5���y�,>�4� Ԭ�#�'�܉��l���!hOl���".��i6�G�;VU���H���B5h�9X-T5�c�7M�g�NyV+�k�8f_xM�B�ϼΎ-(�NO7�}I���0ie� %z�]6���I�@��8�;p�>����:/��_���;o1��͓�I��Z&�G���荥�F5$9ۙ��Dw5�AI�7�^{���vѢJ���6�&Ʊ���F�t�	��q�E�̏?~��b`K���[T�B�rG~��#V�"D�E��?�Ov@��+Qh8[��~�`"��fL�8�<�mV��T�`z;�h�x���T����ķ/jy@����r�q8ɑkƼn4��,V�yO=�us�ЊI	-(�-q	�UG7�9���.~4k�m�KbάS�v���"y��������es5���ޯ޽Z���'��HP��C:oa�%����u�׌��xSMy HY�F���6��M�H�3�%E�˃:���,Z]��d�9��$-��ӡ�<�F��0��t��j���*@��`����p�\�Rs��E���c�J��$���k0��{5OC�+*���2�L��A�����q��Y�|�b�����H̡Lq�,|-�`����9��a��;T�/���Z��/�#���� Rb�Hb��*%ܚ{��X�+@
%+��-H�;��x� �s�!��G�j)��)�����b$>�'9N�rT��M\V�E3aƈA˝�@Ҹ��:�Im@�n.�Fħ������.F���>�]�r�c���l�
}*]]rR��R :�;cGd/��^69� �Pdb(�C�^Z\`kQ���^bՍ�33;=�.����:M�w��%��gb�o����S�Md�l��ID!'�F��`�:{ c�"��p��l���A���ӳJ>����1�/"�Ѿ�I����xP�)b�)lE3��&��DU�aO[b�Ѣ����X�W�s
5M�󢙖l�8�=�)��4���X��zW,��уC�C�F�G�ݯ�2��
�{���I�ݵ���%H^:N�[��%�m��0Pk�ٞ1�ɲ`���w%](��Ү	�Ķ�?���	H�DS���^_n��i�#xF��5�� :���:ݜt`�H-anWjv��i����礉�h0?'_q	�&��O8�l ���|v�]N6�юBP��,�KR���I�N6��OWV�6Mi�Ae�P�	��=�l��s��T��޴��e��,��dfQE'�]a���qԲ���g�A��fa
$�a��~�P�O0���*���ō�Y�lN�Å���q�]�I��)x�t�>�`$�(n<��؎�8�	�뵣�������%���##���V�L�v�p0�}L|�Wo���G��Ǩ}�>�A�8T�)�8��/Zj����KU9J�x<&�fZD_}^p��njJxP��;5�'񝎕�VGě�:���Y�p}Qi���F�!8]`V7'a�f�[<�mgKE� @��&z�"��8���i�K�/�I/����?��z` i�@�T�VY ������*�hDF�zF\�:�0��p�M����/��FM��"�r3Q�C�= RZ��Z�7��&Ou2#}�.���}�4�E���}��.MZxM�6�f�� �}��U�<N�hd'����󠍃Y'���h@-�Ɔ�$�Q=���B����98��vPi ����P�EwP�m�0eL":����b�����ߋ>�2v����� �2~�|G������i�0`�Ht'8z3�lV�d��v�������>�g1�
36Iu��ީ`'A�{�1��,<�n�v�����m>�T��Jz�x��Ŭ�-�~.-���0-�P| �3Fc��и9��Ɠa��;����5� `�H��w��I7?�=�{β��>����c�K����`dAEj��n��T�����G��g&Jl�o�;oܹ�Ã�����K�5�g���EQ96����P�Z<;%v��p�޽#ϓ�ӓ=�7e֣��������W�k�s�c�{�Pi��l a)0VtO�`��ͭ�"Аѳg���8-��0��yhJ���x|D$����h!Gٍ�U.�;4�6��ܔ��!VgD�`�]jw��頣�����b�<�S��a�07���߶���I�x4w)M� ���X %���16%��A��0!�"Z�RЮ���;�0Ə�+��ݫ��� ��VB��ł��q�b������.�n���,�A
N!.^��9���;r�x�V�ް���{m�	�z�xt�P����2���A�)�Y�񁹀�kp}�`�e�i�g�*��G3yz�A�,=�����_�x���*WQ�M��{�s�K��E7�5�8���G�ͤ�a��t�S]5tܐ�I�I*���O���4��e��,������2���������.ҳ@�ZX<�3��S��:;Ȟu����j/���-?N;��ٛ�O �y�01�Dݎoo�}��3����,&b_�6�T
`�.>�K/����b����CmL�������7���?2zۼX\w��K)��qs0�z���n�����>]��Ϸ�p�9�c�C�Q� `U �:�
q=r�8R���&iy���f��˓�ؾ37[�xs M���Y�P���yۡN X��ac$J\���Y�Kp�D�mi~B��5�~D4s�� x]�m���3��Q��`���V����+洺_�^�A��1���$��ōߧ/�Wk�ȓ�v�&a K���*$��~a#��SA<Jv�k�F��@�w�6�0d1��A'� @s�l%(����_1�R�����،�榢��1xEę��.��4+\�	T1��,�����m�60!�~K@O#d�$�175v��E���Z���W��BM�ک�g��9h+�pe@
qv2���}���X9� J����m����\q)nV�fR�@����ޥ�|��w��codT�`%�h��D����|�86E	�#�BkǗb��.Ʒ������E�â�`Tb�#����s*�`�c��z���d�h1�Ɣ�L���	A8���Ul��^P;�/_�Q@�z��ȃY�\��$����,��!��
�z:����0��G�tF���>X�_�N��WY�m'�YRQcӊ7n�x�� �	�J�{���#]u�'�gT0߄��7�z�]���jw-3�&c�c0E�w ��U���->����1�g�A&�%��R�����#�g q	���oR�F��JF�HL�s�4v�X �6485,-./����	{/2J�	C�筒7���K�F)`�# �Q����y��(���Gm0L3g\�J-|�@st~��K�T_��
+��w���:NХ��c[ո�x�.7T1���<a�Օ�?��@�xP�T7һ}AR�����U�j����epOA�I��SO�x�,]ش�sK�/�K�L��|9ɤ�'��i�r�dM�~�n1�x�Hu�1 �F�|H�"e���n|(�4�(Vuou<6�b��bv�.CW�!a�d�M��MQ��)�M�͞),@�O�s�d�J�D|�L��I,��b *y��x��#˜��� 	fzL�R��}n�p�]�?�% ��bFJ%R�R�@:���
���A/�7ڀn_z�dg��g��Ydb�����h�;U;���ݬfA;�NS
�FY��~���/~�?��+���GZ��実��P�oi��@:���U�\���>�\�wI߉��Y�M(�m�)S��	#�;��Ǔ�$�g���D?��O&�}YI!���T��O����%fך9�!�.F(�B����Y�j�[�l�hN�Ic��J�c�w����)������-���=�:��'w' e�k@Sټl[�?���&h���ӞKm��zCq\p���1<c�}Ľ��~�J�{^:ލ��q�c��p���4�9��R�n1cά�#��P<�
�=��8ݬ,b�L��'�)��,|�s��_kI�4�󄟫���Y�O��U���f�O��u��%���C�p��MA_�m\��7��F-�{0K��-�k�X;�{�b�+i�t@Z�M<y�Ѭ#5"0�>��l�����M�\'飙]���JB����a��j��-�5dV��x~TFꢽ� ;P�T֙��6���K$]�6�T����5[(��"&ZŸ�5�~�����Yu�Q�쏏��{̉Gc�����|�r��8����=[�b�Q�j��w�����؁7�&�vԏ�YpƎ"�� ��<�� ��I�|��z�&���c0�i2#�,����p7/�ğ�`;C_6�`�gF*aѳ��pE���_@�����2�� _x���6	����IM mm�!+l 47r�-iL�X���:E{�9lP�l@��vf�.�6���9� Rv�P_�������N2�e3H�Z�Q<]���|�h��n�\s3�!0v0�l^_#�� ���1�K����m��r�����t��e=tQ�+y�נxiik3	��qE��Ů�t��~[?04�'1`����RQDs��¸z�o�P��)�E�A�;�)����n5��	���[�z��(��Dݥ�8X%Jt{��\5`�,�ߕSN�fp�]����,pu�0�q�*
\�ħ�a 5�ɨN��KtW]�Xۅj!l8��c|��P��Q;�S�2+r��&�btӒ4�=�F���oǞt�$��*�h��Z��fx66&i�h��Λ\B/0Ҿ��u��~���j1l��x�q���c@f[.���OyG��p�G�5?�6���%u��v�����:�(�8��I��̶�l�$e߮�)�9� ����`d`��?�M��?�_O��ȶ��>UDxi4�c4���<~j�����-3z��]L���sН���}n�g@��|����8K[b�۾\���zk����\���'�$�iy���F�;7��8j�SG��fZ����([ؚB�I�D-3���:�?�3�����~ڷ4n��|^scs�~�e�<�')s� �a�>³m��%@��v1������?��5ƣ� �;�6�Шv�<G`y�B��u�O����#�σ4J�����	PM䆈>U/���	�˨�	}�٢zȽ��#m�3�rq�)H>�Jl�Ew�C,��飃hX�OdnD?wSl������6a�Q���{��< �t	 G�>*��8~���׀�gI[ly�V!
���D�v��:>��l=#8�8G��{6�v8��\j�y�nF&J���>Z�M#+���0'��,���a3����e�O�v��O�B�6?;;�\�J��mH�~	DGc#��HGj�X�S��6�Jn��?�����z��
�T9����JC��C�C�]�4Jβ�sm�21��i`���ڄʎ������|�U�-���:wo�]��m�> �ȅhA�Q-�q����댯��Ɓ�/ ��wp� ��rI���#�����;b�}�Fuv�p1�����d�b�,�`��j�������g,L$�3��<������"_���J3�΁��AYx�u����9���^=c4�9��Ճ�W,��um���+`;b������ƿo�GW���st�oQ9G&8e6ډ���fC��Lm�����[e��uw�ͯ�(� hj1 �>���8`�q���<a8r�<�E;�o:���Z_qb:(�`��XyL�ܔ�8 �ʢ�2.�e��cp��!#�]���������[���^�7��V]�@K� f_n���f��e\�&k?5�<��,E�:�Ц(�F���rB����la���mV��\
*�Y{�~��9�=���u���Aԁ�sj�y���_�~��8v�9�}i�\&h>o����t �wW����<zǋ�Z�
]��qu����&Z\����G4�L`��7ճ��Y�C�Թ��E6n�S��29��G�L�g��[�lj��Jٷ~4p�pY���[6��MX�`�I�͒�n*���t��Z�.�M>7_�Y��)�VL�w�o�|o���;���M�r�Pl`��U!{g��/��&[far$o<a���:��n�� Ew�zYL��Zb1^�n�Fе��׎,�>7�M���C�ɀY���mp�*�9�����t'�M�jac)����@j��B�r�a^��{�ͦ���{��R�{eڞ�Zw��ڤ�\�^�EGd8콺�z�`~d�G�!��I�� �7��D��u����aB��قwDS+��0�C���=���H��%&�EK߼����E��:+��ƨw��%��#�z�#V&�R�F��<A���R�9�E|��@�؊۞zTz�u�{�-.}�4�5i���i� ������޿2�����?���>/��-%��[�D�$>|���x�� K�p�9�@4~�^�X�� ��~��=/1R��	P��ԘW���n��,V��ڱ�&W�e�4	�د��e'�Os��7�3�����B�� �Xw�`}��5�ՉP 
��&m>F�62п+�Cx���Y1�4���]ǅ`$*G���td=hG��*���f7^L�i�.���h�~׋ξ8h��Ş�aE)6?�kǎ�	@:�4�~�*+-�j��O�<W:0�ة��f�طE/��yv	Qn����c�ʌ���.vL�<ҭ�&��Pq�U�V�PeȮl��)r�]����:�m�������+��G_t�T�a�����K � �O=�0d��x��f�� @Sd��u�3S�9v</�qNxD�w�}89�Z,�՘���C�c���h1�e�fX����������c��Gq!b��m��<)���p��*�4��# ��x}�����$&Lы+��B8�4�
>?�G���q=gz�Y�a�g��+H�Vi��c�xr��^�Ϳ��u�7�=�>��H�JŁ؋j�M6��`%�;	"}��{��f@��M�=� 1�dKWA@	�3��������Rp�kB�[%��s�	2r�Qⳝ?_z6��7c^����v"Fs(�Ntט}DP���5��WQQ0��4L�֢��=O8 uy���(��2�̀�K(�wd��Ζ
C�<��;��#�����zJz6�����C�3�������{����T�h����TO%.��&�F�z�^%�Z7_xf�D����.�h~��K��o�|3������>��q��zv�0�0�{��`Z"C�i�-���F�>Yܥ����+��Ƀ�f�R��d[SH�%�GfJǼ�<3KH�Z�d��ß�WJ�z��w���q����Dk�;�Y�]����'{�l¸��߻���9=�JT�)�'2�N�+����#��O��,UMw|�,7�{��J�{zjY��0j���Z�=Yb�Z��܃чa��$���a�XI�P7��Lc�G@����ٛ��1�����=�^+��k�R��Ō�J�:�X)�P� �'����H@�Ӹ��'O���8���D�1aF!�Ii���D;�kb֠#��ti;�-I՛�UI*QA) d��B"�Ӑ�Vٍ�{��w��zz��u��@�TYp���|���l�{<��X_3X���V��߫���X�]7i�S��΀�Pnwţ����2��M�A�P�����5��{����j<�]I���f��F:n4��Z��g\1S�G�mAk:1}{P���%�r�'$Lц[��� �@���v�~iY&��0)�@����.�U/!|�>/Ɠ�DQ��3Ҹ����V�O7(1 &Gd�3-	�-1��{�u>ivH�t"���F�R��8�J�ܳ��q��גkt�c����i�>U�+a�K�+v�k��%�u���ˁU�rca�@o �z\�O���4�J��}��]-��:N6����ź���"��9�6Aه�	�� �c(y#�Лv��Ƅ����4k�i�s�]ڵ'�^fU��F�����,��A[1Vj��B�Ǖׁ��X���K����v�����Ez���d-�W>\���sK'��4��D=ᖯ��5�x�Tt�7�u�tI<��NbG���@��4�}�vO�y�Vg����f���w�ڷYڮc;#un���}j�X��t�ˮ�l��[��ݳg�ɍu��
q��@m4k=18.�\���hZ�3��?B?������G�GXD�8�:#�X�w����^�؊�x:!��,6��1�K���Z-�[̴�cvYҸ�����������i�<^�׈ۭ���6 �����QL2�WP��%���]�@�a�
s�'��c�3�=C �#91�⟔��:Ê��1"%?�<�n�,ј4��z�e5��~��R�ž�~e`K@܁p��Zߤ�lu=���
u�Ł�A� � ��'j�:�
�a8І���z,��"ѯcvj�;Ϣ�`�1�l��ll�(��w�^�8j���=��C2Cb��Ʃ�=�~�c���zO@
���ryL�Qױ�Ī�%ɓT�S�d�U�����n�x��e�[Ǿjמ�Q����.�xk��(�0v�Ζ��E$�.�tv}�'�c�׵��&J?�$���Ym�Ā����LE'*�}P5���L�bv�b"����-~
��q{�;� ����{��ؾ�^w������$���;�U�5�46i�,�8�����r����Gwǡw�M}�s<~  �Ծ����N\��?��-m���e�n��i����`fRa!�*`�3�$�* ��w|�R�踿]��ڬ�ݖ��xi�u�z�k�KJ�`�I/��]�"���¯��cA.�k�@P�Ϧ;�a���1n$��AT��z��/�čc��& ������6��?�	l�$�����ՁI�8��dկ��8S ���t�X���k��Q�/��ՏetO�W^�
~�\��R� r��p�;�����M�Sd%
r�?��N⥃@ѻ�ٔ�t�:@�j���)9���$�w*�����w��GZ�)]t�y���!1��ë9f��J	���i��֋G��(���F0��/ǵ�Ղ�t���6��E@
���
u,��D���nG���2I= �zH֚��`G��W�滭�A�����G�X���-���+������&�a9Xb0�=5q���s��ݐ&�ף�D��$J]G�@f���Q �jD�$��Z�����KA-h��ͬ�荙����=7�9�"aS��(��̀ H����w��{Q`����<����y�^_�$��5����<�wJ}��T~�����籗��A���D����@ʛ���H�Dן��~W�S���H�\�y�����z�����Lf�O/�k:�X�pr������\Dq�F�M�� U��� c��GRE8���@���&F�
M��h�7��x#�L�ņ�
L���<�~19!�d��.� ީ�����E�L@��^�d���c�Z�8���z��I�d�#��X8B-��YGRJ�D=,<���X�b���z����fOe�Q�ՍVC¹j`2}� �"q����[�:���GuE\��~�>@����EşW wI�t]^��w��L B*�y��Ӂ��Yy�n@���̋@�\��l_w[�1�sSQ��V�|cA'��E6�қ��j^R�Fi>�|5̺6fY!77&j��A�93N����{�\*MǬw�k�� ��%�k�'W��m�ړ�i��A�=�O
�&*�F�y���q����9�l	/�K����$�y�Ǐ�[J#��%1恋��5�:Mc ��	"��{P�%P��f��8�4�;"�SL?�+w6����#�žb��|�s�U���D�����`:YlQ���gi$�޸�۴��1�B��H�U`�ԯ�l�+���Jg���;L"�-�0$�1�[��X�L����b�M��z��&���[��ӳ�T9��&P��r\���z@���V_�{�"8�@��'�qDǺXc��e��&��H����War�@��� !8�v��=�dI���J��θ덉n̠Ӌλ�&�_g�k��n���!�C���ȕe�Y�����u�n�-y|q;�l��B;�{�U��I�##!@s����m "sd0��@��� ��wg�Kki�d�j��=ð2<'3͉��-ň�4����� g:���6�To����9���� ���w]b�׋�y��J���4b֋�?Iu�?��q.�nG|Y�-&��ᦟ8���T��� ]2#��DE��Å�1�
�$����Ã2Le#�s1�9<^ǲ-J�j�U�x�PxS��?�:%�E�f�\R6W�y"�.�1��!�v�Y�l~�Pl��r1.��Z����Z۱�g�N�h�L��̝�.���'�-W���ا���%u>(q1�V��R���z.�_ �f�O%"[X��h���=0�"a�4#]`؜><���c�3�k̮���q(�ބ�e��9��Iw�)��o���yw���6�y&�N�q؃`d�>���3�,��`M$M�����溢$;җ�+.��a��\���j��P�,VF�e�r��b��]��� D��+����})MN2z�@�L�&�(�3��qw���5Ճ� ��l�L>�-�\LV�fj;>-KbS�H�)�|�$Q(2�Rkc��}n�fD4r E[���_�瘞���Q*��+�e[�<�P=�L�@T+�+��:�D9�ˮY[b<q0�����T�P��4]"j�[mA�(a�]�O���6-���9l�A[v�W�i%K}ܺM�#�Y��e�HS�ϓ� �Ya�6��Z<冲}�]=k�.�Z�y��{�N���zk�	猖����_��Q�����@�AȄ�� ��, �[��f����3#%�R)��d� Z#�@4l��!U�A�QM��"�I��+��O����i�ACT*Z�Y_�#�:IY����I��	��C�ω�,Et��;-��Er�].�' ,>9�~�`oL�)�X��Ƭ���a��<Yu��P��E�n�����X��u_��O`�e�p��P�q6	f���o�!QcM9�b�Lm�Z�#%HJ��O\� ��,1�/��,��������3�-6��o	�`5���/X'MX	QD�^�u���D )�#�}
�al��l���%Ϣ��O�cٓho@�hb=�*�.������\��V��CHR�D�k��� ҶI4w�w�$RM����ig[k���XN�ٮ2'g�)�Ӳ��^����C#ӫ9\c�Ne�Ff�cq�ꢀ�M�&}�j��PƋ[1��vI��N�\�,�ҕY7���tSU��X�hX��)���D�����%�K�>R��AU�TQ/	=E3��7@}�����4^��|�[��b���#���R�=oLUＨW� ~<&��ę���C�D]�xR�tڝ��}Y��e`�����y��hC-d�� 1O�n9�����íD�� F[�I\\&U#�r`.�zSm_��U+.L�"�F�ܬo���ͱp�İ0$S�%L�D)t�5��`�S�X���cR�DMn���!IB�~��lRDS1:����^�����hX�T�p�?�	��}���$u��!)غ�[�Y�i�� :Ƈ��Gg�� 13�V2H�N�$�[��{� �����������:Lk�%6�����b ��W̱�iE��B�� �����b6�����PxH1��yt�x��v13���Qi�@�:/��Q�hZ�n�J-L�I]úF S�����/G�E�A�3��I�5\["�-@��y֗�-�D����$n6���	��eu���Ԣ1xf��z�UkW<X|6[dL�V)��ժo&�-�d�U��-v���F�8s�%�=��F��G��*�%���*�k�:0�ثfۍ�2(.�G�D|X0���[1[k:�k3Ь��o�[�=.����54o�s_
�Az�QY�6W� ��gS�����wi�$oDD�.v0?ސ:�����+|d����a�j�{�� ��8�}r�E�4��^/j�L"��%���/�'�us�k0c[����g���7d�ۊ�c�� �n���߾��u��Պ�f�Ƌ�YpR)lV0���G��X� ]M�����1�礛r�7��MXg�����<��l�����tL�~dӽC�	�`���S�q!jz_V�2[lԄ�(ڇi�7���']�b��^Y��]{��m����e������!����r�������h�5 �HZ|�;���6f�����]�&���T�V~ڝ����Y#=ZyY�]�\�nq�,#�I)L���Z&�EAG����{\J�Ȅ��x)iPz&��1e� 5L��@�Ƞ�46�_����\���dS;E��8�4�e�\Nr��J"0�����t ���URq����:Fvz���Wm}��:�Nn�ld�G�T�,.t�^ց^��e�ը?�S]�	W���2.�+�ƀ+J��i�������x~Cɾ���� �]+7�Y��*&�[]�Ǵ�����y۽���>��llPE(I���E�O� ;���c9��me��u����{#�2�A��\�0�*@�mg������ы��`���Nt6����������|d`���Ed��>���'����M�>W�zrd��ű�b`�6�V��'2u������?XT��W�M,Z79҄ �>�QW��ޞE��>���`���T/�Q�������zz1 7�H�:��g�VYad����ԏ �43��N���ʀ�:AxF���(����4ϦUK��U��{�Ć\ש�Oc$���<��1�od
s�RM5�&ߏ6�����f�@��Ԇ �o��A#��@*���q��|���1� �EK
��-�y ���(��; S(Nc�SmkvK�n�����Q�/�l|'�����ėnW+��im6.��4���`1Z�ƛ���A�c|R��T'�<�dc)l����n��iq��:�@X���P	�z\�՘��@��<����]j� ���x��7��6ߕbv�[`Z��4n����� �������B�v4XE3��U����/
����˛ �ag@V�Ӏ�UW�����u�Ii�4c)����  �:#�v؉*�>`��� sR�;���rf;�<2�H�Oq?�St�g��/�l�yE�u�Ha'�]�ە��@8�A�+����T�6"Ոm��t�� @��B�ӹ/w4f5B?_�1/D`��Ls���ؙ�$���%�cs��ݣ�8%��uc���7K�	y<_�9�b���S���Uey^@{}9�ߵ�ї�Qo,�k��H����:vyK�+�����;�� #���&������.1ŨK�p�Y&���h���ĺ'�𬖐wLT�o�b��V�,�U��T�1/����B��9`:n&
�"}+a7ٙJf��ibjʔh#��o� �	��j�� >&V��쎬M�:B��nf�AT&8;�t@:�xA������6Q]j�w��"+���f��= Zy�ٟ�E6�̘~¸FJ����!���"��<KEI��(lg6��e��s#Oʑ(�/�ž��
�®r�Ko��Q�˥^�^w�c��fyU`�Xn�o9N�n2�Ae"����81bg�q�)�>e�@���0U���j�}A4&$f�TS�a�)Q��2أN�X®�PO�]�5�X��P%��e`(X �b���V�uf�b����|�LX�KƆ��nu5.�8H}�o(er�R��#�Ob��X�:���TR��I��u��@h����m۸7Ɵ��5M�M��a�
��7L2�Y��q�S
j2k̂$��ɫ�O$�la��'�.H�@���N�dq���{����*���Z�%��:�s���� J�w)�k�����9XI�h��?��,����?��(�BdW&�rT�P�r`�A �>�����d�Ǧ6���c�4`	�=qd;U�������� 5�,l<�ۢ_6f�hx�M `�>���|��vF���:�za2��c�X̠�50����2�%�����\㇊�Ip�R�t%co��Ԋ��(�`�+-� ��5^�j�ƇHҐ;v`�1�U =���(R��u�y"��S�,��?���3�ϋ}���������ؽ A\��_���k�\�
��ʭL5�����@ �nN����d�T"�؆��ŀ�v�K ����j��*D@et�R����'?�_�7nb�ڊ:h���"���pl`^�:烲���H���ǉm�6���!p6
{ƽ&-l�F��2+U��vuKd�`�	#��kc*3�n��(W��J�Kmb&şL�N5`��
�K��}3� ��x��vaV��AC1�h}L+b�2�U���?��0t��&��w�@z0 �t���M���S�o*�c��+���e�A$oۃ+�f�`��S�	�M���a �F�N��H1�lb5	P]<�;�;N��TU̫�6���,�ؓw0
gw��>&�'�O��M��&����!���3�ƌ�:#Z�И�k�9�j�r���#����� ��<�A6�p�b���-���Y�5��/� 3)��'��<�b{I�6��b�'툷6Y];J��e�8��D�L� x؍g�O5�otD7!Q:���&��iB恽Z��Bd0�T���X�����p��e��\�o��=�>k�^
�Evn���~�i'�5�+N ɂs"��l`���&N�Ln�C��a����KFk �EA�Z���sR-2IO�+ƾ[��վ����@|��p�D0ƄO}�l��q�giy	}+���4Gq
����)�+x氐�f��7�L��+T��=k��V�k��՚z��e��"{�u�̲��H�U�8��L��b26��,E/Z�V[�J�����ԑ-0NЩ.���Ǵ�c�%3B��'�fl����03�5Vߔ�,,�_ї�ɼ�\8�S�l�g��藍e��ĈV{��1���S.`��F
�oԸ�	���)����ph]��jjR��dr��6r�2~կ�� ج�NMM�Ǩ�k/>ѐ�'郓虡th��Y����IT"�X�诀�/���К�?M��6\+?j�#���t 9U�]����t2���
�з�}b?B��ؖY_�8~�e��q��X���c'�Sx�� ���b�?�+z�a��N�-/�0&�{���et����0�}��L5�T|۾�%N�x���;̓%�����0i�S�Q��5�
(u;Ϩ�I�l��#�+�D�]��᢭!�X��~�X�|���Iеgd@ ]�',�<�m�c�� ��l�W�"��i��Vq0qp.�7�?�6D���z��@���@�%��+�F�"i�>m?�G�_,�����-[H��KLxE ���Z�z��-�[��7%����1O����P�`lIa�Lv���N-ww��,�R����ׯ�ą��W[���ͯUl��"��D�R�z�+�bA�U3Q7R9\q�����}�L�����<|�\����f��HW���x\>�7�{���l���C�� |����J	&,KhG0\�o������ٕ��]]d�DSK' ��#z�?q4�q����8�}�
ڴ��-�}����T�@�����#��@�4�0����{���C{� ���^PD�*����YE� SW[#�0* }�Ol��X�����+���%I ��^kT���c_����o�=h�t�ۀ������g���0w�v:\a��%��k}�������,�j��>�����c���3w�<O���1�P_}&��$�̫���&b�1��I<� P�h�x�C����tA&H`B�sLA����YU��HP`Z��?/"�;����N��5V�� 5�ݭ�z���7K�4����Q�yށ}d��N��S�d���G�Q,:vXd�y�C��Tb��G]�+�j��><׼���]�د�K�E���<��B���]�b�#���l�6A�4" oQ����Z�e����b
��d�kx�4XpL�7�eyk�t�p�P�=�+>�@���vn���f:���fP���ÖQ�<^d��մ#�$���WRl�����)D{����� �N�m� �c�;�7��6y�LFś�~.`���e�wtA�!P�?c~(L�D�;��3]�)�Tk���qn���^E�k��zn������:+Ee�s��|X�f� ���\�@�XT&3iS)NU`�H�J�H5��=�>�F	�撴�V~	��\^�/)Ww�m�^x��Mt��^�(&2V�e�tc��`7�)<(Z������������O���w��w���NK)i Krٙ���Np��뒮�SC��%@Z'oӵN��1j8�L�PJ�ګAl�Bװ�������9���q�Q��b��%�R�^�@�n�T䋦�fſ�N�[��Q�C���8��G������
^�>�);���z�0I�w�IF���<��H�X��bt�S�_}��I�J�f�E�ʡ��|`�|�Y6ը�Ѽi�6��Dc6Q�]|G;��ｱ�"�5���S]���`�z������U��:�Jla����u�8�`,����0#}|(�������Ǐ��Ǐ�ݻ�I�e�����������K��c1�������+�aw�e*�:�N�
p�w��Y��ű �r�x�I�V`�~�8^��o%V��t<�R"��!b�G�Hծ�WaK�Lo��u6�T̳��#�aU��b�<���h�;뱂�X�}m�\`�Ffi�	��~o�
V@Ҥ�e,��YNl
��#WŝzyAO:2}ZaF�!��8Oc��^����~D�������W�P�^PFL�V���7G�h1��Y,y|x(���˗/Ogf�^^gf�ylt�,����O�/�RtM;b�"��z쇴���`�
��<1�Q�h�k�.�'w���'��(�[
�1vއ+��w�5�:�(�Bġ=��i�k`¡��1�L`���Ġ����N���FuҧWs���.s��գC�FO1���� #���r�:˱Ks@B?3`�&U��͋n��1��ԶK5]���:��Z�,/2���)����3�bX�$�����	�T,B������G����):��L��ȞŃ���Y{80�i ܟ���i.O����O˗ϟίϞ�ޔ��]<?
�X�,��'Ì҆{2��^����Ϲ�����X�1 jJz�I�8�DxԸ��˦��L�.Պ?���_��^�Yw�[nۦ����5np��s`N�g��g#��pa2���>#op�+(�4�LWq����S��@9���p=[?�^Dc ,R��u��6�%����Z�l�Â3M4�F�H������� ���F�`�e�
�-�$��N�>ߟ����~}W���{��ޝ����G֓�K0���~��P$I�0�|y�R��d))�W��כ�󺲏+|/�o���{�V"�����h��8���,�mɥb|5)�/��?�{<�<=}.��3f������fD�w���R2�-=�	�{������<aխ��I�`��f�Sm���(����	ȑޡ'Gc�kѵ��#�lb�ˑ��eA8G@Y'��*7R޴��tV@�/��������]��xJu^�O����h�0J�Ԇ��U��2�F$��O��X8�`7�R��#�UG�<��N����yޗ����u�O�EtQћDq��Uo kzS��s�������Z�?��p~��|�����/?���3�~�V/�Q��Њ1fi5�VVa̼���o��Q��������K��o��,�k�Ȫ���Y"�F�b���&����(b�r�O,��i�I�X��)��3�O�M٤��,�Va�[�E��h�.��/v���-I�n�@�������̐S��g��S���߼�X�z���&5nЛF�Sm���ꗻ4��=,��h8N[z��[c�@Pk�Zg��q1k`c��u���j��f�H���Kðͼ��N{�K�Ekf�:>H%����s��Z�:#o��={}o�ڀ�Pbx~=0����Qz����N�Tv��|��
 �ޑ�+$�j��<�\h~��j|��k:ˈ�[���ec�]J�\^��{���o�� S�e��w�Ow�1	��)J���:����|����.���S��"�ܰ���N�� ;�u�.Fg�p)����v	�TL��v+�l�٣{q�j�|�x�iK
Њ9]-�V]q��L�A1��6 ʾ�׏�t����5�P8���|�M��A��Z#�@kw�k�n��ʶ��l��`-)[h�}!�$����|�Usvc��Z����#% ���}9�+%&J/��>6~�9B^bi��ؑ�r���Xl��~h�������l�I�<c�]a�:Rp�x��� �u�V���Δ̡ļ��@���L�x� �������,w
������Z�����~k[/�݋ķI1���
�:3Z����HV�������|�IC���	�����N����w��T���Z'�t�:#��$���'	\��K��Teӎ��8]Ms��?w!^,L���ј�TY����g�d&����H�g})��~��'��f�ة~Y^[n�Pz{��u"�Ӈ�0��ꀯ�.΋sR$t����=' ���Z#�"|�E[ د�# �x��k�6��{)��k�0#k��1�G���V�&����x��u׀���F=�n#�됨��V��B��g)=
6�!c�9�(��Fm��ȬPu�v�c��CH �uw��DJ������3�|�� �މh��	,[��&n������oqߦ|���\u]��}�7�P�B�E�I*�k8����l���RR��_�<��3r��2�B+\���GߍV�[����-�A^V[Sd�B��1C@�Y;-e��J��6Ľz�X�EQ�J���K�i�[UȥF>ېv��ԙ=��iz�ݘ�z뮻3�]
�s�7��N���C\:����3x�;��;O�H2�g�H��O��MS� �T"��#L�ޢ|�����Xh�K�� �*Q �>��|>2���� �"6�<g���~sV;�@�g�#��E�%ߡ�*e�X�ԼH_W;��?c�|��n�&{�v��o}�pG{5�1�zQQ3���R%��^� �[VD�0稟�o�wN,rw���{��#g�{�L�4��K6��<��bT�������1�����R�����,�53��A�v#[s���u�5�ì 9'Pt��3��4�]�C �E:�G��V������w�'��/w^���o����/T���˟�߷c����;���}c�^����©�34�3Q~�,T����<��T=��0�ċ/�a�ɞ7 ^�-��O�{<�KKl�?c��i���7��q���� 4~@�o�m�2�f`�� �[��-0uf}2P�	�n�'>���K�����������Z6�c�<������T��U~�v�V|��?�{�����֗�At�3K"<1�;}'%'���,�+y�4��j��1����#�n��T���M�����	���Yd�K��a��3R���4�޳��n��16͠��1��x���{D����l�l�վ��=ՠ)\���=�}[䄅�$\��.��k�������H8�N4~{N (^ Q}�wO˹t{���1��XLZ۲�.V6J�& �=Տ箚�ӡ�q�o�b�@��z�a+m�	w�;�xg���d��d��V��#����H�#'0���F����H{��K�������v�\���u�� ��A�#�@��WL���'j�d��\_���(��u"�@U�J<у��O���\����~z{f�?o�v�|3)�w鴿r���� �3���﻿�Ʊo��62hs	�_�=�*��墊�jn�<~�K"�k7��5{���F�=,���^�ȼ�`�A�Z{8����&_O��A��"D�:��l�����u�K��u�z����/��y�����>�Tx"��S���h!M٫j��� �ob;^�[K��������M��q� ��j??w��wT�Ћԕ��3�H��||�z^�W]�o�	\���ֹ[�M��=HJ�z�Ku�ާ=���}�����+�{%`(������:������F�>L[ɠ�״#C�YO���t���9&RHF G7��z�	Yn�i������EZֺ{�K�z�x���^\d2��(o�#�I�������*����3"�g`����,Ë����Q�)c���x�q��^b��:���G�O�;C���D��'���e�u�{ĝ펯�}�����땍��� ��D��L]�i�_���@sq�]�Z�n{|������|o5z3@}��U���������o�p5��7A!�d}j�\�7��n�6CJ�g��x��bq�5p0�k�߻�rvy���;g�%��5F���"����rS�D��o�!�k"�"e ����o~ΘU�]"1��=�\��1�AB�T]�/��$�u�XVe�}���ۄb\��u{��}�gQ*_��rc҇W �,]��ۖ8���+5 B3��'��JT���ZK�����B/ׁ����
��ˠX��=�o��}��^�V��@Ò]��Y�1d���ϫ�
�� ��g�H�I�C����8� h ����='��ߚ_��s��,�Jo��u�TzpM?��A�ʛ��<<������Zf�ߦ	up�]� �����AͿ䚦9�_G'�駺ү޸!�^˝�ҳG*����.�eN�����'q,�.�{f	�g�<�Rz��ۗ�E`�s�͞�F��R�6v�T/q�o]��"_���B�\���ϼ'��uz�:g���w����c���۸P�EY�l|��`4n���6	��������iF}�gp���fX_���2j�q=]�hAڈ�N�f�a]�K�w/·
����}����W�0�m����Ok��{����W��c�ϗ:+�JI߁h\���ێ �����~����p�����D�M����z\�m� �r�+k=P��&q� ��@�ǟ�Hl׳�_f�9�m����X���IW,7��zU��t�[�_��O�T�	���O�p�j_�\Z�V�Ǥ��=}���ce �<� r/�0�sV �1�S� �{���2������ė�P�$�&Ӫ�~�o�|Q�(k@o������r=��r\'�����`�kF�ϱ��
[�' ��ͨ��/���Q�f�Ժ���V��W*6�q߃���������!T:Nw�mF�z�� ��ҭI���\,}燿�֛���ј	�uF׺��c����=z�A�ZUl���>��|�&ܲ#	�zl�s�3�?sz����F�^���沺�Yʛڑ�W��i���h��a�D[�~�I�NI���[�= ��u�{��=���5@��O�֒/��>���4Ɇk��R�Y}��ڼ.���Ձ��reQ26�֮�~��MKR��K,4g0�`�\�n���F�a��M)�㵀���b�z��&�%]��ѹ�(��nD#���D�c��o�绦'��]���r��Q�~���r�,�>D���y�b���a��s���mW4�c`Y�S��8\3D̉m"я�����w��,�{��@Q����`�-7� ��g�w�:]�k���(~T�D����G �U����ts���{�z���A��-&A~��Kf�u%~�Qu�;�() �����z[㠻1���}r��15�s���y_b�#]�7�7*��X��~"���1����)~�i+끴������%&�븆�&[
`�тF����q}����͆�����:G�%���~�ZL�1�(��l��ؾ�WcQ�(4�Z%�t��CJn���>����%����F��1@Z�j$�c�[4c�r�m�}$��Rz=��ރ�t�E�@o����&V̷�ib)�Z�DCtY��c_���6� \W5��y4n�.l�wP�c����7���55K�#�R-6���V�k�s4����6 E��@j�����ط�K��Z�2�`�uBB��^��y�v?���R��b/�m�h'�]e�%��w�5V~~�
H��z�^�.��{�]�ޗ�u&�������}��6��ۺ�������Wm!��|����s*������o,#M�'��M��p� �W�8�J)����N"�%�-��u�թg�=H^S�X�ݿ\&X�@�/���ҳ_k��A���n;�����.U+�9j��%]�
���$���ܷ�* ��k��7�r�0�y>��\�<��ّ����"��8�4y�ёX�2��k�t�[����І[��t���փ���.�hz���n-ݲ���2�����]��Z}0�os�	@M��u��Kt���/��k��O7��6����"�����2���;h+Q�5�e�`�n)�c�΋okp���V�[@t��8!	�/r��~�U�Ri|Ǜ'�K����)�a�]��7n���@�I��zᘗ ׭j�-"r���@���ko�t�6y_x�׀ӵN�N׮���^[^�[z�j�ƃ���\��}3Ϧ�����'2�[ڧgz(/j�v���z����A�&���x}Em��    IEND�B`�PK
     mdZ��� �� /   images/7b19d218-2217-455d-9a43-b73a208c2c5c.png�PNG

   IHDR   d  �   9s8�  0�iCCPICC Profile  x��||eE���6�ѫt�q�"�����ٰD�ݐd�b	!��l#[`a�.  m�"M�(E�HS�. � MP����ܙ;�w�������w��L;s���;�%ɾc�,�3��$s�-�<��Ǟ{UWz%���K6Jt���-]]	~���{,i��G�i����g����a~���a����_:`���'�}�s��Dc���!z��G��xrzS����
:�jKf����d�:�Ë&ɪ]�i�=<�2���м����3�Θ�$�A"ɬ9���>�Ɯ;����I2��E�ó�dm����}F�5k���6)�L\R��~��.Ӻ���nU�2֜�ff����[��78<4�M�$%Ӵ)KӁsY���L�M�M=Mف����n�ٻG�e�'+�iIW��d��-��N�˒f�J���֎�5��׭�Y�`2���P2�l�4�]�3�M�^�����gI�Ԯ�� T'~{\ˁs1�Y�ѶE{oR,���g�����u����C�f/��@����jM$=	�Bos��;}l���-!����b�$I�`�!������d��c��$k��$��@�y�S��������������)�9�%ɵ�m�ɓɫ��6l� vmاaY���6<��ڨ5Fe���:d�e��]����G_<��1��sژ'�n6v��+��s�wĸV�x�y+�v�MV^��C�LX�;�<Va�+�:c�?�ֹ�]���~�z����rͳ�Zk��������:����i�m����w����~a�/\�aۆ�耍����M��ț�n6c�7p�c��_L�x[�_j����O8cˁ���국��f�/o�����iv��k�}�/��u�|~�8X�Q{���Nݮ�ӷ��C;���_;�岉��>:�;�<y�]���~���t����ԍ�Zw[�}i����O���5{��k�7���ߞ�w��o���)3���f>��}���y��_����^�xs�p���]v�w�:����>��#78���s���vܣ'�w⸓.8����O;��	g����g�t�%�u���Oν���]���W^~�{������|r�S�����r�W�ܺ�����o��󮻮����N|��<<���?^���lz��g|n�秼8��^���]_�ፉo���x�����^�тO��_�?����ڕ\�|���pݨG6��3p�{�ye�A��w�J3W����*7W�^���[��5�Ys�Z�}�:����z^��>�p��&l��&{l�x�S7���W_nL���MZ���լ��ns���������=���7�x�XY���כ�-l�v[5�~�vޱ{����������^8麶;w~l�K������n�!;w�2w�q]��vo�+�+O�j�.����=��/���7_�֊���޺�}��͘3�p���3����{�~WϹ}�C���O�W]�ɢ���/����Z���c>c�%߹��������#�Q����ѳ�Y|�����q?<��.��U'^{�/N����N�|�����?9��3�8�Գ~�c�>�C�=��_��?�`���h�O�^<��/�x�֗�}E�\��U�|�Օkֽv������冎w����C7/�ղ[�����κ��;����~s�o���߽|�w�{���������~�؃?t��w���G��g���������'>�������̎��n������^���F�<�o+�����������vx}�o.}��^����<��'�����>��Ã����n���c��_���a��Fm:�Q���Yc�{����ݱ҂��]����U�d��V;~���8u��ֺb�׹g���{q���0z��7�z�6�}��7;a�K�������Ҹ�Mh�r���n��6�|�'7����[�ro�x�{��-���JfU��v|u���A�زӔ�}�e��C[O���kv���Gwy���]+_���ީ�N���{^�6f���'�����W~����ӷ��{l�&�dm3�����x��C��{�~�Ϲ{�S�^_����٢�Ż/�}�A�����:��e���{�*�m~8;���ݏ����>�S�=���w��p�9�铞;��S^:��察���>��3�;���>�чgp��~x�G���@�%}���.��%���ν��+��򰫎��q??��3����+���w\�����M�����o�ආ�+w����~��o�;w�]�]�w��Y�ιo���>0�����!��c9�ѓ�x�c�?������'yj��s����������em|~�ƾ����x�ٗ��ݯ������?.{���/~�7�x�ތ��ݿ��ƿV|�����m>��x�'�$:�%�5Lj8���Q{��{�}��1?��7��m��+����U6Z����V�r��V?s���<�K׾v��ֽ�����+�_�x�&6]��M�?S�ŭw����O8g��zh뗷�x����m�X��+��˲�ٙ�"q��Uݣ5�ؿm���cvXw�	;�u�̘����I���z�?M~�}��7��t�޹tʏ����\��	���L?b���͞��⛛|K~{J߬��?}�+n����3�����7�>�o�9��m��������?|���.^��%���_?(9x�e㿣���C�]r�I�_r��G>~�kG7�ޱ�/�k9��=~0p�ܓ�|�)�N���CO;�G�~�ǜy�Y��踳O<�sO?����~r��_x�E����G.��e?���+����ّ??���9�ڳ���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\���<���O�磟9�/�?{�s�����x�{/��i/���K_���;���?����o���Vo���޷�}��w��w�n|������~壷>��'� rX8��< �8!I&�+�jŊ��N��]e��X��I�J�s�I�����I2�KI"�a��g�ly0�j9.͹�g�G��1����Ã���צ�L?h�C'�Y<���Z�ޕv�8IF`��'�utT=`M�?���iI2p�{�14��V��@���u�5x� ��������������v`�dc����ߍW��U!pS�0�0{��_�+p|zT/^'����gԅx����xm��7z{�~o�~��ܿ�~��W�zF?�W�3&w�ok��9�v2�@���z�3��i/VJ������hq�>�[�P�Bp�OH%8�����/���� \�������p�e
Ҝ.p�j���|��n]	��Š�o��?If�����W[2%iǘ���|�|�En����&��[S�p,D�2�:�L8�=Ȁ�Au��z�c8���!O��e���7�} �s�;�5-�:��g��?�?�2�\�M#V���+i��A��"N��tm�Aw���$%30����@f$#:W������S�7i�D�� ����?�!� s?�4�@;��J�8�-��SX����e��|�I|�?o:��1� $�)sd���2���K���gA�qs������l��g��A�s�"��m��j�R��������;����2<k�9���9C��/�?���?<kpQu`v���м����������ۧ���:ch�������޶I�ƞ�E����Uf���N��$sՁFL=�����������8�����e��JO���m}��;�zzۺ�'��vv�M�n۳h� ��:z��;�v�u�uU�'O�n���tOn��k����=��mJo�q���E�ա�:	K�ӿ�kx~S�u���Ý���7���|]}�{v�aܝ��zv�6N����Ll�i�k�~��J�(�[OW[kowKGޭcZ'�6;���Z'u�j�5�eƤUkk�k��j��Z��e��2ejwgKG�^m��z���ٗ�i�q϶�����ImS�:�����abwKo��)}]S{z�'v�y���6�TİgGGD��=ugz�Si^Rm�v�����܊ί��D�ڊ�\48�z�Т�A"���k�fk��?oF5?��Ξ*�e5�Xm��a�����)�J�L����=���Y���H�A�;ZZw��!?:��)=nW~3��sw7d�������.�8�����3��z �jc3���s���]F0u������Ӷ۴6K�qjWo{'���	c���S�4�T�2eZ�Ķ�>ld����I=U�E<����og:��JOKgW�S
��n��d���I������������#��i��fZ����A?�c��V�2���'[�F�
+a�ҽ�U�jt�W���^U�ƅIU�����~�������8���R-2�YiҊ�����~�f��k�q����O�����2��~�	f��ʚf�[�O0�
Q1Qz��8(���8:���'%�JM��=����&2�9�Ei)h�V)�T���c�e�k<�R��<2Z�Hוl�����AGͳ*�]��(4�M%�2����*�)�s]iMs�Y4�q����u�r+5�`�Iiy5n�E�م�Y-�)�@g�٪�%�#�%�_������Ό��Ԡ<F�J�J��X�05e��T�B�)����U%�%�1rנ�*Nf$3T/�i%C8ľS�v�Y��̬#�J�F�-6bY�܎>K�MX�6�1�HJ�H�U��&�2l�p�4[��M-5�$*���NA�� �Ժ#��e�F���ƪ�fRn����I�2G.�R�H��
<P�C�G%�Lf��5!�$��j�x�י��5��56��@���0�)l�8�z�k��~��R�Sk+p
��Q�:��Ƥ�ր�{� ��)�T�[��^G0��$��e�TY�#f��p0ZV��dXOp�T�9��@H7�R)�F+s�u���I)@�����r�
$�tMH:�z��mKx��ž�K@�p�D�G�%���ʩ�%]C��T�
ǲ�Gs�Q6+SN�����~*���L���p�8w�9iwRA#�5f��	%�AX���K�uRKK�uk3if=�Fa���K��*\U��y��#2���"�'����&�q4�xMl�i���'~D�T���@+G�$ͬ'������ ���B�%�ZU8|,ܣ%ͬ'�/����;�m��>�"���N���a�dA�t����,U�YUX�ι�:�^��#��0�	`��FA�֕�0�j�:~(+L	��CU�q	Q��u�Dq,����p���?CGQ�h������?�>�����=PH�?C�_�?�*L���ʩE��;�:��*J���+58��Iޖ��	�LC�d/n6�FC��� \��_1�?�$U��N)"�(�4����@���#&��I]�)U�6�2�)p
P{سդ�������z��� ��
�C����{*qR�JM1�T�� �42�U�hB�TJ*t��b5,���h;0�\��Z�F���*p�Z�!�:�t�jx		,��a�`�FT`)��| �#$9bFhf���Q�ë�R��%ͬ'$ia9Eq˒$�TFp\W��a�_G�,Q��$�#�Ru怈�HS5�@)���76�R�Zҹ 2�,�R:J����4��pE���$"��(���p�_G���r��>��P����j�PX��zB�n�w��0#�8y���(�؎$�'�0��C
cB�"�R�iA3R�z�0	�o� $CZ�f̠�p�v�u�!p}�5�#݃[� �Z(|���	x�a�����G��j ,*J�d1����%!�B,a9�8�]E钬!Be��'&���2� h�LI�gD`E��Q����.8 9�([����
�Ԡ�O"e*O%� ��d:EG��e:PFX�i�s�a
���X!�F$�.}0�P�9e,��c}G�U!(kd�FƁ�C&������ܭ�#�i��)�%�j���QĎ��8 ��A�=9X�/ WS���wD<Eg9X�?	��=�ȭ�;

� ,���{���P �K��x�@*�@� Dq��<+֋l�>Y�R�g�C���	r�W �b���A`��SN���D૘+��()���@�vd)*�������� ��)���BN<YuT�Рd�Ry��Dq�jd8��)2��(J9��*3*�0#I�p�BW�,�(���)�T�j2�3G�tQ ��W��(�G,U��bV!����?C �A"�/�-wE�k�b��d�qF p�d�>0� 5����%�*V(��F�RR�wK�;�O��g� "wnX4�T��R��1+���[0��+#sQ��+p���W�@(�"ׁsd��Y�G&+��x�(@ #C^N³!X��
�W��3"��yXE�3tP��U��)����������TE���U%�R)�g�	�����
�е��=�T ,�ܣL��(��q��5 aԹGC�F���pl�{,:
�r�F�s:P�I�-�J������Pmi8a8��Sa���f%=�bIU��gR���TH�>����mZ�6��"���'��DO^�[���"�g�[����� ��(q�Q�3
v�%��(��:��eU�b`���� 	E>��C��YVG.z"�d 䒪3���u�3����w�(���Ѯ~(]-����YVK.zr��T�#+�����jmy�񫥴�CH)ὔs͚`z%+-'�@��`(�%���%�	;��e��ؓ���M�@�=m��=Y�(4�� �1�p�䝡�����KL$J�����մ(u^2@��)�T���2r`K���fN�3.d;��\�I:~$=��@�{�~��*�5z��t�S�V��9�jڧ.q�q���s��"�	U6��eSY���}�eS��)�f�)0�iKzFϔR�I �`��J�+S���@ rZ6�D�ŠU~8��L#��� -���/!o�ی��-[Pi�ϴq��2�Ig��D\���j�yY��y ���%=#A���i��Ǩ"CePڧ,�q�������T3��%
�SOU�5�& ����kAu*�Жt���U���dÆd��	dwH�H��Z=�Z�QIy*�Q0�&+���%^3���q�yBR��w*qpNz�KӘ��`S���K2��Pt��A�����OQ�_S�q�z�(iNV�M�$&H	��1
WlDO	� ��L�Qqr�Ty
��H���cJ��D�7��(�J�¸K�0�0�
=Ed�?'���4��\������`t�L%(9�qZ˭��P�3���� �!����U�'�g��g��=�}�f�P���L�H�EO[�f�����J�r���0�(sy�@���Y�t<�aj�9EV�

M��)���r=YfiNF�G�A�c��KI���I����U�HV��q�Tw�u�J'WyOn4��(K�cOzPĀ%H��H�)a��\�,���B֨W��j��J
o���Y���+�g�łzl��i�S�`���p�����e��}Ҝ��g�'��	�h
���.
�V�;r�p�6��fȊ���,3��	�
���~��C����2+�QT��/zR%�S>'Ҹ~H�����V ��* ����J	�J^�o�O���(��;�×t�R��ۢ'E�T@[2*S�(�I�"�0���#f�̸���P>MZ=DOU�3n�����:=Z�甔��2?�Isfy��V���<�8z�{R�R����K�?�ׄ��ZP}Or 1:F��q�TR��cq����A*0��W�e`��SGeR5��%�z䚹�^=�.iĞP�Y�F��SN�9�O�}~ڛ }̃7K]D�H}��J���(!��P�	 ń�"]D"l�dIt��Đg�(Rq�Q\d�V�ʒ�BfX[
���1����)\�t�����vȅQ.H�o�,�Ӕ��� ���'J�����)[�
MȨX.�#(�ڼgF�L�9�x��=�|�t=��BBz�������&�bR���a��F��q��PyM
�i��!�	I��F����pʤ���<O=	�iQr�q�����N(���)�)���Y&�
27�dqѮB7?���%C���
۳����ڭ�O�[��Mb�rÕMVm�n�y��Ӽ��c�y�u�yfF�~�mD�Ȫ��]:���EP� ���!������&z�Dw�4E�j�������.�=�o���Cs��1���s�.l�6��3�r�VYrIR�\�����$��uH����!��-�G:^�g\DR���ݓWJ:^M7��+i�Ƚ礥��@�x���8�Z�*����ע��b6�K��缔���$2c�tňx��G{�UѩOZ�	��2�-����Ll�HCT�=�����jEh1:��N�|T��2�EhE`t��������9�@��9^ZB��rFO�s[�/�uG��J@�@��Μ��;��?1��N=���%u��RbǫSzt�Zm�]x+��At����n��A� �����,�W�7;���D�I��'qX��E��}+��n
�:W#�V�zU~��x��|H�HԎ�~rAѵM/�@��٬���Đo�n�1�I�9?��x^�$�Z�6�df�r��B�疛�k�I�
z��0������9�L�d<�D��Gb�\�	"o58='��|7�e���,#_$] �����ߦ�3"�d�9��7$��V�$�~�5Г%��*52�Y�u�6�p����,_B� ���U�nЄn��x�Q䭈�~��":Jߍ*z9�SIתa�<�$��|~!��f�i�Pf<)����s��]�kuY�$N%t�����Bb�0y�I-�9�)�r^�?^�V���Ҧ*��X.3�^��`��ZA�����r�_�s��z�Z��yu~������a�s]�ru��_A�xA7a�v�㕩7H�D~�#'�)4]��ym�g��iH�Ck��Y�n2o��o��S(RɜW��H|84�TOB�r��(Z�V#�
$g~�ty]z^�_�r��MV� 	�)��&�F�DM�9'�nN�y�5�\!�N�<
��<	��K* 3HV&��|Λ�f�ji	��6���r�Z%z�@ʠ%�J���7����I
���`o�\+�_�� �K����V1(�w��/�$�c��"ZAx�J2+F��+ϋ�٠.ጵ��S9�k=/9k�j�)�u� (�t�d^��N&2?B�+���
}��a��;F:Mu���v�c�tN�:��PQ&���E� �˱��@������q/�\x���>P+saϓ�z�D��܏�è�U3��PH��IN�]�[\�g��=L��K�)q��0�g�,�"��|	�X�j��_I����\�X�\+�i�z�5{O 2�^�"��­	�2V��~��� �e�_:�˯��7�y�,d�ݵ��D��e�C���r�*@�6tC����C9�*0DAfE�������'����ޠ�{2]|��I�HH��
�L���{��/�� p Y�ܤ�j�N!�d�y��t��n2��0L���u [ɘ�![|΂yO����������0Z"���D��x��0�W��đ����0p�և[�ڛ4'o�<bfl���OhE��yC�@��Z�'��1�GC�8
��{.FW��-0�7�HN�7��Uy_�#��Ⱦ�C:������EuӬ yȬ8��a8D�'��&�V�}��d�0}7�9��1�#	���p~ǰ�=o�a�՟0���1CF��/���{�2{�~܈ahZ�Ρ�2�Z��1��7&�T|���6�WO��er�Y<���_ʲ0��>BrJB��"��xx���ӄ���[`(��a
S!i���+)��H�׳�a���%G���$6ă�D�)Y�D��8A�q#��p�ޭ�L�ԑ���[`��F�{؁��WD�i$�QyI�g�y��g>nR&�]7�����Na96+��n=o�0X:��v�]<� 恷�0Xm�r��y3�yC��T�%|�IY�1t�� �t�6�,b��=�a��>��F�\[�#$��I��ﱧ�BR�UP���h���-0��2��T��c1��[r�S�1kU1�i��R��I���1}އ$��U�5���ɽS �¹�"�z#����,���eIoC"b����Z:pR���E#$���J��] x�*"��y=�T������[`,'�E�	gA7e3�[`,�ER#汧�F�'D �O�;�֟E�0��4��U����ED�� w�n\i)�-0]m�NL�B��)��F��X��_*��AF#�_xCY�&z��-0�>�f�e����GɈa����̼��TH��AF��2���T�j_ޗȈa$2'�}���|��g2b$����&�t����0HWT*�$���1��a\��x�g�"#������0U���x��H�UэPYNbX��2b�n�R�Rg���0�"������K
�y�)�O�%9J����YDC�\�NC7�9D#	q�@j���F��
�xT��XЇ�a��yX$\E8!����1"w�- m�:�ce1��Oɛ@Zx�9��FRu1LL���I�fàՆq�����~܈a�¸D���G����d�0hաbZ�:ݤ�k��R�nP�2�𵷋�a0��A Ï(�㐊FR���`��i�3�[`��S���5ؼJ�x����JB��`��U�0��/sOʀ�1�J��-0ZC�H���С�i=o�a��m`���%�>��������-�'��W�u(�[`�����w�i�k
*bŘ�ABk��MK_�P�(�Wo�
*�}*=��511}ZW�����*b�L�+�����n��T�0���+}���	0��uZ1�E�U�;���>`�y�(�{�!z݁��>�Q�(�[�ިXx����1���?�ʐK��k�y�`AA� |�Qt���Y�0��3�a�*t=bEwȳ� |ȧ:��Q�F�9}(�=F�1�k}~���xo�ȭx�F�3�!X��Ǫ�a�e!��A�@�P�V� �����҆ڕ��ޗ�A�p��V|mEG�+}D媠}p+��a���ح�礦˙��FY�@א��R��ۦ���D�=�?71��k�{���)�C�atV$m��R+��:b
�,�&�&���ǩ:bڭwx��T���WG�黩�s�9i����a�d�^B^�C�<>��h�SAPT��"���k�x���`��l��?�À�{��X�Ky݉F#��O�#���5D�"|2K�T 9=�p��`
�Y<��O�Hn�`
��%@g��@執�a0��nE+���Iz^��FCS���B�J��a�
5��M~M��sވa0E𓚤Zu�Y:bLa}�Hw��,��5DC_�ࡄ�¹�}~�#�q�گ�(N����y7T3<���lz�c"���)'?�:���8d"�A�

Co�2C�R¸�Ak�{����5�bW�G��5T$	�E]��-�뺉�Z�Ã��89o�a���!�׀��͛�a�5���-OZ���Z=ޡ'����%��1�� a�n����/��a{5�C��X@Z_G4��W���W0o"���~oàU�:�!�/H�k�&bËg�=4T������pև(�:i"�!��^ʇ�� �L�0`Pa�z� ^7à5�>�X�¸:�L�0��Z�;��ri��Ɛ����4�<7À�P�pB*?,�[`����-��GHz��kL&b��3���6X<��g&b�{Á��C��x�D�PP!'�q5�k�&b0dv�CӰc��#�1�e� ��]<\��+11��Z!���b#o�a� ���z�J2��[`C�)�Y��z��o�0�M�c f�&�k��+ۈa,}Q^�fC}�����1P�!��.Z��f=o�a�V�<�����]�����{Ɲ3�!7����E1��a�p��`0�c�����Bɹ��l�0"!B
̛��/����0����o����(��2�����xa	��q��_o�0��*�W�����<o�a,U�Āj^�ع�b#���)��R�y%���җn�7@��Oڈa0��
2@*��5R1��uK��wA��<o�a�G%����K�d��-b�3��ᰃ�4�x�-0����n:⃔<&���%�;pt�͇qrPao�XCߐ�I�t֕�r��Xz�x���[��Iϲ��w�Z,]��֥��Rw�$�_�Q���d   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    R  �    ~  ��    x       ASCII   Screenshot�lK  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1662</exif:PixelYDimension>
         <exif:PixelXDimension>338</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
���%  ��IDATx�t�wsd�y�y�gH��+��Ֆݤ�5ÝU�P����kc���~�Մ���H턺�M�a����*
ޤϼ���yϹ@��l�@e޼����S����+
���P*�B�Z���~�F��W�e�7�y���A(����{��9����g���O��W�X̟���o��~���>�ߧ�^i?��5�S��B�\	�lƙ�%d�o6�g��nh�l?�)�Z��1��;�O)�K�VSSS�d4��תzϟ]�z�>�Կ�ݞ��h�3�U�Vt���is ��MOO�iS�F�f7⚴� n��� ��y9�p](��}����}�<!�ߧ�S@��$���{���g�~e#�$�
�7 �0.��H�,�
�������~�`3==z�������~��+������R�:�F��n���b���C�!���/���������011!��e�r���I�I �/0�����R4�q�H��S$C|��I?	� �� �kN?�n��a����䟉C lŸ�V��C��Y6��X1`7�(�L�&''�1�͚N{������VWW�~�ޥ���5��+�r�t:��>�����밷�J��������)�E���O�[B�	Ћo|�u�D- 7�H	xIL����_TB/5�6��u�^�V71��tO�r
�)���d�9���~��E���咉Y�nǈuR�?<<�s�./���NDv&��B���?����WXYY̝МX��T� ���o�����mX_ꍉ�{�)�N��,�Ά��#-�an�ۡ�j@P��diE3
���=�W��"�������u:m�=a��j��ʟ����gÈ���#�FNC ���j-�f���Pww����01Y�Ŝ�qb����P0j�2 p�߱��0$�H��)[/ϫ�R�+:�����0�����f�ik���?�1\�r5�������&�`���q\� ����ógk�Љ0k�<cn��c������B��Yϔd��k�F=��Q2��UJ\����QR�6@� F�L���]1��!���Y#����O��wR"grr*,//��㣰�jSԉ�  	�����ܬ��3��a~~^����ֵsssZ�ٳg��Wv��p X��:��⚙[�v�����OLN������%{o�^��3�������i��8(9Q q�X�~�
�� �`�K�+aqqQTztd�l�=�1 i~vND���?ί��77eI�9�`@r���0ʘ���כ�,�k�	 �~m�� ��� З�����W�k�%��`����S[�Rx��w� <Ar?� Y���W��UX{�,|�����\������Ξ]5.�gm}�Ν[[���Ja��>��}+R�U��>:�$�j�8��Xgݮ�+�bq�5�Z-��5�ɥ7�h����,�P�h�����t���-!�ڨj!+&
�X����]����e�ՍZV@=�i��6����ٙ���m��SS�09?a�Z�1D0(����`��0$��f�Z-k�z��Q�+Q��o�fC?++g� �}6��jќ�p�bx�b]߁8X���C�g2�1B���e��ph�8bтtK
s���"�ܬ�D�C�"8�u�)�)�@�:��Dٌ�鴻:_g�ͩɦ )��{X,20�t�ʕЙ��A/_�4��� P�RG�j�ڂ��07LO7��W._�s�!#[ό���߻'N��_�ҷ/��e��@��@�Hy��D�Q�3��%��M�A��lƲdO�$����K����@뜰�1QeE���A�:��b��:�����G����¢�uh��m��)�3rH�N�6P���h��"�c<y�D�2�ƀ�	0�˻�����A�о��vwvEm��R�[�ˍ�F��[3q�L�mr��7��3�+1b�C�Ǧ�^oJ1vQCq�H�����a�D"��GY�9��M����2{S�s�("�gH1 *������ϟ��7V\6�5�+u��ã�8*9��a_�Al����C7!]�OfL2�6��$�rg6wj�Ȃ�QPX	���Š��h_��W�dY�6��Xל[]�&����E�>�{e�?�7����^�a�(JL���-]�rL@Ƥ�z�Ϣ%M����ɓ���o�#�C�j�b׈��7r-�n��S&��-,�cqQ���gl�:�b���P�錾E�a���Ǿ�D<a�E 3����~s�U�HD4j�.���E�h��b�0��c^3���c76��Lb>�'���x��^���KN���M����ٰo� �����p�r��2 @be<c��#����� ��!�5��{��ލ��#}�XA�E�,'b�bn�P����f�l�1eg<wg�C`D�d��j��dW�BxDw:]�^|�����ƾ����.�9��"I��8��(��R�i��UbMڗa1��E�L�C�\�����}���h ��(��-8���|�p��w �=!?�b�`l��ŋ���Ʉ����1����_H!��$&�PD�DKt��P����r�x
ݬ�?����qʚVWW%����{��T Q �{���80��̭Ȋ2�ʞy`�#��H��~i���G#ʰI�r�*�O�l���MmЧ�3Ƃ!k��sm���3�g��`߃��������08;3z�q(�cf Ϝ0�xl���jz��ޮ �?!��e q)AkkϤO�Pj�G}��w���� pNj�K�.�	�������YKY!{�H@���5t�!��� J��`�ez`b���`��/A"V���q�GI&2:���.�ƒ�p	�� brS�d3�(�y �OX�iJ�e
�������ϝ%q����lCnV.��I�;4��,LΠq�r�<t���Q,�g���eYNl���=C�ŋ�Ddw�����gr_8�G��Qs� ���/��3�_�M(��!���(�Ơ":����n����s�$���'��)���x�k����p�K����{* �������w���h!����s�9Q$�B$�1�L�υ)�tɼ)K6��ƽ�Y +����y��C�� ,./���1ſ��J���1q�%l�b/x.z����B$pHh�H�8�q���Dt�,�D�"Q�T��{���B�z�߉!"�L/�O,�Z�,�@��.y�?ZZ��*a	�ƴ�<��ttӁ�� �,$�������_w�i ET���&�/L�`�/��(Ul�ݚ��Zqy
U�]8E�nH���[�1�`���H����(Ii��M�㔮w"z�2x�������x��������I�H����0	 �v���H2��Q����\0Q��)�(�s
)�hp���&�� �3uD,��ˤPA��������r��u��{z����}���ׯ�� �r��S��a�`SljwoO��XGW��]4�����l���d_�<���ϠT7�l��L,�o�N����t�3Q��YB�m�����\ r�&�TAӐ�.��س���MU�ݴ���D� e ɻT����!�zt���b����Ƒ�]�b�|]�|A��������u�`(�n�t�6�����(����e |���)�eCʖ�ݿ��_�����bc#� �#�|��~O�êa[1y6�x���ل: vJ�7V���7�x×2qH�B/ ;�r�V�S��S��ו���X�>l�3A���W5�`�X��B��3%���I65�ӦW)�!0M��6ͺB���X��9x��[)�nO���gW��^
?��Q�X�n�;$ipCr(�8�=N�t岛��cPHx��<z�8�5~ ��$�*�ΐ�:�N�.�5O�<Ud�?�+N6cV�K�Ք�ȩJi����N���J�ŀ{,�T�G`��XX���!E������D�8%��5<��(��H�&�*7G_���2��{ ˈ�@�������;�H6����p��j�z����)d1g�Čm��O��e�t~�嗹8@�H�Oz����ښ8�?�P��K%z��@*I���eC����w�
8k�FM���	�_��ڂ�x�5��@ �p=y�+DI�xۈ��K<}��!`#�X+�4��-�6I��l����D�֑�!璲�[1%�A�Ŝ�HČ[�r��]���0k@^4j�׀��W�j �]]=gb�g��L�	��u,��s�w(��u�]������s
@b�o��:><R����T�]�8��hbṉ��m���Ŭ!{w7��XWL?�2R�E3n
� ��k�{ ��UWܕŸ�ҭ�,G��z�tL��5�Y5�Ƌ��I)i��zAN�1+g{�#pW�������$�5`@aq���B'�޾<Վ�)��Ƥ<�ho:e����O��ggf�u�m,��|E\� �]s�3�!d����=یQ�){�7�|�{  � �?�DA,�'�=�h2����%��#���BO��Ϟ]�ߵzU2ߨ�dԵkW÷�~k�~G:T{@�,�7
�q�L"�9y��.��?#�x/,M����v횸B�h��ȓp��'"�D��/(��ܒ�үU��Z,R���]�.Y����Ʊ|<����{f�C�����+�VM��^"�h�MJ�"�-S���p�ٳ��" ��Ec��/Dg�8EؿX1e�J�Ư�5���8��4�UP��@%J}��n�� ��I]��d#V��!Y6�67?k"�%��������Q`R�O�sh끈��1���^�0�-(j��޸�4-	�T���_O��ˀxy��P�Ke�M��cC��ޮ����f��@�x�$u<��Ő z��LT�����pw?RaP��!�Z��e���Y:���sCI�&�R7����@��e�2f2�DWa�% {}�e,��������JWd �D")0(X+�Y>�������X{���ck��� �1f���ʣ�f�cEL��ɋ<��گ�(���c�π�պ�f(ׅ�}U� �ub�����2

� 7Wb8RXY���3a�LU�ب���0<��6��#2;	A(\���Wo�sAf�YT+f^�}��P�ô�P�+׺LkއS ^�d��Yu��<�Z��Y1|eģ5JAx�Ϟ>�5�6L|c� �@ �f"����ѣ�yб������7��R!^�4��1ȅ�L��(%���P��c:�X�B��F��g{�,,��MG�c�� �T�K��"ڠ����?�x'�4 #U�4F�`ld� e�LW=~�<\0����+F"� z.2��p����k�E�#7���|���-"$� 0�B�R�2���
q:�o�\�����Q[�	D�	��p����!��0����N���!)�U�ߊY�dM�8�9d��Ҋg 톄7X��{���
`!RH��H�1^�����>�j�&i�7�k�������pG����3/󩅚Yep�Д����O�<����(#�4d!R=߰'�� a8�d���+�ޚ�2 ��@2/[:*���AĀ� �˗.�[�nI
�{�%��r<��>N�
"�(�sf���+Ix(�!��Mq! xt�6`x�m{g[����-�E�"2`�w�}W���=��5B,袉R�Ħ�l�y�jǳ~��OHRa2�R-��H��s_h���:�����#J�&J�HfOG �PD-Nݵ�W�����H��� ��z���e�bأ%"-��d�nˊ�rѪ�G�7"���R�0���F|��*̟rH!�����.������h�����X�X���� d`�ݸqS���������!F)$��6v,DVc�'���b3":]����Ѩ�b+���2�����^�m�^S΂��D,\���w� >6�w�}'��B5˧�22��
n��z�psRD�j�{�b������@@O�bs��'	P�R�!Q�S��.�X��R�h�����9�T�X�5$�q��}��1J�8�F�Ǩ���G2Ѡd�T�}��X�Q�= &&k��G��҄u1��P���}/s��Hr�o+�b�ā�j��8�F�(��b�E�$��.6��|��P�v�����ޫq ;y�	$𣠡qg�I���>��t�B���T��_�Q����X�������ǥ����ū�	��%3Y=�'>��]�R�����_� �@۹s���s�6o�T�/%eH�"J�ݿ+'%�#JWl��(D����vd��Km�X|`��j�����w�M�`T{<�ᡂ�k֍�c�T��\�{��h����zݣ�OMD^�v[�=�2e"�{�QE�7��:���y��I7��6{O�r�1�bVN��%�ć�t���1*Cda��(Q��1�#P7�q�LS�>n���<u6�|�Y�w�(�[
��X�[�u����,��=�>�=���S�(�k `tÉ�2���B�qN�)7q�rp�g�cA��TP�QĞ?�補�	�����ML�{+�W�R],T�%N�.r������S/�%eBOv�h8g�ɻy�fx�b]I|�(�#9%ĮG�<� DGt������t)?��'J|<��#�<Q�� ����zD ��Y)w��7���)w�F������ˉ-K�#�@�W6z?�!^��Ck/�ߐ�T����q�'�t��d�\ �_mz��@"\�r]�Wq1Ux�;R_�g�^��y�h�0H�-���w0�"���%Ʀ�-���;,��SF�ޑ)}Ҳ'���Q1���|���TI��rB�������� ���f����u�xp
?��Se�؄C��͉YY�hø�\�3�����EW{"��W�D8_om��񒥆����Yqׄփ����´��x���O��B�{�cx�S�X�`�'8m�K� ����v�PJj��E�.R(��/c�lQ�gg�z�@�A�b�����fdy�Q���q\�~����d!&���s ޻ﾧr~��ߛQA�c@�e�M�+D}��+��;���N�3��dBW�#ѓDxa��?_�|�Mx���M,�#T�Djq����� ��(���5Ǵ���Id��Hj��B����f�&馈����T3�D���3��8[����?w�lTjn�C9�CU�{>ً�r z\���#�G*P�-����tbRU�/_�
��V�������&|%�NGQ%�ٟ��#�<8�H0@e�V���.b
uC ��>x>��3�q%JG��olo��X�F�rl��dN�lI�g�I����	Q�*�]�ES\P,��`���J?D��P�
��x�I_�&o�>!Ԡt��LSj|ɿ��hK_�z.Y38B�C�������ڱ��.�
  �?7�w̪��?��v�Y#���ס9�O�?>�jt�fjo�X����r.����� vMm�SƄQAo�O�,����O�)��?�ڌ���W���i����H��/#JB�=W��6M�M*�5���֒:�����r1:K��%�SV�΢����~%R��$�}�o���V/t��p��=����wE�� �IG��B�^>k[���H��= �{]X=���T}��f�C����*�΄��n(�L����C����+.���Q��hP��!d� ���%"�U#�%C>ݦqcoߌ�I���q��s��l4�" ZLo��H���2?djrB�����U5���TT8��{Ks�p��m�	#ْ���M8傽�3�'��=�,PP�[険��w���r���I[��8 ���H�TE���#Q噅��2@�H�*�?���Z��pbꦊG���gR|A"}��;�U`��8�g�;Jm�ʭ�P�X��1�:|#"J��؈x�dA�ʿ僈!�r��b�I!�+F�w��� ��d*> �HE��۷r��T��*�r����\��萡�+Y��)@PӾ����x��X~���S"�gYA�yA��3y�y�@Fg���LZ����,Cn(���GO"烅V�޵Z���hi�;>'>�A�����z��I��T�ԿFH�tM�G9_�rM����J,n�➒L�8��/�J���ã	!����s����W�U���)"���ɘ�������r[[{.���������6+f*|��w��Ç�m������M���s������bu�B冐A�{+oa��B��	㪙��"���L�U!4C�[�-����aoǬ�U3��M�-I�:�AT*kV'�ًu��jF<��������eEIE���Μ��(vI�L4�S����&�$��H!�RqT��7 MNM��:&��k����g�^G����r *b�
���W��p�7�p�bf�����y�и휙��aŵ�弊^�����cؚq�@4ܥ�E=�9���g�h�x��wLy�ߢ����:����+�/U+�L���5�^�������"K�Fu�9 g�6@L�1!��\�!��,�;�߿��p[[[�L�`P��U@qP�-"��bY֏�v�#�$B٘�7nݔ���_��/!����#Y3�ؖ�%��
�Lfnl�D��;ъ����
@z����j.��~Ĺ}��i��&�fz�15-qI] �8��&8��SQ]��J�L�]�jI���Q�s���(J���k
�ye�RX{�L50�p�����)�c,�P,g��	�"T�@��%�+���+����f��wR�B���y�?ܹ#�q���\>S^'j���&"�h�����Ϗ�5E�!r�\C4$�����1��YT���!�b��>���#lˏ�a�0�ҙ,7���nGa���Ԕ��` Һ��H��S��'��|���z��5��N?ִ��˞:���ce�"
(�&s��>+A�Al/�#�<�b��(z�0*�\����٭���?|����2��7��*Y��pL��typڤ�jeh)J^j=:l�b��]ZxN��2q�}��z���o�����H2����x��CҼp����b���O��Չ� ������R�������I��I�r��Tyr�[
x�;xB��k����OA���b�O>�Ĩ��p��u��(P�Fg�D�ɗ\�b�v�P^�G~�N4�czF�G�j�M:	 *�H1_��4�,.�WR��<z���R�q�Ç���Ad�?�`̺�8jѡň����6<1�J�n[�ƍ�Ѿ$ �;����H�I�.@�"â�p=\B<o�,����Dc��'��X��@A �
ѥ���ѽ�B��L&,2���ԧ�������+	Z�/�R���hـw����( �䱟=}�����eq��/������'&g$ǹ'b�Pz�.Z�9NQkQ�E�<|�P��ԟK�.+�8E���A��˯����
AU�(����BS/��NʎHNI��A�P7�%kĶ"�J�?�I��[�J �pq��333!���mI�d
�	kC��� ~`w�'��Y&^�O]o&G6O�u�3:
 �!V0��M��#ߝ�J/x%�[Gp)�g %���eh��l'GB=��KsZ�@�"
y�˵���^�8z�6�ݱ�!���ǚ�s��qP;�x��q(�)I�!�����e};�44g�]�iґ��*�y����@�{�~^k�RWa�'e�K�JD�;t!�6Y����8������	.*��� 9�օ�����VN
�"�}�QQ9l�D�jiy^�QG@Y�\&:�/���96nE<��S��!�Ì9�ݖ���ޖ�C�M��J��I�F6�ĲW/�v_LU��a4�׃��MJdU���M�x����|-��
}�؎�y�DH�V�>SЛ='��(�K�/y�=�_�cE2Q���ߪ���䓏?�"�(�ʎ���A(�`��Ca@�tsFE���Z�{��8�MD�Sy���'^v�(~>l��Y���*�O�Z����ѡO������JŔg�&�9�p��+揠�[��2jF��"#1���g��(."��v2an�De�hp���2���ئS��8ZY�-:�'RX ��։�X�a�%�"r������TgE��ֆBț���z�-�6^��*LO3J2=[Gc`�Ox
�M��M*�*�^P柾�ڋ��fOj�AȅX�eD��ҀR=cb1����s�@���\ژTE��	�I��Yo(y�v"��3��.��|��ɔC������U��J����{&i��ΈMɑ���i^ӊ�B�� �а�+Z�X����~�3�>��h1T�B><�/��R KE)BMlB��o;;:n�H�6}q��E)O�$��E�G2��3c�װ!��Ԅ��G1y�M[�B!�-s_��p����5��n1��*���
8���* ��F�0H�b�c�$�I���F5{9>��$B
c9wӱ��ۦ�ѯ��W&��P�����J�P�=e*�=�{�*�9��)Ku!F\B)l ��-u�h.z��A����7d�C�=V�4���0������vh*��b��V�����0�1��o�'$�pf�4��խ�@t%�	iJ�f��f���V�9�N���3�s�\h��]��a�P%�/�z�/i�نX��(ℱG�Dl���U'E���KW�h��e����X��T�Q��]Y�,���/?R�Bg�Q��w�F�[����,�'�H�8���g�,}��>K��3K._��� �C�c�����0�޻']	@h4�厬��ޚN!�Z�j�8�m3���8����'C6��"��cxɞ����l�5&�94�'(��a"�X�y�J�(�Z-����+2#Sʕ�ǭ�7U
�l�+>��Sq���H���j�F����)q�][�1g�>�π���> �J�k�u��US��35%�����I�;��`�bQ����4J�,:��pp%ZTT!..-(��g`���l�����d�1'Ί�
�e�����K�F���?��Z�v����Ӏ�<�82s� >P�^e�pǮm�X!fBP��IsCP���s�Hi�D���Q�yy�l `�j�WRwE	?���L����xaVR���$b �!��
����}�ԇ2�pGj���X(*.��l֮����Q�s,�Z��p�!,7D��-������i�sR-�<��(W����*�jiK#X	�1��zd3�ǿ�7���B�tE�ñ#kH�L���Ϥ��uT����\�?ڱɾcA 淿�'��aq8	dAu<�I�CC׎$>��oK�cU��{q��ݝ~�)��n8����pfA�Z�����xޚF4�����MD�[	�}�Ǵ��:�M�Q�A�6����y�����O�Q���)F�B��{R��9ߞ)�#S�d��)��u�F%��=�{�u���[�5�F�� ��]�}��L?ͪ5��Gm��
IB~���W�\���3/�S�rET�C�X6}`��*��&� �h�?�P TH����s���� ����Uc�(�k=z$���4�!!N(�E��B�y�U��łە������]q?�E��"�����C����J��1�bx^�p �	j��lo(@|�cB����i�F�(K�y�&��q�QO�<��ȿ�Z�Qi�du�PP,}��+"�iL���Q��%�B���� QXV*Q�y���dA���/�I�e�_}���L5�wx ���j'9F�3�ڝG�P����1��7a0��f)#�'�B��ʅ�*�1�Ǳ��D)S�CU9s�ٻﾣ�A�^��~��˚!���/�["LB�͸��0��^��W��Z��X��U8yi�SzR�h��P&��}܁����#q4Ā��Nk����f¥�F�%t�X�P܇,K�PDq�q<�WV�b4�yp1kR��!��ycM��H\�,+S�
���3g���\�b��TKh����= �7�-���A>Hy�6~^�����1�k�9T�8�����' ����Y��hB�A��@,��Ԑɂ�L�g�F(j$��lM���pN[5�Q�io]ʝ�-�N�M�0"�w�;�@�d��i߈����K�0� 0���58��ѯ�`�p�H�vQ��z,�%x��B@l�Ƒ��Գ@������/�@/BK�jP�m1A�~���0���d⺷�z[���G*~�=�Bg<� �AD����\ȕ�`T���u!���R���o߾>��SQ(���i�4��z���=��+g�63r"#�ܚwo���{���3%�: 8�0��*��_��93K^}ЦF�}zC�e�<+(֏`�E��I�t����1Z�����ű���5�j�ƕ?.����U��(C2vs�q��(ޭ���8oP�LL$	x�i"�Xp�������ˍ)������S����,�&��JP�:?pg��aȜE��4gC�`=3/�C��^@����bD/�i�i�ٺ���� �k�n(�"��\�\�;zr�TFU��e�ʍ�����v1BlG���B��Vy�K��z(
�9���>z�O|��pc��>�ţ�U�a�g\oq/�mE�m���7�:5`�ؓ��0���ſU2�����N�eL��sG�3D�����6ۓ�T��h䳳��LWyթ�/�#��s@jr�j�>qʱ���E�В�`��R�tAȋ@hj���RG\Y)J&+�������r��Q�$o4�$���� R����DJ<�2��ը q�@��"�1�S��r�L�K�W�Q|��?�I��4U:�Ue�w~�14�G�=I�b�C (e�P����a���?|[<$�����|�b�k��>�k���Y���I���j�&��wzw��y�Sِ�7c$�G�z���.�p~5Z^�s������*�]>D�,����z��P_�/l23=+dj\�!jSs��xY�#��)���8�]� �\U��}zvvU�����3����b��s��hA#��3�\DS?�WK���&]+��<�	Y,*�i��e�a  J�AP6{ �a�%��P*[&���TOhfva6���1�O��4�u�^�)����q!�hT�1Wa����g������p�#"l#i@> �~�g��|d�j��J�Q��\���iq�w�NH�a>b�oۂ)����4c qQ�;��ߛ�p �H��y*�0ġSh�D$lL �`? `߸y���Uש1��B)�m�4��n�{~(A�S��J:ڢ��Ou�Yb��4;;��ý(V��e�*���A�D���{�נ0
�yr��x�x�
��3\.�Í�>���5��'_���d����w��T#R� bP�*���b�C��< ƍ7L�����h�`�|�����8�z�d2�  �Q��)���]'[bޖd�]{��y!��'�����嫗��Ֆ,$5��y�����a�`���Ռf7߹C"륒]�s �R$�u��Q�)���������<l����\�hn�����[�n��?�\�M�	P`wOx���SH�P �ԨQ @�ģ���NÛ��x�(a�=�6�����D�:�*.q����J;�~�0J5c(b͕��$o�����A��-?���<�y�ܓ�Ha^ӄ8C�`�!eɊ�Ќ:<9\��h��"�4v6��U�:�<���z��a���23Ow�ÇO���T���ޡQ�9[k/L��4����K2q��³�k����3
�=;~&ca1Nz����$v4��ņ�$�p�L�=�����N���-�V|iׅ�����/�_I�<��X�|f~Q�|��a.[r,ød�~V�`?�rfn!/��v��j4z��Κ"\gx?ʤ����C���R��GD�K�$ON�5X�`�P�"�yxpO���޶tWC������Q�"Q.�$	�r��=y�����~���ݻ�@X=>j��k�B��{��#Ǆ��8IgRqTC��GSS��~�v9z:0�By�<���- {��mQ>�W��!lv��`�"Y1$WT��b݇�5��jΆ��������sa�9gD���:�ɸ"�����t4�4hmjʇ�������``;0�a�P!x��\�=a��C"���1X� �B��o�Bsg{ꔶ���
eK�Gvɒ�� !�b����ƱTr_~�:�g0��7r	��~��X�.�t�e2y��7oi�o�\�Q4_�D!���[�ҵ���9#Y&A�7�v miq��0���X�@��ڔu�Ӳt�&��x�`O�EW�NL@]41��)CGz>��(�ux8��HB>R��ߥI��h���Q�<u妘V��6���"��F��%�VUD��~�d}�8eƳX���W��L�Q��Sؚ�At��������`�*3@[֢�ݞFq��+��u�/�E��ܗ��Ȅ�1c�-Y6:�������Xքc��	=#{!����#\�^JS�T%C����]M�M���[~@M�0�����;���V�%��7�L)�S99<���L���@�XR��;���Bɦ����|�A[��Q�\��9���Dhzgr�01k:^iG�=���x�Ǡ`�P�ѡ�� ��ǀx��w���T�����9d4f5ҸG��͏��{cS�;O(��+�`Y��V�4O����gC(X�.I�����Ayhɱ�bq䇎����x��^��1��o"�ϖ��Y�*>L>�1
�4U�"�;B� 24 ؔ5Vu����!Oȸw��Nh�k������]9O�uA� 0/��0��'up �"�Y٫��� �	{<7��C)dv'+.���Y/���4��c���vm?8�H�t0�����Xlǖ>��y�R���I)�Pd9�DN��3��rL�#V��r�>=�2�yr>�	c���"%5`&�0����#�Hڰ`"����ȡ��2��Y�:�̀퓪_���L��P����߹s���R�a���3��5�\���T37Q	F��K���:̧���='�h������9�_1�#�w{�n�0%E��^>�3���}/]��[��9?A��{��2(KQG�9���(�@�<~�T�C/bb&���[��AU)IW0��Y�@' L?��}�̄D�'�#��}���Ԩ/�ͫA��qp��#}����ȿ�T��|˴k�(N�rc"�1X
v��ɫN���c�'p�_�/Ao����G��a�H7����2��8�J9?��Q�	;i��B���·���_�E�2B�H iZ���6����o���A�5�ׯ��vO�_��FT$g��L�p �I,Ϧ���!L��A�O�
W�>N��pxO�Z/o��P�� �F�ii�qx%'L8Χ5���p p�`X���'�X/�x:t?���{��r~Iz�n���R�䔟~�g�"3�6�^29>�G����a�c!�M��F�?x�
By��?�y�K�ǁ��X�R~���R�y���˯�T��Vg0B6�&5�U"{!M�Nsx9֔F�G���c"1�:�d����8�1�)��S��NU!?� ���S���SMS~:�-�C�Lj��������R/���xz��v�X5�MO�a�������3��Xa������J���n{˰=+�@�z1�����/r ���Q:�s�Oq�r���顯��&$ܔ�}xt�<ap���?�R��N�1d4b4Vj��,�a���)�F �Þ���:\�S 8����<�A<��{ 7|*�w�Y$pX��U������U��f�g�!��P�S��H��̀�sr��U񒦶!�YF q嶩�hö�+T�h���v?I�N�pbc �GKL늵aXP�����s�J�I�����c��C�?d�'O?0q��|M�|Ճ����d����3�ʘz#,.W.X�M2��y�t,Sb;{�a*�X1��A���'��x&�;H�������?RN�߃߈bge|��VE�`��&�������Z^@���?�ՕN�
	:"v�C|?����������c{�
j�
�Ӝ.�:���������T�r��m��i�.!? ��K�t8����å�#M)�������ё�70�	��~��89uR����[��R%%���$��Ѵ�hz�j�B���+O�%����n���$�o{����/��WR��ߎ��7oݒ��NH�JfN#�t�$�r��K�Q�ra`>��GAy�ss
�4��4yl�(G�r-Er���?����41���KG�a�<%%y�5)]�F,󉥘�XJ?��bkT����F��׏?Ϯ��f�9�����4�f�b�!jw3%^SFo&�C���Ek�ǀ1ỹ���31gY �=^ɂ�j:Δ�	 �0v��e�nD���Y&k|`ʟ�S�e+�1��O{ÚJ"Q�{+~�-�
�!�q,�k~*VP�U���`�L�L�C�/_��s��D~�L%�}@AԽ�^~v��O��\&{�'���i�;�7��W���߰�|.�7~�DE#)2��6 �Q?��:ܤ`AB*W�6�Ή�(��yP)�Ks��-�U���@b6��0�W�����	\�\7$�p�G���Tl{f����9�i����7��A׏���b0���P�eË�C��^�����(՜�a~���@����� e�NF�u0�~X�G�?1鐟t(�8���Q��U���μ�˽t�3qg�^l�����TBa�;5�m�"j�%� R	E}��ǲH�S�~=/�q,#E������8r�D���^I�8WDی�0����d�r;���z�98�x�����hu�ǝh@܉x#���<��u$���oR�kv����d������s���^-W�Ir�=�6�V��'O�1%5��_���i�h?Ü���
���*��8�x�l���.d� ��C�
����|	��9Vẃ󈬧�&*R:�Dʁ�f/���f�2(��fǄ�A���?k{B48�ٳ�Ⲇq����T�� 3�DME�o4��/<ΨH�c ~�<���ݽ#C� n���X?z S����t�	���z���d�CRo7l�؅^�We���(��ŘΞ�P
T�"�X+P�~��%�^�B�FGS�0>��o�FPp_bY���U\T.������l�i�='�|"6�<�P��JU+�#'��7p�䴧�u�Y�.ʥ��}C��g�D$�I�҉��$�`�v"�8 X�[�q�z1"������o��N���*B�0�{.N��L��#�V�8��T���({���  Ԟ��1K)��3D޿�,(s��^��)�D���T£�F��5B��� �HB�l�/�����|j��`
�D��~I�ȍlr#�-�#}��cn�]�N��ў����Q���:��@~�Έ�ڦV���n�{Ko��F;��{�I�+1!6�ӄC�횕�0Hj�X�Œ�`��cJr�v)s��m���Ac��	�Z���`�n�%G��'�Fo� 	�8z�*|8��u��Y�L�I�r���Ǵ������n��3�AF:�7/x��j�Rz]/��{��z ��(i�NU�&]�9'~��A�!�?ͅ䓭s�����T��ls����id7"��A���ʆ���~�sE��w�����s�U�8G�ٓ��p�N{6�����#&�MEi�4G�a�l��i��P{�(�<G�cn��M�t �A��1b��p�}�`Nr`Oj���=2���^Ҝȁ��1��)��,�oU�R�;qoD}��:�t�>����_f��6v6�0<�	����7A@
����Q��)������ |��Е�*:w~2�kYG�����)�y#���������� �(�ſ��d�%�)�~�#�Z����\��9�ju�8�����o�ƳY/���|V��G����*�Y�(���X�u�.Sh��;��")U���b�ח�>l��
x�x��Ԓm�
��!#{�Yu��*��!
��~���o����w:���L�V������Yq ��  dAi�8�l#׽�!o�������������[Y���,�Ap�t*�=�HM����:MhM��i̘��ׯ��QV'A�t�EE������Ux)�gi�n���K'�3�����,�L�l�'�����R^3�.�YN|��产X�U���O�P5�)���R��F(AI���U�Ky�$�w��1�h;m�`�zs�%�l�r�TH+�[@#�ѩ8�s=K2>���CP��G����ى[��􅘯\�����T���*f�uF�?zC3���|��ION1y6�5��Mg��<>,���}�
?,ޝ��w@�g�8y��������+�%����YB�B!XU�`�Tپ!�L���y0�jp���� M��B�f >�֞(�%v��cDi�)�`�#ǳ2;�i��~�� W������,̫7��ZP� �}�]�O�o,Do����G�������@X��p��e!L�.GbLD�F�{��ώ��4�%��B�����?�3f)�I�����.�) ? �#�P@��l��Z�"?O�# �CR���~(�&[�[�؎�~�I�w^�R&W��@�Cy��{�)�݋S��t��ťF�#��P�[:�w Q��P?8����k�zQ}#D��1������>����<��eᐂqJJ�<�0Z�7(�7Gj�
&;�o���,�L�6�����-{�3��+h��O��;ԧ���H ���7Z%�V=�0uƹ]��� I	�X|�{�u�D�#`&7�C ��/�&�?�����Q��@�B<z{�w�[f 5�W�&���)l*�&���ܐ&�AD���ܑ��d" ����P|#t�r)�W�@�g�����G~���J��:�M��Ea�����hQ-i�-�IS$�rZI�$"��������*I�Є=i�TO�,���9l�D�f������^&� 0���j�*��<�vz!5H�0f�ъT@��Z���r�b�@�u��=�������C~V	H�fv�ƊTވ'��{~w͞�qD{u��B �*�;^^�d��œ�3,^Gvs~��M:[ӡ���$��y�I����P����t��g����1�I�BFt�)p*1�T��_�3ߗcE=D��4�u�rz�W4�#'���=�>�ݩs�Q��v�1P^|ǐ5F�P�L�Z[��y �k�X�gWW��~����{�jMc��,Oҏ���?���A�):�Ͼw��۪�e�I(Dh9�A.C��8^��0n��Y��W� �o���$��cM��Py^ޑՋ����|�������@J�| �G��{ò�WE?G��C<��Z��q{G1K�6���>Q�/>�����Y��h����Lr,>�6�i4���ӜR���y,(y���FmPoYJv�d!�
%���z���lqO�=�hb�r���{N�D�QJ"��Ǎ���$� b��$�.Fc*��׿�g���YX9\����Y�x8�⃨�an6�.AߨG������-�˷�&Ș�;�4U�|�.XYݘ�1;�(�f$�^O�x~�7ި��b]���it��y�:5 �kg�[�H�ˏԟ�|�mx&��i(M�4�H�š/<=[���j	�OD$��b�,b�q@��)zP �m��;�}-$�Vn�h�i<ՌǡuOM���W�]�x�qM	�
4�Y��>D����pp�uV�X��v�C?Sf������h:�4N�\��s�7S.F%B��=l�ZZ�8S��G
�`a*�)E�(� �gŚa1n�����{���E#�UI>c�a�2R�e�Y��UJᓏ?`��{��с�϶������~���O�̝�S	�ah칭����F�G��a܉"&��J^�]����q ���B�����k~��Ο_� �ơ3���8G%q\�O*T�GG"zLw�����~B� k�Yb׮�ɳ��x���a=0C�s0�0�P�n\�L�<[͈����D]�S�pv(���F�`-�e���譲2DN��P<Wa{��O����.�W��r�"s�ΔjB��C"
��8�:Ey�ǈ��ٺ>���q�{G$s�Y�߃8e�4��mm�l�D3�	9��\	��$�f��w��H�����OM�N�#(��I6���iE��ڲ��H�_KD�B2<g�QG��^>�EG�&b�����8ٳSt����-�i��9Xk,��0����7�n����kEg/���B|�����p5��S���r����%��|�ng7���ۨ�g��#�Ux"�����F�0�6<x�bC+�2�A�#�_���S��|�b�x���k/����9�>���R�����Ţ!؍#�Ҍu�?]�($R�L4�J��S�8/��,�Z������~^�&�jN��+E��Ғ�Gd`k�O�a����:�e�
Q���N�P߽q&2�M:e'�!�"�E�d��}�3�8)��ޒ؄�1�iO�@�� ��}���j#����A��2�ʊ�f!�|�Ӥq�x��cM�1�@�5��#�Z��Xe��TS
Ċ��>m�2�4��D�6��Y�X�z֑�������A:(JD�^7�<�U��Ӫ���Ѐ3�P��(0H7^:'6|�^Ws�~(Eӱ͏��6=�B��M�����H�U��7��ɐ@°O8���T�TG>}jjFHK4��lc)�s�Ė�q+S�c[1i�m?x�� ~޶M3��C �*��I;�bl�i�T:)g��|���W�~�bQ�2%��sR�=/wX:p��|�R9
��KZ��KqR�y�⤲�n+�ݰFjF�N�v�6�?\�GN�
��8�B8��R,��MCJ��^x&�T}�U7����$�E��:����X�qQ:��'��cCL��gojJ�{�lͻ�H���JE Ka	��N%�G���Hn�z�s��a�so(�C�%�0Ԍɋ��+W��ڣ���<} j;W��JWc%!T���2D��=�e�=�WZ�<Z��ҖAfk�y<, e?77��� J�8#S��&�	D!c�fu�΋=z�A���*u0;-c�C��i��9D��V7�LxyW������h�S0�mK&�8�}�&��՗_�.��Ce>�- ��'����ԁ���|a2U���ot�v������u�O,6e��C���_4�2'T�>�"K�/~�����]P��=u��^�����)�dq���b(����jЉ��zL-�^(��P�~S㧒ŋ�"�Ʌ�̡�n�6H ��>H�1�[�75��A�:���b>�ZOX{�7�dN�P�<)�Om�>�O���Q Z�����+��]^�tvy�O*H�Uv��͇U�Ÿ�b�]lǒV�|�Z�"�=!\=(1�_5 b=AXU34�/���a=�%`�dS�Zd�a\_�O%5r|�DRn$m�:�C7�I�(�u�2uQ��!����a$�dT7��¿�6����]>�,��+Ȳ�pJ�jޡ#c��x����9��J������/�C�F6���hm|�N��N�C7Qϕ�8VY��*R��ͦ��������n��/s�\��~�I�Q����L�(Ɓn��:C�2{%�p:�gb�h�� ���0���$RQ�9(�%�賒��t��W�	�DުʢV���Z�X-%M؄v(/aN���ޅ�}�~�O)�sYkg�e�f��S.!:�W�.��c�J���ێ�q�;�I@L��Ұ�8y�w�����<ܣh�q���8h�J�G��X�>�X��R4Q�	1�Q�����YU�^�'��r�RɨQ�OSM�O�8=�4��[6�Q�T/&�C���ZF�Τ���x�h�[�c��Gc?#���8Aw�Rk�Qt�µIjrPD`
0j�EDZ�w[���45�&������)�T�n(
ϢB�̑BP��L�8�GU! ��#���x��D��8�ӓTň�R�o*YIM�.G�j���%��*��=╅��'� w����ǉt!;rt�`����9m������	�l����- ��H-F ���T?�C�����A�B|�O����|�JYl��XO1��ˑk���̜�aՓ���+�c�ѯ��â�1�^wI"Q��Iu�����\�8�K`|iƲ:���\�	�y� f�J.U��'91=��u���bDXp�D�H�$!˧y���sW�Y~�obo�ꙅ4 7ł\L��8��-I���{�s��Թq�6~c`�C�(�"J,J���rH'�$�����E�A4.��Gt�
��N��E쥂�A�2-��o��Q�>�C���q!	��zKN�A:��9!��B>�0W��8��/ǡc����q4 h�h�a�\�1�3��2��p��t+�!bĐ�P�ȹ��|�0/8p�qDH�#)�qa��u��
9窍-�.�����(s����l��(�l
��O�M�.F�|h�n>������#��rwE�dr��r<�:�W
.2��Q!���ܙ�H=����F�uS,`(FG����{�pR��S����W�O���.����b�N�`��"�S��Qju�iN8�!�7�*�ur2�ʣ,ϚU5@�)M�D����Q<.QM9v\�#����ƈ�4�����T����I��eD�-�,��#��rѩ�R�J;�g��q���5�sTp+i��0��A4�X�&%��d��|�R.�+���2}{2����L��Բ LSsQ�_'b��0{����~�\�霋8,�O���n6�Iuы��+68�� ��%3����d�Rı�f\r�k��P��`��2�ݔ��,��6[*��Q�xr~ր��!�8s�@���;��[�2�M�<�jMJB� ��Tm��yb��룘ױ��8�O�m��#I\�T(��[l=e���^w�AjŨ����%Y)�_���yv�aw����K
��=�j�m�q��#,7�M�Y��c?��3�K�}�������Fy�T/>�+�G����7.�b�^�H�>�#��@�,ˣ ���yM��8�S,�	㓂����~D� :��)GҥZ��J"��눙UK��t_HzF�Ǜ��(�jM1�BX֍#"���KĲQ^達y&1�gΞ�Ę�R��tbM�%�=xDw�y��tF4����ˣT|�r�?���8u� d���*r!�.����٣�>�}��,W��u��m`!,�Q{ۆ�M|���?S<�ON-�u&��>:9�M�� (��Ũ`	�Z�H�L�����B@	�tԏ�X������M���;����O����$�5��T /�� 5�0)y7T:u^�뙔��NN�so��;k�J%)m�t��'q<>�<�9��j!�����|����(J1���J�����^�8Ώ�(K��R,���j�zf���r;ܘ��>�Ps�C��ygR��"��S��l(��� �գC�����Ƀ*|
[Q��8�E�,��&>�A�#�M���Mބ����P�lDg�Tj�P������ Y��VH�'�ݏ��(��
�vj1j����x�V�t�9��e�8?w@('%�+�c���uMR%F�A)��{���hO�(�y�N�b����A�@����+�c	Յ�(E5�!o1��)�MX�{PR=,Q؝�}}���Tc��X���n��ϗ�\�(,���(F5m(5_��Wj�C�e)�xRz�ɧA.6 2רe�뺂��z��he�w~�r�6�l�9��z/[�h������z�5U;������81�cB�Hytf�Ձ�&�ԻPt�{b��?b(c��L]	k�X_t�ۃ� ��m��(G$�*��7�H�7�s)G~GE�Xڔ3��\Z Sv�<�0�%��2�3�i+�^2 �Y҉%G�GvO�A�#�p����|��/��!n�k ��x��1�]�M22�]D�*�*x� �NEי�}۱���u���n�H5�
�U<�NH}+��1�g���N�XYiP�h��k�w�5v��S/e�?�9��Ee�x ���{�"��-Q��b�4��I��}�U�z�>דC��))q���" �+Q��򖷁w��E��S���V��%
�$R��.f_dIp|R:�!��&oWp�u�LT����E9襋�e��$O����8C�G��>�3���P*�"}h����#P�bO>'�)�F}�������˄b%h2�u�m:��"(������p��9m�jD�/nF�3{���ҏ	0��?&(\O�=�	�K0^��R� �T2�K�����n�R}?�f��@.�'��Ѧ�Xn�h�ٽo*��[j٣�8���d]�c��`���_�^ih���Zbab���81O:b�F�7�By������Z
Tn��US�&sG��l'����0u+e;���)8��2t�N˞y 1S��{~�ӧ�#��}�A�3�\���W<�[��~�I.��!1z|4�A�0^8^����熼�~^�X�4~xpC�n���wT�4􁡈A�Z�,G#�z̡�_I����'[�~��|��)oj_)��X8R�iD�7�:�뀊� dAQԳr�
�z�K�aWӠ��y
P�U6g�=<ؕ����� ���zc��p�����+�����~�����bt0�3䝏�r�j����^�'��0R�zfz³���!#Syk��$�t��)t��Gٜ�;�sF����d�{�aKMMH�t���MK_�Ϥr#)�}���������k,sd�q
y_�<���ʀ�qEt��u����y-X�j%f2co޸�Gi�쎐\�x���t0���r�/����^=������cýX����a/�m�ұQ'2�n�K2��z�:1/.M^wG�e%8��i
Ay���Ǯ�f)��Vq��^�8ܺuM%<h�<����ڵ+����Ҏƒ�_|n�xV��Ұ�'�UjJuN�4A�F�/6츣�_�8q�^��8�
�L��|�6�4��@��nK\yaI���hP��7ߺ®�Sv�4@e2tl�^���qˌD��yΒ!����b���@�nw0̳z�A�����~�䄇8b��P��|����H��!0�Ϻv��:�@4K:}�BJ�uvyA���T�G��̲�Eͩ�OL�'bx�"�M	+F%Eb�b>)+��T�j_s���A��g��=&����XM�3q����5�T5�xͬ*��GD�P���YP�u�qM(3�����`]QnI�֡,�I���	��V�&d�L2�0�2t& rw�fʺ�בy�r$�����:Z��k>?��ci�i���\]Z.����u�d<|�Q�J0���	9ч�ǡc�[^Y�)������.����+D4�-p�
�㈔����g����tzjү�a)��,Mf>��ry�Gq���2�����o@R�FK���L��R)���T:*���w5b���z��d�P@m��**�V��R�)TB5;uP�bC�@V��+��b�%��nt��"랬%�G<>>����r�ʔ�7�no)�7�U���J1�hJ,1�U%��h�W@�m{���38�G��G�T�C8A���cs|�DD�8�c�hC�'�܎I�0fc�6Ⱥ�3�0GG��v�Q<�=~�D�dL�k2�]�>�=(7��k���O�G�M���2�
`�WX���䧩t)Q�����]�NfW �E�(EG4�u\���>�,*��$��qO�����e<Ƒv��{���y���b4`���%D���s�O��#gfbn 7@���l3<Y�*�W.���^<o��M���a��x$����`L�Z�,ǈ�,)�F�S~}�j�g�=/6��m��fJ��u�2�(J96�g�Dm�0u��oV]̓���Kx�����`�a���x!�ŋ�,��x�]Iʜw�_�\�����i=0J�Y��ٙ04��?a�"p��I��b�N�'ad4L/i�Z[�9:*K*��i�����%�!.�q�
5�<��3jx��w¥k�E}>ý�c�Ut�jq������������������ZPn_|��q�81�1�� 0�
B��?�Q]c�m&��O���P��V{�����V�g��8ɱ4��h ���[�:�B��Q�z�Xv��f�S;�S�j,J"��Qu
B�z�|t,�#A:���t
�j*}��D���1�i�S����|�x�j5/�ݑ2��2{��A>��G)�4oc�ǣ�Y>j��J|�����y�f���G��GtO�Ϲw�^̗��I��c{i����S>�1�(}�7�3W���Y���J�1T�(2����bE�C=1����RU����v��¼Dia�nj�Z)L3�!���O��>c�Ӕ������s)=����구�b<��S�'�Xy�0#9��w4*{B,�$DP1y�CH���h �ӏ)%������A?F��Ĭe�؎���ɔP��;wD9L^#�����#�e�@�T�|�����PX3:�>z"ЈC��9���]�tJ���=�6����=oa�h�hDF#l�z�*H`����aX__��u���Q[C�@}Cp����@lMS�X]���@�,c!A1�
��Gf����0�NS����8��	��p�i�tcA22k.���T�d�"�i�ǋNGL��2���$�X>��ЉD��z�؂�%\��J>3�o)�#mp�b�������P-H�C������F.eR�3j*�/����6UO��iN��-[F�+�h�M'�fnO��::�@e�lMIɳ�5q�`��J)/�!�=��g⥁��ZҌ
�k����[���!�U�2\X()��Bqd��7
�5�ik'&z�ށJB�����
�t��aL){����?�@�N_ll f�߸~SG��5Q�e����ǰ��əH�Q\a!5�#kҌ
,/��:��~VV�˟p1}(�bgo_3��~�=��85c@���� <x�T�|7���K""�*׎h��
��gT�!�@�SHHe9��#$Q1]K��W�cӾ
�Ǟ�&!�{2˜=p/޸��=ӂ���P\�Z�2��zw!�i��4߰-6�b��G�-�!������Wr��2��6f(Y�1�^o�TU��K>1th��?��WΞ�u4C�������_�"�x�Nxnb	�
%δ��3��{�,N_����.1�nd��B���˕�t��(�3�������~^�>\��U���e?Sо�f�#�� R�z�}�F2?(<���h�s�Ȓ���V���?�1Ί�_:�	��?ƏY�kb²y�ۦP�D�S��A�VT#�J��g���1�Y͠��<��ta��+U��(T�g��D�ߺuC�QN�"s����[��vk�,����!���F�uO�������O�{p�yfי�͡�V�B!�� ��&;wK#��3K��`���[���n���NlF`�DΨTN7�;����n��� ��������ٛ1��u�o���mStey1|{Kb��#��Uök�"BcTR(�b���NoDTBT�c%<|�Xe�-������z���8&����\�[�-�y$�G���WT��|:��s�g�6E��D-ka;�e5���*:L��+4S�[XB�OA��ƚ�����08l>eb$�{p7L�1��f�f�f,��rPatxhT7�5b�����t�ظ�0j˶�A��m�Ėe�Ǆf�4�Ҍ�|SZ��zر�/�s��7|���~8��@=�
l��]��\4~�M2�?���j���V����p���8��%SJ���0pD�yajH�3s!�ZN���|�P�<�ytU�6�; �l)�+���F�V6�V%`Ak�1�d��)��̟�nԢɌ�[,s ^�ˌW�]3a��h�d2�>�_9X��\J��@f[1�T�aO:��טG�A"R��4g���	ᘿv�eGJ6�T���� �ad�tŒZ�}t9��.����G�h~�VoN�E��+�m::pnu/pþ����ͺ"�۷�I���\i��p��7�w�l� �1����>������ճg�2i��˦T����9�g�y�s�^��~!{E�1;;�B((]`�J��5�P)���l��@�*�u!�:�} K�D	���,9> ���܉ ��~�|C$2N����	�٘-v��I-_Gx�"Y.����Z}!Ac�0	�LJFn��8���vH�Pt	���w�?
ׯ��	ڍ�ÿ�7�'��������C݌Đ��x��I[�ez-,Ǝ��ZW��i�nZ���}/�(������p����{�{_��ǟ|bI�n*��Q�zY�
nF�]W#+�oQS�����a*��zͼ/-��Z��+�l���G0���O�ugD+Hh�����)���|�Hj"�!'^EgT#lf#9Ul>���$`�r[\Q����8�I3acNҚJY�~67jB} "�?ܯ�m��$J̔?s�X9��r�rq��P����)r*�����F�!e�8�v��$!��#3��ͪ�1�q}�'�WWkZ`և[�$�AX�j�ـ�q����T*��J[�:W�RfK��(��\7���ZV����[.�9�!枹�&	9���1����N�G���#c!��}Nj	l&�t���ƒmJUfjr����Q<c��ٳy��J�5[����ܹ�)D��VI:E=�E��w>j~�l~H�v�/]��N��<7?���z����6�W Q��X7�Ұ'?�M� rT|#�-E�GǬu�D+��|�4U�@�'�;�ߔ$���Ʀ�X���<���S�-�L���?�(�L h	 ��Q�=�U�Ʀ����|�+��vL����H�d�"1�� :J������ƂrHn@b��q�I� E��a���E)����A7SȂ���LQ?��O��������?�/é��L�A� ���C��6�:���nr�Ty[PV)�T'+�G1�]�"aG^g#��1I���qQ	Uu��&dq)/S:�9����1�<��?�i  cǗ#�X:�5]KP@�%�Fk�~�fS�R]vѰ�Bj~g3���k ]��>��4���lJ�L�Ӭ�d�k4t0�D�, %����.}�Y+
X�nd e��z�g��v�A�,,��YY&�6$4t !�)�*ab|�����'
|���֟���Ǵ[�-p�L}ZXS��/M��)��rY�G�\�g66�0�[�?��a�0o����<t���X5�MKw��	m��ڢ���\'l�V @�ot�bP6Ӕ��e����-�q22�(��8hQO�L�>�e�f� �i�d�ڼiz"E��G6;������j���/�	33S2)����ɿAO808jA����-�G���'��t��Q���%�5cIi!W�ν���V���e�8����p���H��u5�����8��̖�l���T_m1����<v섈WF�,��5����mˀ��;<�/�,1)���Q��ɰ�~0Ts����!�+����H�9����p!�{���ʚJ���zػk�I��v���&}�n>��Ǔ����޼u':0&ǎ����dfh~zN��ܙ���r��|�[�ߖ�$C���Q�E��<�9�w���U�B���S��+W4ǈ	z��Y[̂��>ۈ;����̌�-H��6����k������(�|V+��en5{��h��=~	f�����!
Zc��Ld�#������77µ�W�)C�̲����];T�X��θ��Q���d�\.��¡C�u�@Ob��7\a���}����_=<��N��R�w�ȑH3&�6�vlt$r��zzT�Z�o��*�|���~m\Z��Z��fL�cv8�����<0dڼ_f�(H@R2�522�葟�ϫT��ߩ8��D�>�v/̈��e��� �q5���9�L�Pm?���6�.J��[��{�����,E�������:eu���H�{P��g3��0m���V�z�L�	'����
,<z�R���t;���姦�%SQ����V���\&fZ	L��*|.�u:�Tc��o���+�.$3=������e��0�:3;'à�L�=�HR�k7	�e���F@E1�P%`�ص�j���4��)^�T*&.�8<�T�P�&����:=0�2>�l����u�����%~��φ�Nm��;2Җ��jAע��l�}^T��XtS��^�������-��m�	�x%����ɓ�Tp$� :$��7	��/_()��ہ�����n�a+
F�p�+F*�\~\�+�G�y��z�PC�����ٳK�.�Y����l$u;�N���5މ%F6$��e�E�'�ȇ�g��P��;!�̶Ɏv<���=lW��DYQ�.�V��k����6���'�����RZ��0*�9PZ3+$ev�\�&HΝ;�ȇ���������֡��>�͇���,��R����q1C�)f;|�w����I3��2�E	�x&9>�M�g���g�ӟQ,fz�LQݶ��:d�DyD�B�ح����&c|�!�
	������5P�T�k6�z�]�t>"ͽpV�-���S�&s�%����V���8���=z��!��-����ߗ	,\�!�����>ᯡ7�c�D�C��oߦ<Hbő茛�g���W��{�.�R�,�����0e?#	O�SF�(�:3��z3$*8�Хp��Q�Z���Q	�V�Wl]�,�\�H��x���r0�[Z->;�MH�&_�vټ��M��Wi�E5��7u}�lw�w�4<��ia3�='Y���^�ܾ�(���^Y����*̦L��-��FH�H<��zS�{�� %(yN5�e>k���� �!JBb׮:eW�]~��K�#����Bo�L��BSJ�O-�����|�>Qq��9��[J1i4�8��0�\Q_�k��B�a����̏��*M����(kA.����ĕшk��҆l���T��~� ��{w���H\�E��nO{yI m���踅��ʲ����r�z	���A��aS�d�bP���[��`D`�%�l�#��a��=��8�J� �D!���W�Tm�!ϔp*�����N�M����I�oܸ�>�6w�,ü-dZ5��JV�3�o8�13i��Æ�r��5�*�К�&y���(�3����=3�S��6��z�X����5K�-[�n���]�`����ȕ��n�"c�G�T(���Ǉ�}�JB*�~�&"#�b�fN��D��|��O`���#����E�з��J�ݻ?��^9����ou@H���#��q�琉����b!��ɵ�6�@(�����^j��'��?��S��0�T�	<\TyE3��Eh\90=�z@���Wכ{b˳��ڑ��;I�������z��^��T����I3�EC����RDSo4z	t�@����LrҢ���Q�ՉS��U;$�R�5�.����1�1���k�����J�h��29 ��4 %ZY��px�ZP���&�f�6%�y�0��"��߉�h��w���hkˑ<�5x�O�L��0D�����{�<�8VMohj���R:�E�"M6�n�{�(>[��KP�#U�E=���)G|�.F��9�':EP/�� 	�Z��ʪ�#	�M�?nkG4����b8`\ZU�VXYZK�������?�|iTP!ăA@�@D/|;�i�d&D>��><']�B�&��y�T��?T�#憬��T�m��c����سxؚ��1i@E�eb?˧�й�����U���%���]G$q�=S�H� R�,zr�/f���e��9t�px��u�AV����[�Zh4���..U�ЅW�n��/���=L	t"�eD��Y'~�|V�F����{[@K��kk�2,D���|T���8�l?����V3*DL�����W�
�.^�w��)�3�V�W�'H��~&�sjŧ{��v0^:}ZU_�'aO��YV[a��\jyn�E��q<������Vc�SRR���Ȕ�#��� �N�f�<��3�Aʆ"���qRʀ���9�tj8���~���f6�T`S�V���V�Dp5�Y�3�w����3�U�����yĶg�.��K0Ծ��tUڂU���tj1d�о^��'�
�0��{̊s�CXw�౦�N�?$��	e'<�q�)6�E�C�����!ª���**�֪>�OR��H�Q�H�U��f�q`ǵ��#�[;˷zܳR��On��2f���q�7)1V6i��af���a��frNٟ�j���ܶ]�6��fT�⦺������a(�]��C�\���J$�_>����c^�H���\��䓲&��)���~��G7dHξ�l�6�7��(��GL�@���84r����?�קB/(��o 7'�̒�n�I���:cE"�����(p����)�M!�#�����S7f؍EA�jq����:@7ڷTz�-�CFb�2�.]�T�{�o��w�牪���q��Bɵ0 y�v(�)�:��W�������+g\�A>��b�䷿��ݖ1-��@]����~���T�?�^�GX���9���x�r��&�O��㺃 :V���W��R�ҩ�~�KeV���e)��Z�7-��%�;�����Ő걎r���m9�Ro����5i��o��>	���߈�	�<��t�ٽ�p�x�B�Ǐ���'
Y=	�]g�'o�:�B�tZ:�_]�(�Wa�#�ȑXJx{A��S�#�M��،Z�)�D@�z�L-�29�.J��C��CH՘�R��_�Á�xK��I��n3� �N�0,�"�rc���H0��aC|Ī��fQ�YY��:�~A��Y��/��o8�X�SG%g�FJ?{������>��i	R�����;u�D�o���8�z��p��qs���1�WR��d���m�|�+{������߆3g��e[��}������}��pĜ4K �q�FrK�b���:�������m3q7����z$x�kz^ ܇�������>��/D�#ڝ%��A�/�Zd��w&�����" ��F��e��o۹�%&��tl�Q8�)�:=(��9��]��̆�;�'9��s���
co�:�Ν3�O��w����<�s�m�Z�%j��aͮ��Y�fr�����ۊ��T*99R�B��54��`@���4N^�概|��w�M����2<4��]�D�WOr��1�N�����	}� �'U\�DP8s��m�DA�Z|X�9�0�!1�6j��JN��y�!K��We�>��I�=)?g#��H|�3Fdcs#Һ�ʂ��S�0D�5�y���f�[fw�<�{���_�);p8�<{N�Y�DI:KB��"��gΆsg_�+�ϦB�ʹ��w���Q������HGP�O���5s�͟=��k�v�^1�[�h�����9E�>֝UB�p�3���:���yU��|bfG�"���I�B���F��$̷������DH>�?��ޘ��:[��^ٙ�D�H� 8c�k�%gE��U�L��.ڝ���|�����Ri \�r#�U���ᚙX4�)(��Z�|��8E�;*��}]���e�WT'K�������������X'4Ge�Ν;zY�2�E�7N�yYP�'O�*BLyuuC84:�X 6�⡦�]Y��0Qp�������[�K�К�#0b�24�,�czwՂ�+w$����	������2r^�"r"-N;�F2p�H�fO
�T�Μ&`m_ɂ){��rea�B��Po}"�W����l�ێ�t�^Y��,
�{g��f=�F����D�>�Mc��֒0�XKY�@�c�> �Ϥ0A�gl�/j��z��K_��d�))m���̟h��A/���Qϐ  ���v�u/���u�Zcw����zb�G5i���v2D:U�Wr�f�����f�9�P}��o�u�ٜ酧�sF°݊9:N�6|f���"��`eI~
�/�C[��KG+˥+f�������#������ӧO�$R�k�������Ӄ9z���R �3}�}φ�A�=H��F�5Rx�(���q�4�*�F�%�kd���=��s�#7}Nj�>�������2'j&�\���i �o�^��gs�Yp����`��@k��E�z�(�,BN�BsQ#	t+��h��P}�md�!��ȃQ��+�(Z���|�N�>���'?�������G@���f~�� @������Y^]r	��
,$��cy�*�Df7�nQ�y7�DZ�h�0I�v� ���&�r��8;��J��@m�I��t��*�t"�-�k
����� ���搳�8����`;̎��:#\ϩol��@F ;��AJn�3ā���a�Q���$
����!4	P%�BG�y���dN)�pp���9levN%����^P����z�9;\�6�Iԭ��6�g#}�W#�0m����d{��,8��gy�|���H��<g�OB*�
��nyK A.3碧Ol�50��� {MQ��EnZ�.H*���cԢ$�r`ݐ�,�,R�L2i>;t"���5Cc� p���SK�#,��$�bڶ}TO�I��Y��̡�r��]�-n�tpJd����9$�ΘW�3�p$�e3[��5��T���Q�$�D�v�Ӭ��
��ea��q&׼�MSbY����([�1�l �!�����a�ўH�q]����]/�W�TT����cn0WRHF?��39,������ʼ>�/3�|a^�a$�lԉ�&��vE��R]H��6���Y;�)Ao��l4&`I��5�0����%	>?�%�J(���'�D���:t
�?h�����e-�@�s�}�L������ㅛ��z#lJ]�M��w ?����뫵�ȁ'%�$��&��Nۉ#1O^2��`�E�&4<6��G?n��,�:�}�bJ�3�A�l�.^�`�΢���6^�ȑ
��}{��|L=}���9Wș����XT�	��h[�'yCu������?�zyP������q�p����[�БC�~�~��0k*�on����QA� �Y��x��N��T����3�B:6�ÞD^}b���f`��Aj��8�d;��D�G���zVމr��N?6T������&W�.R�����r�=Y����|t�T
!�۬������^{U�Q6�&�d�,�������%>SQ�ߠ0'Q�L1���):�'|������_�\?v4<�P���_�QE�֭�Q/�-a��j�_���0�{HrA�p��%�Z�y׫�$���&����`(ȋ�^K#��z�#4����|]7���r���g�n������ 	Ǣ~�VA�E���CJ%y-,�&NHP�F�ـ=� q���Ts�}^\N�Ç�\�)	���������$���{W��xͲ��;-Y���O���|C3��r0��C�_�B$�)�8)Ⱏ>���]U�)�xyd%�`N��?1Ŭ��g���jQ���@���V���Y?���׺P�qrO�eJtW^���9�D4E7�Įي�Q��>��f���	�l�:���b��7���];5���1]��Ǐ�g�b~����p��d�'F���A��'ɶYPn�ܵ5L�zX�lz�n�.��SQ�R�b8�ƶ�ο�Ţľ��޳g_�/�r���gN�E��h��'"Y�0y�+$&}Byn]B��;�"%!X�n|�Y�m�ZL�&s��
u�?�[>#�/���!=�����PJIW�+Ƶ�q��qhǹE�,^w��la���nȫ��&�	q�����~;)L1s�K�ᓶ��	4$��G b<�!�����.d��@/�����m����/.�O>�Ğ�����'�Փ'�#q�ŋ�d�&�~���o���;
O������
��:d���1��F��M�)a�9��0وNR�6'��B.�����T���,1.��D�r�;�J�e7'wMD]�EMAu ����K�VTE�6D��?~�s1�:x |���2	8�=�h�J�D@����5պM�.>��~��脝�gv[��P`&I�-��}����I��Ɉܮ�;�N���@*�'}a��t���f�&ë�N�Aѓwb�cef����rرP��NۃnrB�/���~3f�lDXly��ہ��Г�.bˇ���h�5��:��-����퍜���$�v�صW�D{4��՟.�!f�DowS����M�I6���|qU��g���)��{�7����B�8;0&���K+c����7n
x�}�v�X�]�F��ᣇ�F�D���ů_����RtP�������xX�Ϲt���M3�9�2�7j� B+y{O��@��pk!��AH��t$N�|$m�H -lN]�S[O~��0���*Ӄ�n�`�by��Ji�S�9նO�������.Ӱ^_�d\AT�!Mf�½������UA���EH���ۏu�0{ ��X߾;ܾ�4<zz=����m���V�[{��Ec��N����̈́�v'�7C@��޺uCu�m���-"kFނ�y�-�g<z�<�	W�t3ܴ@Rɍ�A�i/[�Q�O3Z�T&�\cieEEW�6`%"*�Td��Vun�ر-)SC$�3��}֒�O+�����ZOm�E�6'��v4�?&"�ݮ�l��`�Ʒ�rn��U�����7{@	B[�N9� ���D7�چBjj\���r�EB7<��ei��l&��� �{�n(o�;各5ԋύw�1\C��-8�t��q�g���m8���[H$��:����#Nz+Va��Di��"�A�aN�� �
�X�X���^�À)%��*P-�o���W���D�N����Y���IHIt��y��Z����e���^��nW�U�E�Iؘ[wnhc���҃]��?�LC�26R�����H8�-�o�6#�o��������e�h�j�}D�<k	g��@�|���p����gD=S�$zT;U����aˡh@u��n����2�tչ5]�������ʪ֢l���z`��錞�e;�U*�_�7$���Q�%�U���O:� RF�&z�_��6N���S����;$fѩ�1�J<N-��2�!B�������h�-yjy��n�[���ݒ�xl�S�[j-�38����67��>[��(�����ʴ�� �G�{�5Ad]	t ���tG���(¥�����"�̍���l3�������E�t�B�w;����oޕȔ�-x��)$y���>\"�g��$sT`;�v���ł2mg1X�Os:Y�z��B����3@��rc�䤢7jW�Q/~�ĉ02^	�͟z>~��2퉨���1�T�Ep�|l6�Az�ϜSDR��5'Wr�0�I(%�UQ�+<{��Q�J#>?��7{} �M��U�/y�9�N��#�����y�$�N\�����E��7���T�A�_l�N�ܱ}��O��Vv�O��pR<$sF�M�5�]���D�����򻗢��3S/]��k^}2���-X��בk0�IY��_M�`͈�,N�����)��_�5փEP�\��lޞ�.=��jY��P�댳�7 �憳���u(�3N���g��k�:�L�5Q��|�7��-�����Jd���8�83����7i��Q��m	��-,�ں� %u	�>�����J�΄��y?�28�HI��l���������{SϞZT��=>s��L7q3`;%��e"��Um�`!�D�Ad�-��%Ε��8_6I�k�OR��As81a�(?�XP��萸L��Ll5������X	����3Y*,F ^Ƒ�N'�ðpDL,�
���GN����s��_��_�_|>��c-t���o�!��'�.|uS>����D�:yJ'�������>��ɓ�Qi�q�S����O��%	�s瞙���5%J��THĸ�]V��p{���uM����3J�hdtT������j�F� ��K��J�ԤM�\t�
>�~F5�x�Yk��L�{Ԇ\�ć^:`��5$����8���x�:+^YehdT7�b�)=~��#�$-�@_)���Yu	��'h���Q!Ů�>a��4���}J�u���)����*��cz�� 8B��N��������Z�3D��r���P�@�i3c�l
�y��.��Lͳq�œb�!}D�?f��A�x�N�O�(�B�fc�%)bÎ��3g�ʌ��=]n��kJ��^�C�Q���ڬ��8N=�n��Y�c��FQ�b��Ͻ����Tg�gc]��d Ԏl�C'�����'�:����*W@�����C�4A&>�k� j�����+S��,��E�DTZ�ߌ�-�Y#0TZ1'�ɚ�CDȩ~����]_0�F��D� "K>��`�6Z�Ul��Ƌ�2���$@C��� 慲�6%�#���T��X���E�D�;���4},l�sx�,����'N����2�8u�%%o7�|�?�ף$�Yן��|	961�����9aq�ج/��2L��N�)k�X�&�`�|Ms}S���t��lg\*��Dm�I`�-����Bĝ�D��+?�U�k%V�ki��ڕ+������� �HG ���f��TȽ09���ı�c#�]���5,�a0�� �M]�p@�_|&���N�n�-�}�:l'��8�dȝ�s�cx���z�w�9�8fֆ1�,x]n'����ᙙ�;���������
�ю�O��q�u�5C�@��~S�_�'�C�f��qțG�\|u*��[���S^� 8��r����㊝1uȻ���z��6��"�!݄&<���ܚ(��/m\����|1��s�	�g���m�'�S�?aЅ� @�[�n�M�m���/���G}
X"���7�юlv{�����kq���h�I]�7����\c����9L�^Lű���,*�"�a��	?���,y�Nr���Bu�ç�Cr�����oVj@��4�u}}Z�SD�*1�ZQWtG�,[LL��@B���3[���k�6��u�-Zlv3���uK��NI����3p��˯�?�h�|S�@�e˝����g����4��y��M	/M@q�~�P@A	@O=�j�@�lKcJ��}B��K��Mi��\���x��|)�;ک���ީKYdd�#�fÇ�A��� e�T*%?��St��m�L��z��wyO��2W�зnH'��%��p�`�٘s���-���?r$%Ȑ_KG��	y�R�i�qh�V�ʥ�Fm��f&`�چ��ɘ�e��+��ڍ���I�S7箓e7�-(�:�%w����C�?#��Ug�8�C(����m� ��k>��YS��	E����s�$ө��`=|(,;&?�F�ɨƆyO��T�=|6�������-�޺Ɋ6�'i��|���)���Vϝk��`aZ�3�H>�� ���/
Z}ue#\�v]�3zd��?��	3���`�CN�0���e��΁ba�>�E��a�drǤP���2W���P��y��rK��`sS܆5�h����&}��?7e��CՉ�Tf��vi�"$s1bcXra����^��M�9bji[p[����@A�����zѱ����S���5��hF�e��2;�V�3��"��k�Y!�U�o��Z`�m�F,�X�L�d����� �ܳk�mD�,)����������p��U]�};��/g�d=`v���_���G}�l�՗_Ӝ�̓�a6m7�L!�ڴ%�]W�#�h�)�#��Io�HK�xx����x�M���
W�7z	ԁ�t=�fۍ��;��%x�BथK��J ���,-
�:L�x|$X3����9��D�PNk1F-�=���C(�q��s@,�s֘%�_|��}�4�N{��e%�(�1X�ƭP��cZ
[{���:�3��ݻs�e��\ ��#�X�Җ��42<(��i�Y� *�� <��K�y��f�0'�ĹBׯ���UR���O�=뮶�ͪD�2�Q%y�7�L�.ܒU�-8��u"��(��/�xYQ֘c�1�xQ���z��g"r��M=X+U?#�̘*)���^���s�|��m!8xD�S�f��-�4����e�@� ,'l�\�A��ԥ8�O�>���8yB�����R�K���U2�U����)��`3Q���҃G���4��NE�� ���y.�LO����f$��:�Q,*:>mS_��6T)ljV����5���Խ��R���EyGև�A�^v�jG{�F^��C�u^�u�M.�y����^u��99z%�N���e�ˉˡ�r�Rl:���ǎ)˽y��~br�|�}����|4 5N" ��$c�3�r�G����ơ���1��O�(�, �g4"t'2Įiaª�]r�8��-�5~դ���F�D���r�>9t3Z[I�Q� ��;�߫ȊM�Hͅd�iu��Aj]u�J�9@vh���2L?#�x9��&v(��fZzpƚA���j#�֦�*��y��/�l��l�7���*��^��D�	GN�|�QrJ%�@
��*�1�����ko�Y���Ĕ�����@УÃ�Y[[��R��"�w�9�A�s>��/����=f=[���~g���t������,IPt�f[�&bt]u����sջ�c��E��=�ܪ�k�=����b/�r���m �Y~����dZ�R��@�:�@+�.C��)A�������yCv�E��,�+>LѲZ���i���>�ĉ�A�(��(�1�� � lH����U<+'9	�D!I�^}��t�F.6����VW��tr� ��	�ǟ� �'GI�$�"��{4NN�P���7��J�E>�/MiY�e�z��E�'�o�ů�b��wĝ�
jP�C��rG�A�o� 7��Ih�W�i���9-r�2�pZlHB�F@��S+(|Pa0 ����-�K�,�`&�((�p�Yʮ�f6]Z��F��S��@ՀM�Ɔ��X��W���0��W�FScE�#r9&����%`KT<1l�z�[֝�iE̗3������a��?�[�F����O�3�	�è[-U��v�ĈN��l���}z� u��M��S*��P�n|���G��"�80���c���:��`9��|7�Ee�1��bNkқ�+LuLD���Uu�k&�A���g��sr�kHP���r`N$�Ѣ �;C+�SKQ��y
���9X)-�Da�uI��E���CCZ�Uшe�d���q`�8�U*9�����^�̙�D0À�!{I� Շe����a�+�U�(W'XY6_���4=��?~���%�R"�SF�-���'��S/�
?��_h�;@��t�}T�y���Qa`��γh}�9A~�!I���`Y��M-4�8�DzC��Į��k��J
L�E.N7<��%���\[r��	�B���8�d9�\ nVr[�h�SQ�I��E 0�Y�	�Cʯ����U۰��z���{Nk76,n,����ŢK�;r��Ȳx�e]�+�DCw�ݕI�{ϭ8z䨐�!��qiN1�Ʉr�l�����F���Q]��܎!KE�KG��P����F��?_��i/6�Ky�P�o�S	<2v�&$�I�L$��q�iYKz5�x���%M��J���\viml,INT�3s֯��3�1h>�F}��Í;42���n�_:�S��������20	�3SX,�e��� +D�t��Ԍ�!h�@���R��l���"f&Q��	��\R#����3��;�S�p��������8JR� ���fcS�EdAbK��LzTc����� @_����fI�̡�u��CR[�_�����g�7׏䆯�eIy9]������:���l�@�D��pJ4mk7fuyM���r:eNQ��W2�o���]�.#��	���;o��g03>T֯�����аc��rG�. ��OY�8����"6/a� �IF�y������Zn'��z�m�UG�"�Q~�ji���ZCo0���7c��u�|ʁ�#��:Uio�
\ݏ�gFΖ�Hß����+*�0��/xyiJ	���P9���'����a%YQUS���9����ݾ{[������-����&mPj�#�@�X�����Y���8z0�濎�!�Mbt�'�b�l�3��l&��_rrP��[�����8�dR�9߽6X���P���ǲT,���Z��M�U/0ʅ�Q�8��,�9\���i%i$�����">)�؟kݒ�fYhs�l��k��v���kW����ɫ�we�tn�T�j7��?�^�\�r%LM?��BmGC7�#���pFs���?����ܣ�����Y��w�M��9ɑ^vscQ'���Oߞی	8Wml*��ϒ����6��t��.FznV�A�	��Jt��nD�H7��RY�
m��� H�QQ��W�iY@h���o�OY��'�U�P|8���Vo������-|��j�O(�7��F����t�-&:�MNUv�@�;5wZ�N2$�<�\���S)Ü0�N����s* Ҝkv:"�-.�rqA&X5���o�����Ci_#�v=�-7�uÄ�~��/�,�N�)>]��z���&*#�jY��N2���I&�ySX���=���6}����6�:���H�R�-�����o�D@v�>�#{չ�	&���`f
��J�_��OH�Dk�]k����ZS�t�Y��왩]a����mA�f����ٸx$��mW�T��+	�.	k�n�{c���bW��������5!M�Uws�PNѥpoMף�&D���^#m�C[2A�`'� �XRdT���Ke3لj�'�.�� 
;_��-[���Ed�rHem���Pb��a	e�\Լ��p���A9}e�9���jL�g�7P�ry�L�h.b+��RI&bh�����ID�ڨo�_�u��JR�lS��dj��������s]�s�D�O���DQ�ވ"�C�M|�*u'�I�� vK&a��:22	��s1b{CR��=r�`�Z��u�U�WVEY������<�M���l�e���t>��F�[ͨ7�����RR�v�lx����R��	�'�ia�0Oj/��f�e�Pʻ.�CAS�2es6#ysG}���X�S����<�W)+�\]_Sv�4��tjO�s����p{��oc��0������."7+9�������U�|��˗ͬ?R��2��Q���iVh�P~�׷/�b�V���*��O8�A]��9G7���v1ϱ��պ������dםT��i�\��o7����R�Ļ�Ҝ8�UYܻw(���V;�qM'?Ģ;zT�4��`��17�K_)_���b����F��䔍?q�4��֭{2%���5��N߻O>%��w���UR�\���NpP�:�(ʹ��@O������.Bw��Ƌ��<KL@��TL�z1m]U� �h��H/w�����'����������^�jg&�	����#�p*j�7��y͎�A�կ���Dm&�ga�~��߅_��*����?������҄�����{�|����֏?�$|j��O~�S�U�V��;�� 5Bz�$��G�2�i�ic�>%ib%`�#хNǵV���r�=ԉz��t�:-��ShK�V���4&%,� �M[���Q9�Z��~1]@M��w����([�I�["9���W���	��9��8�]w@���r���^_^��y������V�Q,#1΀L�TH�$$�I�~ �r�6e|@����w�:t ��2���E�Y���p٩���x{6�����ѷ���=J?'��$���,��r^�T��l���ɾ!�`1=wsm)��iY��v�Y<N��m�J�8U��	=Y�n�����<I���u������ח��f
Q.��6����h&��CI�$m�s^C����l�/�P�P]���~��H�r��~�-U}V�7r�ڈ_�FN��FZp�e����]�'��w1����s�X����ӽ)��x$H�'��R�^�(���l?�Y�}���@I��/��@�(�|As�]�Q�A�IT�K�������`b���hS���$�,:9�+�����=0��>O�7�8�
a�0%v���������[�o)	��^����� a /��,#���@ȌCT,����lQ����݆u��e��OHW������0�}���0-��=`C'j�'
;�o9u�cJ�=޲U�_P<~��E��w��#�@C�$�hB��y����N+N�ü�W���ܒ@q�%��nN�M�ܴnS%a^�\����^~��-��p��Eoq����@�zXn���J���j�8D��Lݹ};�r�L�|.��/u�����N��k9��eՈ���KϤ�?�ֱ��ș"���ٔ�(f�TU ^fZ�Oӽ�'��j;!Ջ�<ܗ�g�{�媲��(���|#����ʈ!`�v옔i���(YAݾ�bv2uBL��d�����s��~EY}Rm[���)��|_��8LK ��ӧU�Y��VK5�FNI�駟)�z�7�1% !8`�U�K'O��X_o�j�J�vBiJ5�n�q9��8�&	�I~�!T(hx��?���{���h2��Dg���Ӌ��s`{�^b�Ad%�v��4�S��>i�/�p��/6�eƃ����l%�����s:QR]�f{�2'Lg�G?�����&$C�����ً~�{��^x38��=#���__���o��I�p�ԋ>�M��w?PO\%�bI���\^�ЦB�3�}�����>rG�bJ�V�I�ZXjU��V{|Z2�(�F`k+s6�wO�XΠ�qfk����Ǹ:LF�H�:5پB���2���ⱓ5��7e� 3����iF�|LV��S9%^A�_~)�M���揟	����K/��'�oiE�Y��3/�������~�.7�ŅRXx��75c�,b+
؋P�����C�O� ��V��mb���Q5�k��f�� ��q�-������j��� �VO�;�8�\�P�	g3��"S�7�d�F-@}�}PJ�?	��<@�&U�''���ݩ�W8���9�;!{!�%������"۴'��HHb���F��XgK���M�"��?R�șB��@>���C���^W��7��W2vx��肋�9uI�N��R�C1f�W�����U?�]���TQ�(mQI%�VH�z��ܽ�7F�+E��TlۦTB��|���N*��:#��!��8+AuR)� u�fHD�|�ں#KT^��vSQ�z?������a�k+
�Q�~���] &������I�K14j?��T{�9Z�8�S�z����g��TvQ�8���C��ƜECpZ؍MU�}a��c���:@x����j#�Hx��5�t\K�[S�lfJ>ty��Dl�p��:�C�����Q�ᠸM��D��H�%>�lZx"�&�qf�,./��bQX�D���aKQW�M�"�h0a�9�8r��G?��K�ơ~~r�(b���G<,/�9u��C{�|���eY�E�]���w��^�^�ߑ�G��3��*�s���H�ڻ庢MBf�@d�r��0OH�½�Ŀi�@T%�|^��ߙ���Jw܇$�V�A�IIxe��Ռi�C���rkF�FE|M����S��"���T�)K�l%^.��eL87���DD �ON��{v�lb*xH���P�%��0��D9⾵g_1_Gy���^Ӏ)��-V��x�;�9*dd�K����	�i<��k�l���M^��'ԫ=	$x8�Ç�`��D��&���e����P�C8��PFI̥�F;[\'��44�P �
l'׉+z��q�J&|�W�
.��U���p�&@0# ��T���]�0uAc�Е9���q2�y�w�r��q�n���ί�?���Iņ�Mߛ���\�)�4~κ
ȭ�]��\{0��IJE>��u֊�23w��U\H��(	�u�f�lv���=������]z�Y���.��H�����m��"fJ���xs�+��E�J8�I���>�Д��M6F'�2��^@LiC�M���2���PS۶��%Z#���ӏ�W%�lI,���S������zVA��eߢ�6s�-�e`�c�W���P-�:�F6��Q��g�ܵ3LK�oA����~/g�hdx<J}�s$$�_E��;�I=zr��x�}�cfyG�g�@�ݎD5��ԅ���r�T\3x�E���#}�&n��Lےec^<�g��0EÖ�'vO=K��"
��f��?َ�
W��yo��D�@�+�3E��a&jn6L�����B��t����͛a����e�<���lؿwG����~�{Im�>bNxL�٘P*����q��U+�έ+*͜�8�Y&�2�޵�f��������J:�%��9����Xߌ$�^����E�t&�%�Ő���c�ָ����>�.��G��4���])�a��\�7��)-� u�J@���YR���A�\0�kLÚ�%4'�U~�]��0-�M{dr��1U߁t���G����������N���q��s;�y�-����i��%�C�v������ �����1�o���rL7��,��AΔ���aL�軫aA5�-r�C��e�
�m4]e'�<p	�k��O>$�^�g�N5�?a�������,��k��'"�D-{�C���v^$,�����	XkY�X1#
}���*���H�4���S�*b�OK諸�?.{����8�(��g^o�)z����]er�N�8e���Ls��{0Q}�C��Z}QJ�U{gpÜtz>RE�v{ �|T�fʗ?c�9����+^��	�o�~]��%�)16���bÖZ��@��:#�	�1�a��� ��Iv�5�@y�Ŕ��%����[p 1asߠ�[�����J�q�U������F	4 n�ޔd)?���.�ѵ�~��0I�v=��?����y�o'���6��
�Tp�7L��;�{�*��C��т&� LG^�m+H�x�gL��\37����b�k�ԉćy��)�]'Ά�~V�6�����m��nB��3 ��P/ǱJ�R�y3-8pgڌ�@��N[�����$B�T	V���f�`m
DVA��b'���ڭq��N좹0rUy�#GN�5�s�ݵӿW_�g�妏�qFS�#��*[g���*�W�f���7l7 �nL�=#��c��l�����b���x��,���|�,���Oj9���զ]�o���Аw4~�}q�d�����Ǖtj�%ѐ��!WD�
{���
:"�O�!]�4��i��3�hAf�9q�`�a }>���|u:i1�b��H�)nd�5��Rš�0ag�`��,��ȏ�hutG2�h��'3.���}.���}^;j��k�9�cAQ����>V�aU�Y[tiUU%��a"ء�3�XJAUI1�-�ګ*w;"=�|4�v�f��N=��$Yu�ےy*�ʒU'�I!_,�ה�B�z]?�%��1�q�uM�GI��ʶp�a�@�0�q����}-������E�p�]o�,�VPBa�XL4��j2�э8'�&�k038qrߖs�0�ֽ�A���vn$u�~��,��J�`��E�q"�,0��wM�p�?$�$��k^*J�[��z�%*E�7�+�5�z8G8\,9_5�y���I,��n�W���Ph�pɖJ��O+b򩨼&v��ح�� E�_؂#A�Q�ϱ���ۅ~I�kYԖ��6����F����s� 3	X��V���Ƶ���Ʊc�*(�r�}Q�=U�ڣ�eͤMckzJ����5���󨹞|﷼y��U�Ai�q�FP�"s56/�ї�Jݳ!~&��[X��qt^W]<gj�~�����!�ނ��I$�Į�3;�W��^ɚ�'T<%Md���9	ɩ��OL�wT9ئ�`���6Re�����t#�伉�&�m����:]r�2"��#�qUDnc�Iar��;�Xl�G�
Ж�A��c=HH��xN~ :��lꅾ���rxj�	������i��pG~��Y����l��X���a`F4��re�D��d�� � s(�(]t%7���M'�p���_=��P*���Q��A�쨏K���]S���Y���B7'��ԅ7��x�M�}�v�T3$���z�	�ygmq����I*щ�a����HK����lܸ�GG@�.H�z���kɊ�<%SRb�4�#���t\�QH�\1,Uk�Y���N[���ZW!�qe拾Iy0�����0��zQS��$?|�3��z8� ��\6P�zh[�>�J��Bbf�T�qf�$�{q�mjw�|�چ��,�c�-�u&���4�ޮf�],��H|��$|kB�D��Ej�z�h�~��f���
��v�W.	яo�#DP1v����VÌyE�>���ؐ��>��D!��3��f8Ô��-U�&�_� ('��5�:\�.��X� �5n7�
���F�9���8p�*��\6D"��G��y}���eͱ3R���2��Q��X7�7�������m|W��3���O���إ����E}2+������mA��a�:N�p����Ӊ�y}��!��Q+%�,{Ϟ�"=��/k�`}mY;�T�e�;��Jߠ� �>&����k}��7�����IQ�j3�c�rg��� ��@��dm.�U�Π�C$��F�-.�(-��u.WTU�pؘ7�3a�cAx_����!�O?���r��v��`G�݌�j7���gX��K���L���̖CT�KPFUޮ��-.��,(��f���\V�fc}E�DQ��SU=�m!Acqv��f��=Q]��C��.?����AC��p��Q�;MM=Q����K�$WA��
1*6�R����y���&	��;��>mV���5����&`b��`��i1Vͯ��5�����k!�2N\�`8�p�;�CV�	>�^Kf�6Dq�G� ;�}�~��{$BU"H����\*��  @L��5)�#G�)z���)���â%u׮|���w��n�i{j���L�K���	@b��-������ͅ�=���8|W���LՄ���>�(�U>��Z뉩���7��@�KP��8?փ��W����y������u��'	����ߢn���u�@��^��ֆh~!�C1d�f+YtL�݈��{w͎�*�����^
��a(%L���G���}��_U��"�LN7��K'�*}f����kN04J$����Kd\�Si��3�=�a9�:}�j�d�!���>x(�%��v�w�K+�!qJ1}v�=ñS���QW�F�e�>׎�X��J���	-��e7��;����E�%Y������Sw��Llo:�V�C��J��5.�)j�0?|_�@E�L��H'KGprl�����+4m$N�
����zU����>o�RиY
�h�v�Nq��!_[���y�Q��M��YELc�*>��Q��f

:p���2�� 6�@$m~o}Ӊl:���MY����� i��o�m���9fn�ڦ��������75��)L"+j[�5R����:}l5N\��ƾ�Q�n6����[�M�X۰��:�& u�O/E,���4�9��@�0�FՕ���O���/���ߔ��VTt�G��e�(��1]U	�Ͼ"�=��b|bW�l}�r� �
}f�Ɯ6)�3~����V�s���N }��Y�5"a��^-�W��p����e�Z��l�t#��S]ZD!,�/h�}G�����_�W�#�Z9D����	�G��8uV,�]�n�ە狉0p°$P��c;�'����.�ױ|���=�v}�k�Veo�dDX�vΓ��$���{���ҥ�4{��%�%�c��Աѷ��
׮^�ii�/���X���cH^SK9��_��ZUdH.E~ѵ��42,�<�������@K��H(�P���C,_�P-�a(��Ą6�*��6O�(��#P�H�V�#"WR�J
��etI���o�q�0W����5ۉ#�Ţ���y�~�b҂#aa� �PrdN���i^
n�|Q�8�����3ܹsWa-��ӥ��D��F��[(��8��ͺ"����M�i��!�L����JvM���UZ��0��>�\QD�>s^����n���xO���gR��ϋXC	"��:�ŶY�d�H��B����T�,�&�x��|!�td"�vU�vM���BمX�2,�=n��6U���^�[�_T��B� ��b����kX3W��y�E)�:E��Y��X �ʊ��9I��SU�+
BR5�Rc❧���Ui��PZ�E��<G�oE(�@B�I��@�
���9����~ex�>:�Q`@�:��vSxF�/�LhL�"�m$cw��Fe���^7J�#a:�d��t����ĭp���ܸf�,�h8�	�@hǦ	��|�H.
��T��-��nz���x1��H	&�cu-����	ϳ&���8L#����N��SO��d������=r�Bg�PH�N�0���WW���:�kɬA���e��g'��\�DA���1�k/4��s9��I��ŭeϿ�n:�I�'O*&=��зRЍ��vT��i�����H�NH����݊�<��ڑ��I�c�XK�+�[Jђ�Ƕ���x9G��A�3xy�j�n��)���?8v���˱@y�ĉ�01���m�: $�� #0�(R�>}��%'6��:^e޽kG��=ba9yLqW��`��#�v���a�f�M����X6��;U"�|��+��B�B��\����3
����R�^��%mÌ�N����w����|���'�w"�g�_�ue�~��^�������-ju�V��خ�(n�_^����Ț���ɉp��I�(k�������^9|����o���G�a���=���?�X�num%�o�'GDg�~뼝�R��/��r�{**�=󲸹|�5<nܸ.^��h�rN7C�Dw��q�ɪ��-�K��������z�~���4�WA�����	�ץ��t�ժ_N�ƀb��E�}��uy����M$>z����#�ѳk/&Q��yHj@��;͎N�өGfg;�MG��r=�7<2n޺!24����>���~�;oi���
���$�#)�0���	Kbɑ<�/�`Bln2���\W�_��v �ȥ|��k:DT `����@t��@��=�V�y�@S����PӴ֢�^�g�A��EK%	��umH"
��Ԯ!Nkt� �%�gfZ�<_��r�┱!| ��wd����@́V�}��������d-(�=����}���~�M����R~������aZt�nؕ�������s����߻�|�M�������ۚ���Er�?�(�@�D�ލaP�������pY����]���\AA]IG#V��4�fӧ��4�5�̳R���e�G��vR�^�.Ay���q�Û�e+��f��A��>%?�(���)��Μ^�N;u,2~G��^����cGUf (X�fYs�#���}�yط�	��|Y�l��Uk~>C2�dƥK��V�o�y��-5���D�:u-���1C��a8���v�IQ���H�P����&Q	���	h�Tf_�{=~�Ă��g��f�Du��r+<���Q��'�lIб#�^ީ�;��Z�}ϔ`��z�RȲ�?`:�@�_׃q��q������j]�?3��ˢ+nU�K�.
E��3B_��@����l�gs��#	%��V��R3�Dg�UVA߄S/yX*����!~�{�W���_�*�M�ץ�������+{�<�b%6�9a����TM*�p��FF���A��a���-���cGZt�����Bᆶ��;͎3��\���E�ĩ'4���eqv��쑠q�=f_�]
����>*?�g�$M���O�,s����̂�5@�L�D8���oh<m���U��1j���`7��@�� ��B%����d�ͣ9�ɓH�:WV�ڃ�h@4�d\�Ň~(�`�=$��Bi]7K�e����գ�#+7?��3�Ȱ��~١�I	��+Hd�\!,!��*@`,!b����p�5�K��zGH@�!���b�B1\w����d���hqi�B����ڈ���A����7�Uc�!OX�n�}yI��g���A�p�oݺ����B�5!�L��~n&�	^*�2��L
s�m�T}�l]`��0O"f �r���;��b$�N���2I�KB��,n�c���Jt-����\G3bg1?t�ঢ���`?��Ca��]�����?�vP�'���[?���T��~���1�d��OW�/~���#h��+8�����P�O{D�����
Oũh�A��{@{���r��>�B�Åz���9N{tdL_���%w���y��s��O��t��m9�5��%��/�H�F~�RO���]Z��G�P�Dtm�գx��/�d�+���&�)�.;4\�Qݙ�sϦ5=D�y�bx�J3�O��ap��GO�����M�Mq����O�D8���̎؅m��s�Th:�5-_ea$�O6�Z]
��!M�I�6��ۉ"��)��c,	��U�Ǭ��>��|�S���4��<"/�m�k�B^�K$��e�f|#�;���k&Ae��)�4#E,7�AD�)��D�m���]+�3s�,Sm��� �����g�Qs���'>G� BM9]��-� l�#� ��֮�Cɵ�W!DG�%)!�~�X���v&�(�Sl;���,	Q��5�k���A�p�fS��Zw���QQu����#6�|F�60$mD#�b��@ 8Q�V�Q�ٚ�+p�1W����AY*L#K%�ܧ��r~�G݈�Y��#ݸC�:.Y�s�Nԏ�nPK�Hԇ��R���x����]�ѣ{��ݹs\}|�J
�`��*��8a%~dfv.<�'8x����p�tI-؊J-M1Ul��!ۆJa�n�&���}���325�ܾ}K4���gG��Q�l�h>�N���p8����H�Ӱ�G앳�q�l�O/��']�X8[I�P=�֗�B��mVQ�2�u Q��0�*��o�
�]y�1�Qm�⌸�Ԥ��xS���Y�#�hayi^W]��;«�^���N?����N/���֞����n	'��1�|�;����4?���f��5	�6��Ս�(g�C�ڟ>y��A��?��L$]K���͈!���i<y�޹�o~�����'��i.�q�L�_�n�*-Uz	퉈�>h��t�V���(�CwޒLƩr�<��LDa� �"��� gzfJ>��M�W����q��e����?p0?�9�D�]"ŶL�!$cӰt�>�h�>�����pТ)"�n��3�T?�geD��n۶�p��~����|�j7Ys��eS
IY�?Y6��{ vڸQO����е#����d��mgϝs���p#��)��I�{瞝�k��K�u8��h��á��p�q���eQ�Ty�uex@#:?�CQ*��a5����p�Wg	���O�)�EU�=R�A�jI��KN��Үs*gf��t�}�m�x;�F�A�'�|cr�v��$<�LG�A[����ǎH+?���������(VR�������mρ����͆v�@�����0��f��~
?FYg���Ӛ s��Q��f�&�(�l�]�&�����)DE�0��	�t�|����C2�����CR����8a5��;NO?��Y���$��<����������&�T-�GƠ������*���L&�2/xPW�Av+n�{B��|E{��V��q"�u�P��5-T���z(R:՛Np��h>�M���}>�t��y�|lܼ��%Q����͛�����;&�������ɨ�t��U�0`��3���*���G?P���ǟ
�J$�ĕ�Q���mc����^G!��bU:AM&���t��v�S��LQ�E���/4����G�`)�)��Ȇr
>x<����X\>߶�zY���Ν�Lb��0d-�ܝ;w��8(�^=�%�����ǁ��yX[��K ��U�~����pއV09�$��n�7�9��>>7���k�n����ۑ��ԩS�F�շ��������z�r�){�=2�T�Y�%��ej��h�0rV���L�q �	>�wfR9P�u#�'%~]�1�-,����,y��'N(<DP�����e&-�%88`6z����%L���in�yx���e���g¹s��-X�I��Ѿ�s�Ϻ~�9�q3���80h�}媅ާ�o� +��NVN�
_4鰙���~G&�\�}�%���ޅh��={��0N�o����ݻ�����h��r����M�8� ��U#�rA>��$i�V�V��2�Lt�lF!o�����S��O�&���+)Ab��g/ �j'�t��n*!I"x���~��_����f����1:y�X@���՛ͷϣH����fԪ��k�n�kd�ν��Y�$7��� _|�m�AM�޿W�I�Dd����ѱ�鍚�Ub�5�l�e�1�u�D$��]A�C*嬦SSs��T��C��#)����o�L��ݓj�5[=Z��%��&��%�[�=�Wg��DF&�Q2�!�t鶦|G����qs��
��m��֛*�(�ܾu3ܲh��#)�0)u{i^� �&�&tE�:L\���N:|��Ө�\R���!�Pb�5l�IaN�� �lzf6|bQ���)�gQ��0\����&(�r:<x��մȵZ����y��GT*a���}�4�����_r]ٕ��	�$@�,��R�L/�4���^3�]�dk���V���r,��b����3û9�}�}	����23��{��{�>�,�!~��������{��]sE�E���df�Ʋ<�n���Jg����C�'�����4ڼ���|FzW� ��� R~k{W����
��0�c��掤�i	,�3!,������e�2:tK�YA=������4g��T
�<����81]�?R���i�3��!� �f�\�v��5]\�z��:��%Q�!p�/��_�|�؊ך�R�Y�tk�� 	��t'��J58dr'A��K��=����,���Dw�E�e'&�U�҈긑����YU�v�j� d�-J��B�)�0�LJ�P�9*\sC�avv;�����KN�"�����I�?�F�=���z;��R�'�	.
$Ԝ�����{]u�j�S����0DgX�Y��:]����ú2˻���|�k*�c�9I"�)W$�����ի��4������- 98�׿e�%܃���=I<zA4����>,W؄<�])�bJ��a��-<�b�Ç��5T�9:N�1�N'� �����-�X�����Y�Y�=�@�+��sR4�3�nwnC'h&#�)�ć�Ӎ�[��}��@�։V|öi���CO�>�v��Sjdww���S3�d��n�[#����"SQ�gICÖ�Z\Wi:h�|Z�H�_8RC���jz[�\ ý�8T��T<m�d
�LK�d��"�7�uv�-�&�u������8ڑxf��ƿAr�J���u��cIg9z�4�T*,�dyɁ55���, �����+�{��%Ye��[��~֝F(�y9*�M�KPWl�����	7��v�"B����/�������L@3-�P��sQ^(���Z���ͩ��ɳ-u��$G�]��Q^LpS�D�㇗D2g�t|c�����2�șs(fіz��A'�GH`q[Z�����	��+�gԂ��7�N��WFJ�Ý�	�����'��Fu�t́ ��1!� 3�J�SF��pp?M����- ��<?��k�u¹	��(A]eOk�#9��X�Q��MP�Ѥ�{1R ����c2P;�X�A�wFN�c��s:�nʓ�{ӾF�L��*U:���������1Kd��͛±���[[���7k��
�k'[�!��Ym�+�+�;�,U��?��2-�ڤ�|^
ϓ��jMҏxgfJ�����iNCj
�@��ϗu�ZШ�@���'E��*M�u���L5>����i.Py���43�;R]>Q�Ѵ m����.N���;>s�d+�ֿwv��0�dhH��!��D���ډ��$+��4�����N�6��{�1�̬�Q�H���ɉpsZ�ۍ�k�ye��E�d�	�W�>�:���U��vt�!:0��8e�M@��sa�iRWi��ө������P��]x��Y-�� (.���X�(UC!�jgcSI<��4���8�E��g�ϴ�<<w�0���aWղ��9i��xp��l1 �<�=����E/Q?�����G%=ά!9,m����LR�u�Q;q�C�S�`������B����eWmxE%��Om�u���E�z^���B>|�@�F��A,�Q�N/ڱ;�����:���K�.k-p��ZE��˶)�� �b�},uU�1f�hr'c1� ���gH���g>R��E��}���AƭVUQ��[�qL��s3ke'���N�d�c��3D�M�i�`nZToΚ����Z�=;9Ͳy4�>}Zt�;5=�%�*ʩ���>3wA�׎(��z�RKl:�U\b�Lp��$4��[����X�T\_��G� ���?p�$��h׵�h���T.g�XG��G�88��}y#�4�sbw�i��%�Ƀ��^���ÚT���N�R����ݒ1a�¤�T	4�a¼�f��C:f�"���iF�Q2&2���;|���֨�z��{�a�����]un�i� ���.�*C�<�RPwxK�T����-:Rme%P��j �	�	�Z�̣E}GE=�=o"�zАj��[4�d�'O�V}^�����CAZ<��d��H��^F���]�ˡZ
��zx5n���y9���q??r0�J��ŷN�n�T���鍜%yqxo�w"\�xᬮ�e*�9,l ���	=�|�;wa4�an4�P2_���ɗ�E/Ϳ2o���eUKlAP��Q�J�n�B�XCt$��ak|���]��� ����'������bS�y�a�cq <���0Hy�8�?~��2���mJ�A��g4���t>]�~M fH(�޿{Ӥ`�>|��@ې�s�8VM߁�GzJW���2i��6����鿿25����W�\�u<�o�S'�K-��Z\�S-c0����8��(�˻�ڛ{x�&^�=r�ד��+;Tɸ�R�$������q�Ą%y}$_���:Ԑ�`"��$Fq3�$4�&�y����B���	9B��u�9x��4��VP(��IpP��)�h���i"�@l��G���~�$����:�O�~�E!�?�㧺��?�Y�|劣�5���Z7�w�r�Z�B��?���C�<�8=�Ϝ.�g�-��q.`�U��(�q���ݰ���3�tFy���+!0�-o��A�����u�A B�4�R�MJ�G���QC1L�������f����R�#�i*J��{�<��)u������zn���7�H������X�a@h�I�o2�m�j�{�����
��T����A�ӤTN����^���%-��'r��>�T�2���@���Ғs���a�x�G>o�B�q�I}h��� �M��8�Q�o6�9�6�3�qU��Dۈ��F��k�򸊊��H�:�?w�t��-ϵL�j�ʜ&D���:C�� [�+��^7�x%�Z�g�%�+J*?y*�^ߔz!���:����1��E$���_�2��+�D�'Meb���!o����Q_H_~��l	��"}�F�S�ɜWW�*K�{��Fy%��b`%?KA��.�*�y*�tO���n����pҚ��6���rL�� ��U��<EN³ @��~�j뵸����𖧑"(�4ۨϧ�>�P:�l�Y;��$�����gSǌ���M㫇����� վn���ɟB�}�&�ל͂���xn~Ʉ஦�ANP�͘p�B��fWQ�}8��y����~�^we�U�u��!\sa4r�X2ߢ���X�9�|.բs��|l+ϺzvU�C�Ɂ��>�N�����c�EA�G��`x� �[�<Bb8�=w������v����7B�`7�Wr�.\8/�9P��`��\}�)g�����;i{���Ѥd��\:t��E��hͧ�������^��4�� �o~����{�p��t��C%0�׫��m�����m��4�WR�#��O�<
��K��=-8����6�x�&PR�t��w��c��C'�'UC�� ��s��7���RI
 ˥�?𸊖65@��hʅ�UY�ޘ��I0���G��ePAp�����>-Bx�����Ͽn	��ͷNbO]���	��+��!0�Mf��=x�*�F:p�pzi�ɖ����Pc#V1�"=�l��Ի��e�nܸfц
E�/��Z%Yrc9S]	9�:�sT 2�T��P��ʽ}��Q�6�7���P*�b�M�ۂA������P��P�f���`��E!>�ۛ�>�*�E�����7�5�g΀V�k0{J� �SP{Ϟ��hϴ�������{AB�d��4�����=M[p�X�)� ��w�9SO��p��Ӂc���%4�9м�~�y�@̃�+_�Y#�>�s#Wu��kR�J�����Zuqy�*�>�IZ=�,���NTS�F�^G����y� gw����b���#i#�y1t/��m�*�-,B�H�+�,���{�ʝ��B[<
uQ)Y��5�2:�>?g���IArqY�p|
Xإw�~G�d��߉��R>x���.�%d��AC�j����@�X?u2W�`��F���Z���^7`�I���5����Q�����`�+@n��vp(>w��ʕ��0���a�xgNM~N$12����u�Fإ���;J���)W�	?���'K��������(��
�F�(������R�E��(l`�',v �B{3�?�7iZ�͓�i�.�&��`��NJ���b���0�CY
�ջ�&o���5�g�8RxD��7�|��B27�K�Z��A���1;lY � ��W�f���v-hQy�� H��-b�ZKS���I	�N� 1)�Gs��K th��v��Z�53���H9��������G�ff@{���U���YEJ)�v�3��jj&��&�MPȀa"��|�K���{��^�d��Rqm���y�{�ܥ���Ȼ��P-����J/;�S�k	�\v�.*�/�F���^����l)§\�~t�沩 ٜ&��L�F��r s^��y�UE˵�EF��8%��#��tp���}^�p-m�?ƚ�,��3������@/�FPpHK�I&�ϐJ��H)E,6C�p�� @�Ũ*�l���=��A]C��ӷ�&pN��Qvjԧ����$�����M߈�t� �����Z8	��g?��a����a}𣫚,���c��@�#8?�����a��@�Esj.���YQe�c��^g�4�q�PoL9�F��81��?�x	OAgm�r&Q��<)�w�f��*�3�>z�kߒg���E
Q,6��;��G�Y�ݶ�L2���7��	�9��;�\T���Gu������1��_��|~�ڽ���.ؾR8͙�����Ϊwc2��K�k��;�������'I���3>S��;r�ŷ�%G �!�AA �OMz��3A�/�-(�_b�������(k��y���N1�(佉=�mҚ�fZ�AB�B]9�	�Wu���d�8�Jk�][��3�"�2I��i��u�4�|+mm�� �-������<�v�,�8<�Ξ?������ǏS�>g}{[��/"�1�淿��G�s�b��n�K�|B��I>�՘K���Ry�,��vlmt�`��_z�C�Jy�:U��r�����N�(����U�0�JG��ύ������OjyR�*��52@͙.�g�^˛z��W�k� ��1���%Z��Ղ�`H`{@��b���%ҿ�h�TV��R�6��J4���UQ��!������i"�o��Ƽ�gf�ү��o ]O��������:�hK���μ{* !D�À��e�I&R�n������n|^�N�O ���c%:�������/ҷ����?��2�7�<ely��-xF�W���?�v�!�f8 mpH���cAXkb2u��Oݜ ��͠%g0���T$,_�Fx���x$G���16�c��~S�D�^wX?s�H>�Ac_�-��P0�T�gL�L�VK�Dm�5����ҕ+�r������b�94�פ��T��^?����	 T#�:z�D�[p��g����t���>n�������β�&�K�P�����f2Q�\��#'�����������,1dj�sY�<�D���uA�V����X�}}P�d�������*��.���
�+R��5uO��ǰ�w&һxP���I�܁����>;���MSߧ���_J�����=Rv����\��'ω5�v9J��yEp��*�ؼ b`;����z��ͨ�@1x��eע�/t
4��l�|�����m!��	���ٿ���Q'����ש�f.�A�!��-,��;fO��sWϹ����ډ���Q�9e_H,�c5�LE����!��n���؈]|r��NE�O�A��s]e���(�H.�sjC���H,��G���0�ZH�
�Qѥ����W�
=��@n����m0�χ�����єk�t,,�f���C�1!:{)�Ŏ���L%x���-�.ᇙ^@j���`?
N�q�G�ş��Xe�J��#n�����e#�պ����2ȸ2�|�!���%����I�A�?gB |	A����
(iq�{Z<n��7Ŕkl�F��IE1�$3�yl�墿���Q��3�x�R5
Z4UsH[q�S�f��B~���I�U��.n��^,���H�*�c��A׮gB��M�ꌄ��$�8,��Z��x:Vnj0���Ъ:�ȞR�lssc^c��4A�G�7����$͈eG�!v�+W�����w����C�uĂ��R�"#Վpp Z\}��߼y���I�W)ЉD�<���>�j��y��^��w:�>�L ��Qڣ���;�4�|ڎ�k��z%������n^���e�M�7�7�B�)�����n�;>	Ȁ�e������7w�߰*��L*��ֆv��2��.[�#Gh.䜰YTL��t�'�>?� FVE��u�q ���(1��4�x�m�2�b_kR�Dd	�ɚ�¦���L� ���/� ��J���PΫv�-�A��J��^�ҧ�\.��y�ˏvZ�� Xc|6����L�0u������?��f`o�5m6��	[\z[�Q�	`g��T�F�v�܊���H}�6�����4{Й�Z35Mək�����R�(�B�&�NQ'Z�*�����X�F�q���- �&�G����>rH�]{s���)��1ԣ9>ǤݸqK��������������0����eknK�5���zѬ#�^�+��t���?�m�h9(�}KAY��U�Pܙ3'-8�-m`Q񻪝������Q�z��)g�t�\�� �y��9�L`�Á�u�3Ft�T�;w�t/�q\�O?�4���h�u�'�t4��W��4�X��s��Qe���no�mkNȥKu�X`��/]zG�I�>}d��"@�m�_N������~��i����;{F���<�;�p��^��?T��kL�͌ax��J[b���+�����z�X�u0t��Oc[Ї
���k+����=3����C*RW�_~�5Ҁ<r��R�P�rTq{i�سr`)����Q�Ǌ3�r� c��w�E|���qɧw#���	9}�zQ��P��6U0I]P�!9��_}`��A�H�B����5{������ 3���!2�������l�M�'.=z\ �O?��l�ց<��8z�l �I����v3�o�G�8:�ߩ��`��bK�g�o�n�������	lc��抖J#���đ~ДΝ=����C��9��H
b&U���x��� ��h[���x���;�˩��N�m�߿�n�v��s�&�Fx�Y]�q
I��1���'���8�~�+��]���9	d*[Ї��fP�C����?N'N�Jx��n	܁���	,W�}I�kb;Nۊm��n;�6|p�x4. �E�a)��qI��\��'A�1Ѝ�a�X�n�HO�<�I;����N�dd���I�c�f�>�/�".�qzbj�bxYT��c��}�����?�ې��E��~�P�fFNMވ��H,W\_�{Ho|g�x�Q��	_�|����b�I�CZY��J���c'<;~���[`��#�8��<:�M:�D*	F���X�(ஔ�q?(P�ݩ��)6��9��a�4�Lʝ�_�i�v_�H�"�ƌ�?����W�1ޱS����//��@K��4�D�[����խ;߇+</)%�%�c^mÄCS��T��\Ť����wӣ���w�iz���J]�����/�'M���)�0�3�e���Z�)�8�z�!��u��4}�6ֶ�����Z�����E�k�+%���qI1]��m	���M���p:��ʈ�j%��1gC9��I�K�LN�>�,���O�v�'�ǈn;굻�Ŭ@��Q�/�������sH�:~��'���E�� �)	���uy/gO��j#�Y͹�5Z�!O�ۻ��:|{R.dY����Mu��,+��W���>��3�isc�N�s9�^����#J�3�� t�ѮC}��@5�r��sQ�4����A/�dr�zE&?�O��&����T������GS���S�z�ۢ�`-�JD��i�k*洮����� ��3[p!����Ddf1�Җ~�6jdj౽���dF��$�};�R_t�פ������3r���n�{��Z3���5�+"��,�ᘼ\Sj���띳���Y�n�O=~�T�\�v��$X͛�Y��B�Gb���|�4�J����GՐEv+���>wؔ�X���\���)E��ݤ��@m\�I��X�[R7-�cIP��޽�F�A8����5�W��1�{ocہh�&}v�jOX��,�JqH������ǿ����ߧ{�t��{J�|��ע��VQ�8h�/@�����:j�ц�$9:��`�ٌs�U�+�&.-v��嫊qn޸)8�'�jJ�����ϨY�)�X7l�w�}��}"�B���'���R/�ߚ|x�"������f57|EY�=5]z�:�lSp�]�%[�.]���]�6큔7wr�)@h�k�d2o���W2�$������4S21/�������,7��~à`�� �X^�K��.�ZX������<�/S�<����v�}�F���mKMΈ8�.�>FZ��PF�1��d�G;s�IhU��6�����Du6�4~�QMm�o-,18�����\�=��N���*�2ZYiҸ�a�i��{#�F�$�����y�>�P�%x�3�Q�����jw�N0��a-�H՜��5�E8\ֱ�B�o꫻�T�K*s��Y���Y�������1նϙ�h�u:~b��¡t�Ԫ�>�������J�Ƶb��5�[��a����j���qM�c�h��6�۔m%=g[��~�J��gϺi�U�)[��'RN��x����lH��@�>��{
SJD�JG��O����H=����4DQS���e(>o�$�읶(@t��S��d~��(1T&-�!�1�	/�葚c �w��yE��fVS\"��Κ6��\Р���J�ʼ�]ض�����ɳ�=� Mel�������pц�hkTT!{�(��{�*�Ǐ=���,j�͟�u�uv�H�T?�80�j{�#uǿA�$��)s�!E D�6��	? ����M�ĀEb`�Y]P�4P�? ����W"@�X_e,��ٞ���=�_�*�C^nTR�����WX2��i��4����9yc��t7�����7�w�6���U�:P���T_�ISS��N��a�`��rDi���m!G|ښ�.�[ڣ����H��
4�B�����&5�ܦ:}1m5�E�?����ZP�<���B���$!K!�͍ϙi�&����6�����������r5�˭���O׵!&��գ����%E��^���L8"����k����Z�զ��p�h�����YP5yp���MgO���tcc[�;���8l���lP[}�=��#aٔ�U�M�T?q�~۽Gث�ǩ�D6B�8{ޖ&D$�!��w�&�J&x��F��ؑ�}Q�W�~������s��j��K��ao���i�3y#�K鑟Q�@���Y\F3Ȼ�H߅�_�᪌=���+t���%z�RI���)��^u�z��6��ѭM��S�HX��I��T�K;����w��[�ӘS���,;bA�nE��c����S�Xj�;P'�w��b��~p��  zIDAT���YZ���$6�L�#��5;@�}E@;����i؟����Grm�@N��[�aR��=�l�Dڨh](����3+��G�0<�z�Gt��!��7�_	��hx����;ҟ�-o��V�Vb����Rr�k�~��rZ��ZԐ���P�Am~8�ʦ�^4b�~���������#	OC�ۺ'@�4�(p��w84A�w��B��n���.�J�a伺1a���醴/^�N�j������������kgX������5����n�8��)�K9����{��M���ǋ�)��T�9��PW�#G	 ;��4ov:v��V������H}i�l�g�r�uw��z�l���'ц�4a@m� �i?��lC���\`N�������_��A"2[dی1���@�,^׫W�>Bv�5��6����-�_?�MY�^͌�e��(ݾ}Cx�a� �j�P2���v?��یy���,�L��������<Y��)j����SD�w,��w�Պ�YaԳAW|�ŒJt�Vb�B��V����K�
���>������w۞X���P�T,�5�uWEy�H3�;�H;�LOhzz�
\Ռ�{&�/�Zէ���}�;�ҩ��+p��O�T0G` �Ra��qyx�\����j>T�t��
�vwwSu:�Hy�2ϋ	��s'Sg�v��;������~8�Ǐ�ɀ�������hJ����'������V�L/�h��C������ZFq�Ng3h��m?�yT�*otb��d����]�w}t^�6�no#����N�3��f�Gl�$?~�6vQ��ܒS�ɾC����gO���)� H���!��J]���ޯ����t�ѭ�3��{��/v5L[�����{�呶4/˄�?J�ע�S˝m2	M��c��L=&����Rr>M�}�u�X$�������gD[����*�U0Eӣy��t5鳬��}g��NoWE�cսb��Euq��D��(T��z�aߋٲ$�f�gt��+���#]�Ce���V�H
�gd`ɤ���+��6S���$�3A|�)UK8��[��>,��p��$�Мۺ<,�h���9��y�N,���*�Z#8_��D(z��U�{�H�'�hK�jA��o�6g�NǊ蕐(�%A��|�r���<���SwFR/�VM��, ���f�ˠۨ9��O�)�`?(���1����^�d�	s^��U��`�����N�t�WD�v?�Q5l1���m�oj���b��ʪa_�:o_���(�1!��?(�\�<R�U�Pɤ�jF�+��]2f'%-�^tQ�7�/9��:��7f$���E$��}��|p�[���aPIN���'��N����g�$j6mdGEj��\WxZ�H�^z��"lo���́8�;E�ԛ-G:�� p��(S�1��$G�,��C��Ҥ���9a5&��嫴t`�;�*S��[���P`�Hɐtur4�~���NV-`�]
��Y�}���lorjO^�1D�'���in�~g*���rzl���[����<҇X^��I���`(�o1\�{ΏB� �%���nG	M��"v��~NК�k�.ܖ�U�QD�^95�`[�@�r__����aT���܏%#���B��D���E�R�t��ܗ�'��Ȇ�)\!8L��e�����v�\�!�>�'Ͼ�ܿ�e�8�&�6d�w��z��źs!��EM���Q*�3�ӀB��n1�(���^
S���t� �{��Ն�)�*�[.;G�;�hދ�P�ks� *`SX�A��asZ8�n�T�7�l ���#y}�v_P��_{���]?)E��5M���-xug�����^�$��M@Y����N�EN�<�R9xq������?R�gb��q����>��M��Inc�!H�/�x�����&*�==���'����|-C�L���gO�)��G��>NZ�#L������]�ا�$��G��tK&����-���f�;� ���;��U����q?7.�Ո��Iwx����HX�q0��f�'�`�����5#�U��99�t���rn߾��?tp!�%�0J���,z�����F��j��!��#NXt�Xx82��ʞ�?����?�/�����7���)����i,\ۼ ��c���E.�ni)���>"�Lqu�k1UC��N!J�@�����|h��i �b6��`1N9��MԌ�Pc�:����_�rrl���*C ��ş<{�,��dy�`���-���Q���BT'�X�"�jq���1̌?��d�1XL¤d{�RJ���O���?��)9F�ŗ�����1�S�����ܑ�C�3 ��SȢ�a���~��݇ϴ��(��(������U����(<�˵�4�l�ӠIG~��w��1��YP|k��꨻Z����5?���Ӵ_�m�q��O_lo�&A�pvx.��ǎ�P/.��$������$[�8Y�4a��)c��}LEY�GT]�v��BJ�p$�G�țM�@@v|�=�Q$����ZzB�#�0j�G��<�a��8Y����$Ѹ����ple�8�Ɇ1�H�;6!�E� N������9�33:�pj�����ť5m.��
0^v�E�	1gJ��u����k�j��;@���V�	�Q��k��{���*�xl��HN"�&�w�7��N"�@�]H'\A�7���#����cg	�t�q�����o,�6�_�(���"i<4�&.#9��ԛLl�D4=�;�3��՟���y�J�t^D�/�"K��wr*R�(�1�ӷ��]��/��)���>�Gɣ�3���Q�����p�ɽ��xnh����zC�d�R�H�|��r=Ng=1>T��~eČ�8�o��&��>o*�B�ݼ�#G�,��% !���TNԗ���,<#��I� �����8=��,�5�j!�hQ�zo< ga�i��1��%�6�R��詶�i��&og]��D��R��w�b79t�a:=����q��
B��	C�/�Z��^TNv�;�]e*��� ��z���}6`�%�<7��/X-xy�$�) ���)hL�mll��55Uo�K��Ҿ$�歛��5�Sk ������84� JjbϢ�,��/�ԧ���w�o�J3��g�����G='����y�&Բ�!4 ���TQ����T���щ�}�����PRi�A�oq��\��j>e���;uՋE��l�� H���qH("��N�����참:���S�%�/i'��}^H||N�4�M�dcX<%}�y[[�Mnʨ*�=��Q�#x5m�B�����~������4\���CS�;�PJ�ՈQ�n���Pk*	/�&���*Pu��n�Ȇ��6!�xo��<):��fx�$Hh�T`�+��� X�nϯRS��unj
 D�i7��%��ǇW�s#R3vrT��u^�9��/�m���]��TI���&��F�D�U  D�:�J8dgRM�t����Y�԰���������\«z�4+26�2cN����SI=IS1��bM��#�
i_P�����d� ��_qC��E`��X��}��z�<��9=�ܕ��|j�\eN�� W�i��4zA<�c���"͈��+$EzZd�M"�0�G93iY5�<v)����R�Læ�}�8����ӥJ_W�J��5gN�>�/�i�7x&y�d�q��`�]O���m*G�I���b�As��+�H팂���GH�qJ�v�!������(<��:g�-(���K!ޗ�q2��\+Ԝ�4�a��ڜae�� Hw�j��B�m@�>�>��J��b�����n������'����Fm:O&���r=%�B�TcXL��]���)��T��U�Q��%��r��2����u/��q�{6�ެ;@B���W9�^TVJsz�8"'�}�����I�C��OUI;̂�wN���T�	OHT�Zw�DmAL:cow���S�U��0_!����E�vP�����c=TFkdr~U�έ�G�c�F�P���j:E��!�k@!�{�LQ���]���gZ�������	'�B�[���%ي��d+^I�'o����gX.ܼ�F�I1�!��WE��q�Nռ��8<���h�E��MƱ�X�J,$�N�T�Z��c�S&B�h�n���@�Y.=E���v.u��|9V���YkL#��v)�,1�@u`�#'Qȵ�ܓɺMs#2��4���}@1�V`���}�8�V�z��Δ�%eDv��1ڭ��# K�ގ������xQ�0�I��a�V�u��>#��7_#���2i�U�|^�R0�j���WU�����25Hn;.}��v����T�(�MC;�&�������}����{@�1�>�Z�f�I��ѯ��*�W���f�\94ŨTu��˳��d0,�7�h�~C4�;���d;�>��R����><�f�vdv���sHl�0�o)�B^�NVY�Z�(�k�_�)oC�����>q��`sK������X��"Cರ�k��Q��\*�W�,��8�U7���%#ٮR�h빂6�*T�MSR������� ��fU'�a��?2ԍ�~�u� F��Z�Fͥ���ۣ/�����A�Z,1N�=�ז0��N����ٰ;����p�s5��t�A�l-�=�dk@�н�i�A*L�2�n�~Pq��K����lS�k��Q�W*m~��4K~�R�?r�B��&�kǨ�}p�OM}�[G��w0�(��WFu�i�ƾ��Ѥ'��Zi���=��E�}��4�'M'1:�I�( ᆧSt�)��m�h:u)<3�e<��騘q�W]p�f�b\��R~Cz5�1�<�� r�c�U3�qD�KʟQ�^�Gu<��ǤP�?�e��,E
��ԉ�t<(n�AjJM��T�P����)�S/���*��g���S_�i)6M���c䈎�c_*X����)�7���)6^��zK��**OݙF$:>�?s��G1�+����B(D�c�N��d�I��8�<A֊��dx.��r�甔�̓\�m�t?0�AU�H=��.]N��>Ô�]d�BL�9[ �ȃ�JMpTk�ϩ�m�mkj�(��N���$����NK�(��u��.�*bjpiv�/����ڌ�����>��y[���H:�J]AW�A-�:�~��@��o$��T�8	W�C$���P�#�f!�'0�5�����"�t$z�tyq>֢*�n�4���h7KSU�@���T�D�0?
@���^�.{qf�|��C2;���{�	CՓ5�Q���C �#�#�
�	���NK%T�X��-���Y|�Lz?�0/�M��>�(z�3]����It#	��"şp>�Уwy���QS�x��I�:�K)E]�=�R��c���d��;:�^!A`����A��	��8�[��6��:6w��C�Hc���T=2���qF�pc�n!KN 3���Z������*b��rsK")�L�խF<�im�A�M�&�f����U�=r=#�>� �4�'�=�`9s�c�L0=����Ź��yӧ��@�R�E�
-�']�J�:AV��k�!�!�����<��9����MI��X�����? �4�#���j�}w�졨�e.$�2���N��aFjf��Q���IN%�r8�G�(�N��%{�p����H1ͬ�S�^����>\[}#�Z�!��Z
���½PU����L//�ۅ�vd"颹���+�S�D����&��6L��n:s�l�,N�X�!���E��"���ժnH$�v��v㐓��Ͽ%�FM�'SIG��>��ލ% ����d�h
Rڜ'G�z#�ǎϥ=����V8�yyA�"$E)t%�)~�z����7�Ƒ��i�x�{s�B�3ڛϤ��m�`5M���I2qf�.
	�$A��F9*���2��&��Ec�����O{ǹ�rp"@Y����Mg&��?}�4�:�x|Ig����rH�E���hH�aC�#"XN{��]���\r�.
_��7�*�֪]�G�L�� ��h����Iԃ�|L��|4ZV�q��8�ЁP�c���p]8u��	KXhtE�>�4����=�l*�uѬ`uy-�*�rd��!\3�Zj�������i�|��1/Nj��g�8CD�=Q�P�'�rbݴ��Ciފ��Ѩ�M`B��%��~UT�H&���?�~���34�I��3i���AmQG� /� ����=��i\�I)�˽������^:rD3���꣮ͩsVЙB=Rf&8��H/m�\��H�v��D~�$omy�],�[C �,ɫ{���"�qT�g�p||�4��a���ȋ��-	9 d1�@��J�� �3�?����ReI�K-ƖrQ�v{�ݻ�K����k+[���͖����i�ݲsm9�{$��?}.'�U�J�!(�fO�EQn�5�ݣɯЍ��:�Vp�hE����0	�=��9h�=T������� �3�TF ��8]إA GA�	�v	`�0J�V��q<j�����"y�WQ�\�.�z�=��У�>x�x"5��#��ҳ�6�mz��xh��=Se|��H'x0zB p��b�1uz��	���Z�ʠI6f��TN�&}~< ����ۏ��6�@�&&p�e�xzᲾu��> �*�O=��?j��]�WHc'U�v���}eԡ��L�ϰ[g��=�\m6E���h4�̪h\m`GÓ���R�:
B�N�Io�uQ�B�Pm��!ahM�25��=�x�!M��e�[W��+i������ԁ`A���,6�4N �w�kjj>:�� �a�����+� 4�P��յ���*�Q���ĴT2:���bY�.rQ �6�U��ZGQ�[�ʕ"�S���\1z�X�\���y$u�&P�d���Vӻ��=�b�4�N]d=�O<+Ȍ/]���z>��pc�x��f��m�#�+��o��)��rJ>��#y7Hl��2���h�ul�Tp{�'&͸�G�D޾};}��?�S�c��fϊ�E�Y8m�9�Ҩi�9\6���|G�0s�Ν<%g������G�2#�>;�� r�3q�ʺ.�z�sKl1��T��J�#�fx�m�~]	�/�L
8�.^�4r��hG�8�t"��_�d���Y|Eʳs��S�p�t<�9>x�c}Tc�=�䨣�P�^�\ ��_����ء+%��\��- ����_��l��Q�ƀK6��g��~>��G��ބ� ��P��-v%$r64xrQ��5�.���Z��h6��\�v��h���Sw��(��Fݦ�N�؂�B½V\��Ulb7/:�k/Ȍ�1��H���g������`iC23�V���կϰ ^oF��z�����p�e-��Y�gؗ�"�F��������s��,�n�mq ����+4a��sT%�����lîc����OV���>�E���Al8Ϙk<\W@s���Z�8�����f��IfIyA)�V��z0T�[�t���v�_����5_���!Y|F=74�B���*���p�ӄ�V����� !C���,>��;7ų�n�SyN8�e�����9y9@(8�4���|Զ7� ���D��[o�%)F�w^tN�j�î�+l��{����5dMm~��M��6���_})0�����O�Q�S����n| �K��pKT@�y�`��=�#�@s3rMi|\��M!��yGHF(e�;Q���L��5	�O@��
��0�����*�dQ@�sm����4�\�F$�{夡6ܙp>�R�9u5�}$����n�_q�<�Lwp�p��[�|�nw�P���J�<�M�!�
!����_̓�&QT�\��b��V��˗�uά�9����S��A*�� �<z9�fB�Q7l>�￿kq[lne��끷ű���\��i�nnaV짨I�MAxx1���������< �,6 o��8 ��iN�����ذ����9��@��I,8'���ӄ�,�`��L|�!�0��9+g��F$3Ȣ�{s�AW)y�%���a'pל�Ш���CM�s&� 5L����pN������:xF�)e�Lz)2H!�"\E�v������M��V�}�����l�5i��$�a9*�3�(?xV6������J3�õ<��ϼ�S�b�|'6�N0��q���>�Nw��w���m|n"���S�J�OvD��CR��	2����)���ka�ƮRl��hNӂ�0	���3 �BC6�����8\Y�$Z¨�)yeS�W&�A9�,��O1��O(^y����CѕK*[���m$��ƖlB*���=UF�j�B�2��a�p�Y�K��Ǌ4�Z�4MtE�Fk3��I��@�S�=�|=��\�������]��Fog5;��r���-1����;���T�V�|���4&'|��׊�����K��\c� 3�j�FGS^���%࣏>��������˗ӭ�7�� �$F@-���
Y�N�a��$_8�L�E8a��o����%���Q���g8��AC];��Dס��g�l����kb���n�e|��\�W*��������F�Օg(ї�h) �!�:��XF�i�/�a�W�H΄o��/�g�qd{UרENlہp���i���t�6����8}괌�][lN�@��S����O�ܧ�����<���٧Ϝ��l�)_\^Կ��k���u�%ZX2�~*��u2��28 Yp�S؆v�i�u�{�^z`�|��$kJ��]`���,����^l?������A	�_�w�*M��_&Uf�Y�HKӼ���Q/CS�����Wp���B� ~(�\��6�����v�*r�KRLZ���x@�\`N&�[0/��Ġ^������Цw�!�lC�<��`S�ښI�sO���q�,�-�In����l��^��io�-�rI�,���q��p�1�LBm��	CC�?��(�Q���Ι�C�J8+Q�b�(*k�R���x:H���tq���2Q:�A��#H�nv��т?~%�����=y�Q��|ԓ'��EqMM��ĺ��Ǥ��d�m��g�ׄ}��{:��m�Q��s�E�UR���L��]�/�	ʪΌ4��i�(<<(�S��ɷn�*&z�||��>�"�^�ԍH��{!���Ɔ8��>��)�GJm&0� Ţ�Kn�I+�c���e��A�ΐ8��^*�V��}���IH���h��(bG�H��&N~�SP�i��Rx�h&N%S7�}� �{	��yz�I��腖	��M��c���Ę�i�4�qTy����W����M���g��R}���pz�T���f�i���E'}���-[�b�!'�N���Ot�y���g[u��Բ��O�Q*��E
��{꼧���W��eXII0��o�������8��@}CI�!c�LTj�[���~�YL�?��ʩ�H��h��Nز6���2*��{�u�,\FU<Q��������cӽz8�Y����N�8!|M��	q�o��`U�
s�e7}����0$ �Dzp1�"�ܖ
a�Ο?��;?#��+A��J]�$&��ht\dj/�*t{�n$�,��-Er�����+ޒ�ͣ���l®���4��'�H�d�Nbc�Q�׾�N��@�sUH�d�K�*c㼯pd���'-õ��&�:�y�h����}w��*�m��������Iơ�(����p2L��P_�0j���@\�ԑ.!�駟�k׮�������X	C�$qp� $������7n(�ŽxHUjq&�A~8H�K�<0����}�$����H�����`�3�g��DGӜWW�<|���"?y�4�r�< ��T�6�~~��w��5PϷ���p��������ZGs8����7������$���>(^�G�C�J��-��հ'+�8J�|/cL�x�13�M��g�#���ykK�|��D���� Di���ϖ�x�7���&�R&��-��[�)ԀJM�Yr	��
h.)��V���$*�'�h�8m�NhE�g�xF�9�K�bC��d/��M���0i�(��Ln#\my�\ڧ�ȹՄӴ�#��{J��c�6����[�	��?�$�k�����	�-F�S�s}P�ۍq|�1�����k��7�rZ8x:�q��`:mۊA�P[���f��j1�7�dL�6�7�!��0T�3�Ϥ��%c�r��Y�!ۓ���s��y�vٔw.]�b�d4H|�d� *����9����7�o$�T�5��$Į<}�l�q�1ب$�M8q���d������I���\��W�H��$����_}-��
�Z;���`?�"�K�R�+��I�������D�S�CB�Y���W_}��L�9�EP��-\QT�Z�#[�=�X���sF��G7�M�io���M��p|]+�� �ǵ�Niׄ��/J�����3ʯD-87r&M���GJ"t(�G��7�^Hu����,<�|of�cPc�Q��nJ����&�Py���85�e3�Xd
~��_�yv��7|a��첻�[�t%q��=  '${0|�����F��'��!,h^�Mpv8gt�c#�z��[����'��d���ϊ8h/�����i�?�X*��o�}��ܠ�z�+�:y���$�H*����䑷G��:N���I�;�M��A�Q�>��]�!$���}|\]�N�7������K:�>�e�PK��|-@��bF:��&#|���3��Y3"�*v�UF�~`�pH8��l�`K�ௗ�މ�=T3��өre,^�w&`W�\��RWo9c�!,)��PY��}^�#[�S]yQ�#ܜ��$aH%7�^e�	9A����O{ܺs[z��YU������@A���=�e�sɕ�9/G��=�&Q�$}��>���؋�<���-�Z����r�9�˵X����͝���W�"U�O�6ւX<HR�,��J>��<�=�{��.ƾ 6��Q��?��2�B�-�/I���v4o޺^лR��P�*�x=nZ�Ň�4p`.�͛7�J*w��K�Y 6M���7��I��2�p���Q�Eu��SfՌ2^؋y���D�:�qVS����9�$A��3�k���L�cF(r��0����1�H--֜&�ʅ0R��Au�6ɕ�}����T0�������ϻ�+i�1�0��W�*�4C��K{&�e��
<�=B��c�=�^� D�C����>}�Lj��L�dʧ<{����&7b0���Q���h�ʌ�D��=|�H�#�O��{Y>pP�N*���� G��g'wռ;�.3�3�?�Uڞ��<��'�\9tPD0�·Mc8��8&����ܿ\��=a����س����8r�qv�/k�d���sX��U�6X���c�%&��2YT;�I0|/^T�N#�ۙ�H������s��9)Q��bE�*�t�T^��M����%O%mEFU�מ$$���#?��BЉ}��f��a��DANC6�"��!Ӏ���#u�!�-\6#WEmO��?q�-Ҫ����iDKH��)�Kl6�����(���W��2i�ِnEW�t����~�=n&y$)�M��6cU�AI��&��d<�-{���{�h��Ұ-�V��������!��qc!s��թmw����tR���s݌3��us}|0��@D���5�ϙ���k��D�,����#4+�Ÿ9����YR
��N,��k9}�y�pmlEn���#��r��!{��i4�{������	��F{0	��D���E�(��z j$�� v�	��~��N�,C٨EI�l�1�i�+c_��'��a�����.��X�qPo���g$5�`����T��p:����6#M��U˚�'u=N<P���;�R}I������u���A��盌�`s'H�G���&���y�̞Qt�z�4P'��kE�ή�Du���O>�D�AFU|�0����]\��,��Z�u�BF� ��-.�t�q��kZ����w@9OWoؕ>'AH��<[�f���"���C �P��h23�˝-ԼzZ�+��{���1�}9,@��r�K�s7�fP�;����A��Ov@�Ī	W6�R ���ے���=�u`.�<'=��vv>It$~��۷�Ҍd�	�N�����;�	/�F�z[1��A����Kj6�+-����IWQ{����pG9�
֎�Ho�H�����%K���[��U��-�A�f��س��^�!GG.I=sz�Nm�(��N3(̠h���.J�)�d�ƙMf�p��A�nn��N��&R��zSS�������M�Un�����%R�����U�͹����,<���==7���cE-��:���%5Iˤ�<��Y������2�����k������ٴjt�ζ�!v��՚>��|f'�Ae�h��DѠ]�X��̅d;���q�s�ޚ�]�M۶�NfyDk�I�'��c9X�����%zq2����H���c|d� ���u
���AT,*m]*XӼz6TJA�膌h׉W��9O��Ls�Y���7W�Sbt!I7�0l�w�'��}�⹂=R���!9.�'���8IO�7�fA�r�I� h��Ӿ�!�S�Tb��u�+�+�9�l��p��-Nx֑��S�J�ãv�|M��J�J)�h�X�q.��۽�\�0mǹ��s�[�h)���a��TI��]D�<uVL��*Αr�z�L���E�p�}m
=w� ���'e�H���Il��k{HM�����њ��q��`���~c��r�X�x8!It�����+Z ��b�9Y}�'+����!e�<PʝQ��X��*��=F�"��WH��?4�z��	�ؿF�9`�WK�JJ~j����uD%UN^,��a@��5�ɬ7HKƛ�f�Pq�R�頨�n0�B]?�l�%��n�u�'#̀b��q-��ی��N3��q���
�[�)l�5�ǌ+A)]��@Z����jFZ�� x��H�l���ٵp��z:����Y�B8_��E����Ɓ��l����gz�'R첳���"v��E|Y~�X�a�F#��Pp�&�O�zm]�{����H7�w�u1�ǜ�N_���q�`&#Y��C2(
)7�t nc�"s���k���U與8�|q�4��t:F]L� �L���;�v{˯I G���`�ݟ���\��<[Nڐ�����IA�V��|gFp1����h4~b�(��.�y{�zrrXA+T��jg(��H�H�:�d��=�sz(b$O;���Dj��xcS�#�� �R*7�"aWp)9�dQՏa��4����q.���h
�!��7�p� }V��쑰lI�R�x��$��) }"OhE����KA���=�I�0��M�G���8���B;�֋��f�2�]��Jo���/��o�ԋ�\Rb_�-i��FHDA%��N���S�\��t��a�r�����M�ίB�G٘k�|�4�������"Lm�H^^����Zz����5�*��X��u�.�S0):[{�|i^�L�G�niaob��k�6?��Tw8/
�K�ǳb?P����ic[�A��s[�j#�: �j�������H������.ʾá-*��x�Ç'rMِL��8�Uu��U`f�>x���y<3'���������;�4?�@�4`&R���͠����sH�A'x���i�R�B�t2�Y��C�)`����L{�v1�̳�I�4�v��*�y5q.8d��gL�7���ćy��+y��K��h�������Y�.^L����n_��>���ͫ&�)AE�h,>7��s�����͐��V��I\ޏ�˜��{�~��m�PrL( LSR����O� ���@mSD�����.3��N��c��h5�p�=sN��i����`e�]����[�YKE�}VS��ozo�
F*6Ա7}B,���Ey�ė��\����)$�]%V�xs��((�T	��֑�==�&6�Oj�t¼'$mqeQ@�ۦwŨ`�G�9�kN��/��f �X��ex�:��<�Y\|O|��=}&I�K��Q�]�}r�=sr�%�j�]q��Ncc�~��Ps�j��ŷ.:�M �1�d	��<�X�
e�xn����3R[RW�Z�{�&0G��C��t��Yi��3'I��if�p��f���0N���~��t@�"6�l��5����� sJ��s����d~�{�︱�2�S�^Q5N%�+N�(�l�޽򮮅Z:q��e�/ⴡ�H$��	@�������pb� 
h�3 bNx��'�\9�E -�ݲ6��ao8��z��N�s���`�-
EM}*��0@�۷n�4�|��J�q����~��󵪁�S :|�<D�l�}��]�0�nbG���G������3X��G��z��zˣ�I�y㺻�A|������n�=�z��{���O�M�ͷ_�+�^ѽ<y���ܩ�(-��%���8/[w��!	q�
dC�\27���ި�
������>Nb7◮�i���>����O~�S�����=��U�Gt6}��_���rp[�#�7gt<�Bb�?�G)��L����%�(N�5�i�x�â��B��u�E��&:)�4�&ɦ ֙� ��93c����>�  a,� �5��5!��8帹)��yr��ٵq>nݺ)!'euEBG.������[�\�e��^0�9fm��"R���ꪬb;J����q6F�ZH�S����8"O�!��J����B�O�{](7�w:=ى��C�ҽ����0��,0^��̙�EC�L�zEF8��E���wGa�Vp���G�H�G��L|��Lr��zk*ե@����;qx-A*����Δ�$�*6j-=�F"ٵJ�o�����=��C���)ӷ������溛���YI�͢^z�L��a����&w�.�f�u�f�O|���7�ҳ9�L�����'�n{&)�a ��h�}!�.)s����$)�m:�/)�^�9��p1�`N�&�Ta�Q�J��8B��5}��HjlS{]ѐ�L�h��������G|`��%�i[q��9�rsџ�ڕ=2U�]ٍfUx��l4�쫬�rZՒ�:�֞��b_`�y��x�����Q��	5�#I֗.�Kё76�@�o�9 lN7�#]n脲PM���J� ���.���p�����,"��o������?ӂ	Nc38ul�3�J��&�--4^Yb�-�a�@�����ƍ�z^�[�BR�s�"Ђ��¯mx�홝|l���@���'��x%�}�k'�7�F�BP�4z�S7�:6*�kBL��gQ4� .óHѩ���R/T9�D�ݖt���, ?O��r{�7*w�N[l�W�:R+������ը���ن�l�wD-��'�r/9������6��+a���qo�(���K��?ԏ{�ɟL�l�����辰aK������F�ðc�p[�?R����_UczCVY���kt%x���L�K--B��߸�>���鬸�2��(R3?�E#��c���˺6�1�ln��x�|�;<�y�Ҩ7Tʪ�+�*.M"����*�jѻ�*���s��U)��x���1h�����
Olg{���;;y'�e4��}T?��%'w&>��L�h����F$�\��OJ��K�>�U1��y}$	)Y��$����S|B�ѣ�1-����^U����G͜S�k�I1����yGۋ�/�@��%K�Z❸îEƕH��+��]}O�� �RT��{0�>�%�A�Aoee&������� ���g��箭y�C���f#��.TtNC�{�M���N-V���H�hxv<u�k�S��M�0�\4GTm!2l�D��m���.X,�_�&M�� �Q��u��6��u����E ��M��o�oJz�,�p6Ժ��%���ۗ�m�{�:k�*=�=v��/�-7�,�;w�9.�%���!�]��eù#ힹ���c>

g��wO(�N�D�gA]5͢M�����|'�r���-����h;�j8�TJ1!��p�|N|͙����2�\�&1�Hp3}���j2�:h' Fkl�=4Q7i�<_�Bՠ&�]=z�D�������m��PO����ay���$�u�㫯�V2��l���)�<�uX`��N��.�u��6������=�3�zMν�>|"}���ҵ��ub����*ZG͑�%{ґ�*�5�l��pb�;K��fy#�HF�M����8�}��M��3��y�JӒ�,ۻ2T��T��pЇ豦ւyuJ����Z��*�M ^���m�����0>�vqiA���9�O���C��C}.Xvhg��o ;f�w�����Vb��؁b�ٗ������ٰ5��~�$���u�p�p��#l��ZÜz��º!,>�\8!��:4M�����(ƃ�#p�IKωs)�M+k(�^��]�~CN݃���.�*�O�)�v��Q/]�f�͑#A��?tu��S��͡�Q,^N�Q8R��$��r����s�`����;õ���|�i�%<)�(:c�r�P.��h̉���\�oW����\v4�6A�-�>�r�lr�~gr�p{�`���,�O�\�4�_X���@��;����"2W���s.�O���3�泧�I�>t����Q$���m{�RH����J�Ϛ�����N�f6[��}Y�'д�`�_��xdK-msJ���'[�����A6�"�B"�xUcf�`��F�BO����Ltt��w��U���.�iő��7�B�J�������4�-eK9��!s� 7N)���
�0e��x>�\���ǜq�(.)RE���	'?�T�8�,�� -�n"ej2]]�g�;�-�;��`�0��35)X�3Sρ��x��l؜B��E%̓3C]ELwͦ�� w�U���� �If� 4�0Q�<h���ްWl@v��AP�7�� ����~����KaT�Z��7'���(�v��Y��q�b4��E�OY��ثgl�n�(N�g��'�[��A�6	 u�Be�k���a�.��R���*�*(�_�	ł��x�'�������zŖ�
�����}�88��XjJ��^�~�3�M��o���W4"8���b2���7��?�R�T�Q%�������L��5a|`Q2�.��p�*!@���q������I�;ܼn�k��M�S	�[�+rd��@��0�-_�A�ƒQ��,^�w��ݘY��x|����	!4���K�Еv}<,��8�^*��1|���A���|6�U�*�ٸ�{��m������S'��6o��UL��e�i>JH87C����,*A_'X��dj��~WYZ��)b�) �n�H��9�]k˂�{z=Ɩ�D��\�.���`wg]��S+�ή����e�1[k�Y3u�Zi~�I���g�@�0�:�4��{R�f�._9+��> �>�Z�i{nj-�U�
��+�7Ri;=�K��a�X#��"9a�~[�Z��ڽq\I3��x�l/�i��N��آ9:�o\s������uB�{1k��$���ܢ�#�K=a��'��yb�6�A�9,�apW1jl�����NH��cS��&���`Sh��X�cKi��R������뼺�������?��ȝ�=1��f��������93���}�5sR��J�J��}vG_�
�������gϜM�N[ƺJK����[R��ϊ:�nB���ك�w54rcmC�Ña@>g%یlC�9pa���
���ć���gC����(ꉈwu�ג@��B�:��tz���\B~$ے"w����,>��jp��z�o��Z����Pr>�,w�4��QO��Lh��w��5l#�7��8���	f��z�����G���~l�n��r��ܻ�@���˞	ʊ98&5uG%m0]�+�R���ͺ�<���߈Ld&B��{����eG��:���E7j�N_7������L��������|H���U����D���aqG�z��ё�؆���������\����?M_��$���w�}cj���X�#���~�D�.��u�f��m��8�����W���k�Ν[ⅼl��<%G��[n����3� ��onx����n�ϝ�%}�888#[��Z���`
p\v��i�J�k%����r
P0��vѻ��QaޤinaIFV����"��u��F쵽ae8��W�;�-"հ���#�-/_>W �ꀱ�������_�E���_�B����<�ٵ5���E=���׾5�q1�_����N?�u�:���j���`�q���XҨ��>�D5�e����Z��k��ܷ�����&���TQ�Kʮ9@lQ�O!R�Ӆ��N��uv��zUWz���<�"!	C�����1�N��I�����|I�G�������*N��v�;1��n�A� @h�hIw��d����yϽ��o�@���^{��z�:�:6�WD�3GeW���U�s���Ā�fr�b3"��b�^aӣ��$�MR���(���g�&�"j<3<�3g�v۔c����j�6�yR�+<�Υ��	��|��O��Y`��YW�w6���j*�$�;��I��vv��_����=�D^�yM bcv�7�hw-/i�P5�[�_�Jr��B:~�pV������ޅ��&1ʎ�6�K�HN�8 5��ڇ��lKww��6$H�T%pf:v�ί�p�uGjwy{�Z���T��8��$¾qsU2,�ѧj�Z;]�.,�0$|F�i6��� ��g�B�t�2�`��Y�,vs��N���qz�_~�g �q�e-��Ӵ��>��gA�97w�׳��y�������y1��ܓ��#8���C��Ս���M���/�������ͣ�j��
����^V���9�j�)/�ڇ�^L��F���r��O����V�\ͻ�Γ/�#v����'l�����&8�{��T.����/2��q|yv�UMZ��gtJh!f�V��Dh#�pF���8���9i#�Ct|������@P���I	���H��>I�!)��j>����_��<!f����=��8���z8����i�F� �be�J:��yU�Q?ۂ�������B���׾����L��~=}��SЈ�D ֳM�ti:�Q����QƩ( �ȁ���5�Y�i}�Mo����8�e5��d7��X��>R���˧_��O�����47����h�d��G���Sgi�������O��"kk�ɧ.���y��x��x!��=�#Yj�=�=�����N��ޗ�Ȣf�nfv>]�b8cN�h�N�A_I_�U���C�n���g�C�<�^�7��߼b�7?��lW�dU�o��Bz񥗅3���c"E�����~>TR�̙^z5;�<��1\l�4o���y�[x垍>rUe#Л��Z��P&6��EG�ƃ�aB��M�FXv�J��s1��撒5����$.�����4U�L11��ӿ˺wWF�, ����/��s�U:n����N���sMW8�7sI#�j A�%��q��^d6V�n��\�G��=��^^��,�粇DPz+{I���W��@�04����)�HT>�϶e#�Hfs��E	'pT������蠍�i�;iK^��+J#�.�4�������~�b��koO^	C�)aC�;�.���5'�1�O��[�P)��^oC� 3.bY���v&�]�TL�.l?�P��3O>����~�wrq��&!������H��vs�����9#T��xO������0Y"^�[��I ]C�pR#�/_KG����_��r)�����9sS��ЧN��w���G�B��eݺ�f�X��65ǫ-�)�,+T~�(�ې�2��3&e�����Q��4M`v�jP�^��{4��R�^`� �*��&j+�2�!O����s �D��f0Ⱦc��)���I|����[�;]^^4���'r���E�"���-�0���t4�Q9B���~�����.%���sS&��7�j�����O����*=��/������\�ҡEC��?pi]H���z:u�Io~5����yeg�ֽ5�S	��S�!�3�^V��)Z& �Q*~�H��?� Oi1��j@q^HJ�h�Ե,��`]L�Jm��7U�[�NU�S9\���o*�� w��i��t3���x�ߧ鹑�'F�7�C���a� m��ż�d �e��X�[�֕��]��"�
�w�y/=���g��m��mar-a�������'�Ns�3Ug�aM��Q��O#�Q��~;SE�]ؐ�(&��?��ڲMcF�q��G�t��~�ݬh�ٮ��>�(����8M�X�����Tvq��]��(u��ϟ�|](4|�~�����-#�4�z��k����.�3�y\�+xoY�N}��X'.fնF���|��(�4����8�	*���ګ����A��h�z�����X(�-��~��kJ����tV��}�s�^*����L��a�ޒ'�ĺ�
�e�x��T��@=���Ta�qkm�-b��7^��x�,*�5�f�呤M��ThSQQ���:I���X���M�s����度�q��.�_I���w���)��/|!=��s2�����t������i�}��i&K����WY�}�z����d��I#N8�7���\��!�r`�v ֙��~);����';	��{�=~�l)93b�	����]�� it��a&�^�n�Z'��S��mDd{�
�߆D
�&>�����8|��^<ʧ���ZH��}���=PT[��՗6�~���=LEm����Ϟ��AR��H�A�y��SD�z����hޟ=1�}�w��_����a)�T��B������Uf��=G����y��ϪB�d3�ŗ~�N��ռ��]z��3�<v�f`��#�s$>*�m��dUF��>w��f*k�\e���/�o���n��+�p�b�0�
���G?65u����!4@��1���qSJx9t�]G�����D>)Y��L�$5�����#��M���֙��4S�Uռ���ڣG�9:*�|��9�;�~���4(x�1�q���u�y�]vd�$5o���{l�/��2E�މ{�DI�5��_������U�vm*61��#����'*
��� ��Y�} 盳c�{Y�?!)���&��b"���pY[ۛ ��.�/������cGus��^U)�:�^�b�i��ܝ~%K]gbR�-�9O4���h�v>X�*�t�ұ{�W.�s+��o��N昨7Tj��/}%}��ǔ&���}/��ץ"���re�����jD��Le^��d���Dpԣ~��\��WO���� 1��⛢��ů�9}�U���ݪP�\� ��S"ٔ�{�[���7�-)%o��$SSm����ʨw��JZS[qR�UN
�}��4��,b�q�p{�>掜.*��Q�������`xj�Ȗ��f��q'!�d���b�X�dSi�/�߭Z�I��:��x7��ގ�0��~,���_~Y��g.2�.4����n�����CF ����R�b�qG�<�j���>�	q��m�8�+�ӵ�g�r�
��|�.y�F�14�n<VZ7f�$��w�&�T^95z�Pl��b[�����$4CU��z~��r`@e\��u39�/�4>��u�0k�8xSw�$A!�\���I'�\��*leWui��E!������K�G�c�*����n�-�΢2��i�fO��l��)�./l(ǅ�ԔAh9�9�ٹ�#�v�َ�)_�j�;Wx�|_���Y4"kl�~��l���FNO�`������i���k��3x:� Q5�،��-k�%Ŭ�����ݫڸ='D�Q�����W��=�|�sOʆ\�|U����P�o��N��#�K�K�Ig3ϼ������)�| ʅ�=���UU�rJJ"ٽ�~��AJ{��i�:ɿ�����;ޥ�W%���,d���OF���t�׷$�ׯh��k ԰��^5M4FKE��mF=() �n;	�zn�v�a�9О�J�߶aZ�
l�J�1O�o�9M�-H'�Ŝ��y�>�`z�D���N���p���ƠF�O�,My�IWЯRBnH��׽o-h�K��j��f
�Y�o
�j��RE����Moբ�tͥ|�.X�:�.��H�`�w����裏+��^���
g3q�� ��Z���~Q�}��׾�I �!˻fʾ�P9�,�Z}��d���B^��^5r��t]� T�Zȼ���;�v�,��|(�������kO��占��`���Ni(�KW���J�S�d��69��@��l��|���pY$pZ��Ͽ�m�?�3o��BvC6ϲ9�sם�"5��0��ݔ�1�0P#F���<���a�T׳*k; J<?����!��4f
�<C��v�H�g�䝷n'�2�B���A�/�Ҷ�|]YǑ������ZבGj�l~��GU�?����H/H���Y���彲Pl��mt�����/9G�O�gdcs����B��1?���2H�fm�aVm���� Z-������=;=�S�����/�g��S	�M���Oq�(���f�ī�&���4
=Ć�?C��0���X3����+�k<��y'��B�ǔ��Y����:��)`��d N'����T����Ϳ�=^z�e�| Ck�j��:�=ɽAٓ;�MY^X�����g9ZV�s��PCaTϠ�O=������H� �Vl�Z��f���q�Q&g�eCٌ�����i�қ�G�Yx'� ^&�Fj4xo�֨T��=vyI 1q���r�*�ɕ�=L�9 ?G���B�ڸ;�09)�I�&@e��$�2w�qb,*v�jH}p]x߱+����|⊶AhhJ���	<*6���7��y8g��,��,t
�vr2;ׯd�.c*=�������埾�^y�%B1�$;������.\�y~�l�3����<&p7v� ����D2��!����YqH�YP�k����(���rhӇM
Q�|ĈɄ�]�y�\��@��>D�⯽qC:<�.�ay�I]�{qʈ�I^�5��Og���̌b�(-hH�^���v�;48��=��x�sUS�:�F���5�SD��.?��C�mP�T� L�/��^�ɋ�^)�'���2�P�L�q���o�� ,y�9em��EU�u��HB`b�P�˱Aw/+U�E����Դ��#�l+�����'c���[��	Ժ�f��H��!��3�9h��^!]o���L�Y��Ii���x�8w���g�{��� T-������6niW������;꺑oh�n��	i��o}K(j�4j�h4��&�n�!�-`�N�|@�TЙd3x {S�k�s4:ن��7�V�OV�8c��;>!q@H��+�ӱ�1�;��.ZvI�`��=��}+m�E^��ZZ�N�0؄Xd^,��䯺=������`�/Xֹ%�L���e �)���1��Z���$�>6�nB��axE���hW�^J�m�@ǽ�����\p�=u�1�Aj� @���/n�r~6�V
��%C)"�8=��h�+)3��r�-�a�|�g-W��f��p}V*�159m�]N�w��D��XHp�4�QqY�j�4/E�"�G��͢'��Ǣ�^������5Eg���9�G�BO6Ӈ�SC ���B$58�W�ʍfK�U��F�K���x��z8obKe`ZӠP�𞬹f��N��=��x^~f7�sg�B#pF�yB���+����%�Y�|�9F����Dvw��8d�2"_"Y�HS�)7�6l�4B�͋A�#h��G��E���X*��KblqyH�kH�2[6o:�<
E��9eؒ�I9�&��7��nN�~Z�&>�J�����VxW�5�H����8ZvEńK|A�"*È������� �VF8������r�����MK���0�6ڷQ�Ua*�n��ڏ�6��ٙY��XW>��]G�:/�=����J��&x6�����5���=r�Ps�($	�ـ�ѓZ�MԼ��u�8R
��vD�m�`� �������Ԇ�a����c�2��'��3�{mH��`"l�����9;����]�Pޟm�ة�u���M��8x�\�`XP�AO6����~��RgY9!�RD�N�g�*�Wm����j�ɟ)p�$�H�е\A�st�H��'��G?91���7+ra���-��M� J���:�5���&�8+v� </:Ɣ�A����3K�%ӳ&\�J�lZ���q�)~���jT%�j��i:$yI����YJp��ά�DhM�������3s�)�6�c�`q�����Os�@��E�&�G�jZ����<��fvcNhH�ɓ�˰��*�<'�FT�f]�m���$���M�hbC����V�B`|):q�5�"���̾ʞ�z�,�.���bhQY��2�]̟a4��"�߳����V�΋$f�w@^��2���Y��p��~v��H�_`f
em*�����@C�m�[���h��,�V��� �L΁��0�&$�N�K�b`�B��c�t���i2�"�)�(𫨟�H�a#�.y6�
���A�r��T3/�u��U���CRK��ˆqM#X+}N�ا��@:���Re|�~ޑ��G���|����暢n��Ն��R�\s�h���+��(�7?�8�?D�Gr,F?��O����ny�'/�OG��"���	H�䭿�
�m�[��RO��s�}\�=��]^8ҹ6Eƺl��,yF�.F2QO�W�uwRܤ�A��Rxnj�(G2� "yIlX�b =��m����6]���ިf�X��^E"��r�tgR@�M]G�F�fÏ���6،g���I�jW�=T�R6X ��l�/���ᗻ������z��8��k��U��d�����߉�Qa�`��uv���q[���U�r���/О��2�����3�= ?}�דtF��ɓ3>�}���<ڔm��1ݟl )N"��1�� c~���v%8m�!�PBa{�7l��h��#�r�k� 5V�j��n�����]�H��؄�9�$�#O�������u��!� �G��f��t$�S�����G�x��wk-��fH�+��{�%<��M��2���Άp��C���B�zF�P)�!�����o�a�_��O�%�Ϟ���HF��sx����C��w�dh6J�{�r{+��2fd7>9����Ʋ�+ҙ���H�eQ09cҊ����h�����x2_�$�tPU�S�\^<K��hs#=c|v�`z�}�jq�M���^�~F�A�8p/rʐx�������������kZ��Y�zW���R#���C��0��R��k�G��kC�l�ۣ��Ȯ=�F��]T9#�5P��ZbQ�,\�ʎ�:��r�����Rk���q�gZ���-��^5��^����q�:�%�+G����}A-�߀&$��n�[�1����{�/�������H]�N���i{e;�fg{ۇ�,9�_�����$aC�sJ��w��7R:�MZ ;�0��?�6;~�� �^���N�e��֋qRa�wސ���L�p4�#m�׉i;{�����lז5R1�PsG��|�i�jzvZ�\i�6E�eۻTA��mv���2�� �Ɵ4��F�Pc8!���*J&�ŽAHb�����j�80v,���|JN�_�g���-E�s��?�0b4�k�>&�SD2�� �����a��H8mB�4uBj��٨��	����:gb�Դ���v�Mmm���T�L��\Aw�)X��Ń�M+, �o`�\7T_ ���t�
XP�A؛��XR渭!/NXF C����`pJ��k$�</�b���mm2]�l����~���u	{p]���qb�F4#{0ǰ�)Ù�y���N�6�������0fsɓ�l�@/V���U�g�"J4NOI��߶��ㆴᚢf�|���]��!�N���]�|���m��m�!=\�"��]V��m�NnF'�2<�)|W���QU,<)���^��(����]��J�	@��iTjSj���*>9;�T%��C#�4/p���H���g��@ᡞɼ1�*�S�4,������SY�ƖCj���F`{����%�� �3�z8�[cG+L�Mb�/h<�$QAc�[�sy�I�@߭&.cw�7t⢮��1X$5d:�P�/OS��R�X}#b���r��k��6��p?5d��M���m��"?�F6h�77�U5�S�)A�o ��B������M>�p��s]�2�Ե���,d 1X��򉊋�ρ��mJ�)��V���I����э����u�^��7�?t�yf�P��Y(����=�.��,���g�����Ą�
+v-G�R�������2Ww0��}��mh��*zYļ�&�:�w�����Ĝv�4��(��76o{�J�܏MA��ݽm��zR�M	M*�]bRji��a��#�O��tBJ����p���w81YD"nz;4��$��;�_0�5��}%��;Ө얌�
NM�;jE�n�Ԉ��q��iP��h�f~�E��h���X����q�7��q�Q"j6�R2�{��֟���>�J*��(�-���7���fώ�D�2L�/F[�~ii!V��3ڀ8Q�����; =�i����Мu4"g��`�����-�~�
^ר��(\�CΗk���"U���������ѭ;�j����CQ�hZ�ں��(V���=�Th6��Q�F���3�9{����5v����E"�]�q�+�o��|%�g�i�z6�@G�|���$w�m&��?yD���Ysx�
���j=r��qvAً�A�n�M�Pgv���6���d��r*f�#u�(0�$٘ �]��5/����C�瓺z��`�G��īa}v7z7*#��mx����Wll7d��t^��f��� ���5��>{2�l� $5��Q��IMQc�T%.,%6��m�0VVAd�9�J��L���y�}�A�Z�ъ�4:ޡ��60IX��<<��0�D6I;Udf"륂�p�	x��wD��i�Y�PC��l��4(m�ٛB��(8�H�؛� �2����I��֝;%�6������ AW���7מ��d8�sb�i8�W� rL�vNK�;����"p�5����坔���G?�sh ���մriE�+6�g��Ϥ�Fz/M:%@�W���F���}A�#�{ާ^:H��S_ �G�p�����Q}X6Ed�RCVGfXD6���,іt{]�skÈk���4�&�f�$6A6e��}�9�p�2�g����F��m7��eH^�)����*[�n�I	h$:V5�s]�ɚa7x�M߁�
���)���6�Z��mf3=��#:�*ߪU���R6cR'��Qw^�9���c���T�4&>��Ӣ�
|��<��s��T��[�[��>��+�!�H��w��Б�������C���o����&��Jc���
9襉�ImK2��/�inn�G�N�ԅl5:�	�\���Q*�?����*Y8�lR|�g��4�ܚ7y~�IYfc�\�w|��Al��?��z��U��u�$�ϘX��ߍ����n�"��U�$��c�[ؓhn��mڼ�Kl��0D�����mw5��b�^�ͫ�D��ZP
��.m+�ܑ�P��n��k�+����$�*f��1r5��w=5�Q;B��>�j=սMM�"�ü~�w�pqEj�����G�e��b����6��ʠ���U��Ơ�j�����j��8	�&�T� �������0u�'=��ea���ţ̽ex0s; >J�I�|���Ȣ#}e2����-��t�X�FUb.�/�ܪ��Os�g�G����R�+(���Y�mM�1N�N'�� �N��G'�'J����L��j=�ZU��}�i�P��.74&�8�=��� m�?�� ��D�x� ��7��h����NvÆ�t"-���܋Z�f�*�!��Ѡ7*��RY��{5�JuD�Px� �o�QGWKj��Г�����R�]-*�\�Fs���5Yh�J(�Yi�(�Յ'��>f���!�S�jgcC����g�t�����<\m������u��N���i�Ջj-mûrJP�a\Q���YX�z���z�4jf��:6�1$��5��LN��}��N-��}y��h8:U�J�|�v7�7��v����5(�V%$�~Y��`U�6#�F��چ���i+A�CxN��/��|}y�����,ÊGjO��=yH[��)���s�.b׶���P��In��R�D@f��4*�b�yVbK]���{c�U%��F� �)Oɪ���^��F.�p4V��5������O����_4�0�$c���S��(�e9p���w���[r�q����AE�2L�BW)�8�3n��i9�p�{��嘬����J�t�sD�8"hk�Ɉ���o4���)�jH�X|FN3m؁����ưu+ �b̷�@���/Y��У��W�9%;�='������g���`�H�3P����:�h�z�����j�:X���.���~�F�����*1��Aa��7��
D����da�'��n�2Ζ���>'(R�:�>�.�_}����e���u�O	��������";v�}_3��X���"(i*x��U�+�\�6U����nLG��6��V���,��s���k�/OPJJ�k�y��	��w}6	P	M*ܞYu4l˄��M�{=�_�0Q95^���d�Gs8�^W1�{"Q��ؠW���pb���m;����K^�lVO�mT��S� 8d�m�­�����M�te�v|@�I��'��4��V(���(#�B����"~l�-R�]ؾ}�дwl�d��@.��~7�r��R�%��}a�����Q� �5q6ʱ ׽��>�� �;a��m�>��Z}{�H��	��Uގ��M���u�D��~,��\�E��z�>Xxd�t�Z�G��[�M7£���Hd/���B�4To�P��x7٬�3�z�+$n-iTѸ��pz�9�=TQ����p�tp3�36��Y�n�V��ꧥ�O�Ƒ��@���@��nM��#�"2_��py9PI^�1�a�6
�=����T���o���WPYt�d�ʚ�-}��ʍfur��#�: ���޶׾w��D߽f�2�q�r�cݚ���Z�g����*4w�!w:6w��W 8>���`>9{Y�F=���M��Ƣ��rM=��d�����-b奆#�u8Ђu����+}�B����9p+j�dc�9
�/�Qc٩��:���)�)��� Y�@�8h�Z����"�t*�@��	)*�OQe��i���b��c�7ڕAj�m�q���	�����J���ӕ7��j�o�*�� �f�-qh6ʒo}?��Xr�}Fa]E��N��T��H�X[uO�S�96����*���F��1V��-�B�Z�99ʊ\�fmdT1.8ݮ��r��Sk�#T��oH�����=�(�l'�6ia��wD�mSЌ�!�;FZ����|�,���Y-�F�v��hY#�y6�R��1�6�6$��֤!w6��J�GG��M����&���k檛�6�P)|�`د��P��p$�MsqU�7F̎�u{QZ�T�2��6��~��ؔ8)�&�J�YM�����y��ݪy��UF!g�{PZ;ND�"����
���L�傶��"����@i��yK܅�Hfy49��H���ć�	充��Q �؋�m�����j�T&�~�}��0�SR�)�i��I��G��*�}TD��F2��UU7��{���<�._�,����;h�|�i��&1�J
�{�֌����B�/fy����փ��	�(�Bhz���G���Zt��&��s]@%��C�,��>x:u�T~���P6����>>c�h؎�ߔ�mz����P�����oR���N��'� �5kj�xR���L����=N�	{
�J�T.x=5Q�.�l�a}3R���RޮWO���/�\�ɴ^�V -�~������ee�LIZ)�~��'���q�hd�c�A�	غͨ�Z��>w���~U�K����D����u����mSw]��� ,3ސAe���"�M�k���7&<�ؤHQ���'|R�~�sMj�3ڳ����[�'���2D�$�1��������>���'5[�6�OT��}��X�˚{<��'�==w�cC�߷���pWKF��_�Ro,T}C����lc��=�kۛRu�-����]O�F������~i�}C>�;�!��]~Ԗ��΢��z��5�SW��������7�����t���3��<i�aޯ�M���cI"������̦|䆘�{]�oH��d|���-w9�e��rI�r_4�=x�o�%�鄌b����Z�S��G�3@2�>S�_ڲE��^F�ُ=%��R��z<r�k�X�(�X%�Dc/Ζ��ޯg��'��U������O�mu�;�J�¹���I���*^�c�FUb�Q�޽�>�iS>vC"Zϫ�?�DDa�٨Ƌ4��|;���f�Ft�5�kσ�Q�s�2������L�~�������z�#��q��;0ݿ���|��	i�b�۔E�?�}�anĝ���y�RQ�Oe���[������������8e�����>�l�M5��;]��<������	]1X�Bi�    IEND�B`�PK
     mdZ�&�y`  y`  /   images/8c2f1315-cf23-4ba8-a920-becb97f13280.png�PNG

   IHDR  �  �   ��ߊ  NiCCPicc  (�c``RI,(�aa``��+)
rwR���R`����b
����>@%0|����/��:%5�I�^��b��Ջ�D�0գ ����d ��S��JS�l����):
Ȟb�C�@�$�XMH�3�}�VH�H�����IBOGbC�n��ₜ�J� c�%��V��h���ʢ��G`(�*x�%��(�30����s 8,�� Ě�30������n���~��@�\;b��'v$%�����)-����r�H�@=��i�F`yF'�{��Vc``����w�������w1P��y !e��?C    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs  %  %IR$�   tIME�WxG  �zTXtRaw profile type icc  8��S[n�0��)z^�8~$R��b;^eWݪ��HQb�0$|�>�� D�h`�dZ@�&F�Ąb�9��m��P=Eec������O8��`��Й�f�
�Q�A:���{�xt�k��7�����������-eP/���\!�����jS�u�mۃ��Qa;��B�["�,FدCl֤�	�����/�&�S�T�c��\���~�y�_���D6:J&�D�z����f5u�R�����Ye:�010�����?1:9�����{��5nH����^υZ�w�R��WU(5G�Ӫu2j�fo�-���)�:&c*+q�y&�"J��G��|/��d�c?&s&]����VG��^q���@����줁/0�   orNTϢw�  [5IDATx���w|e���3[�����!�XQ�	6�g׻��;�ӟ�SO�]�Slxީ��)6Գ��^C��m7����cӳ��؅|ޯ����y����S�y """"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""�P �t뎇yX��s*�+��������L����>����<�r�ݵ/�ϯj>��ߌ�	�\51�;Z�w�e[�L�>��( ��R�	�NUo��W{��v��	댍
�_�f�|����Io[����7�9	s� W�>����&A����@��H��t@U���"^ n@U���^}z/[�j�[�*)9����n͚?VTV����� �*�, 4 ��{!��yLDDtX2�I�+�|���5]�dݸy����S�NMX�˯����^!"Z�SNDDDው�]8|�+LUU�S�
�n�u=&҉"""�����]bc�L������H'����ZND��fK�<�M��DDD p�ݚf���*(w��CDDD��%�$ϷX��'0���������p��a���ʓ<���#������	E��Qn������iӶ/[�lBaaAV�`�Դ48��vX�6�-fh�	�R�4J)(�L�O""":t��r�];���T�r:��'O�����z��:<7<O�����F�ۍ��*����v����"�_A��jf"��r�|��������Z�����=v�m����X5z4LZx�Ͱ�����QCrTAii)~[�+¹1k���e�E���;���^�&���� ""��:Z،m�tV��r�}^_��✕Nx�^�m�H�Q�6�5�_�6���At�z�^{�7].��#�WDDD������[u�ޤ�r9�q{"�F"""j����"b�-��t:]p{8�Q��JJK��x��.��o�\.x<,�E9�

�i*^=x@w��NDD��VPX �������}U�z<p�\�N'5C++)���r��~S�7}>*++#�F"""j� n��&"M����|��`@'""�f
�����D����>�,�E5AM	��������r��t:���(4��r� Ȉx>�N�3҉$""�������3ƌm��.�x��N%�������/ �y9�9Q���M������NDD�4 PJٍ�������(��@([�6t �z}0z������h 4��^�����(�i�ee����h�����(�iK�-W*D@�1�E=m����R�b� �Љ�����_�� t�"A��#""����+ �ϡ�ʝ��(�VZV��H�*w/D�H'����B�*�˕@LFx}>��NDD��VQY�D�Y�NDD����
��q@���;Q��*]N��!��%t�t""�h%М��J�u�h_u�8>�FDD��9�����_g/w""�h�UU���S�����G:�DDDdD��j5���~?K�DDDQK ��p�tݯCg�;Q4�b��b�W]t�)���(�i�����]��:QT�L���]ס�|
���(�i��LP�0��܉������2�fJ�r'""�j�)(���ua�;Q��bR
!:�܉���� �DD���ʝ��(�iգ�i0�OM�r'""�v͖�u]X�NDD��u*��^]B��܉����V=u��-�p`""��&uݸ�΁e������h~����*w""�����z���*w""��%���u%Ͷ���NDD�4�߯A� �+�C�)���(�i�߯��ϡE9i��5v�#""�~���J`\�.�NqDDD�N��	�)NNDD��l6[�����DDDQ�l65�`@oW�3[j^���&��Q ""#f��dX�~0�d������%سgv�؅��TTT������PJ�n�!11�������dt���D��@��!"�:��i!K�pr�V��"((,Ěu��ӏ?a�����ۊ����^�'��P�Q�4M�f��EJj*�w�#�c���5j��2a�4v":�(���fM�̡2N �ro!���b�ڵ���O���o�v�Z@��hI��� �z������ck�f,��������ӦM������b6��'�#�P\Z
�łX�#��9|Ĭ�BV�C�ϡ�I��x�d�R�=�m|�ɧض5��Q��V����TT�c�o��t����o�����_���{�]-��O7���������Wa�QG��f���x�� ��ZM�mݶ/�y�y��صk'�5�촭ܚ��-�7���Ǘ�č�wfL����/ 6j���m؀_|	�����xp�e�F:i�10�\�˄� ��n|��x�����Ͽ���"�U�&-��]��ۢ_񧫯��͛q�5� 1>�A����PXT�w�{���?�r�
��Gjj:T���d�B�*w�U����r�~�<��S((؏�L�Z���jVb��d�ɤA�4�������!�/�fK!��PX���gݏ��"�|�M蔖ƠNDQ������3�������rV�u!�a���|�8������x����sꝌ0�@n�� 33]�vEnn.�v���D���#&&�*������ �6m�m�6��
?Ȫ�ବ��g�����w/:��3�Q�Q �-[���x6oڈ��/��̀�B����F�}��nǿ��:�^�O�@�edfb�ر�:u
Ǝ���,$$$�j6n�p��(..ƪի��O�����c���5&������ks�"�S:��v8�vu"�:%�%ؿ?����p�Y X�6��҉G}���u��g��Ĥd�:}:���J�1	qq��6�|o�n�!+#Y�p�	���+0g��{�-��0�{=x���w�޸䒋�)~Y�(�(@)��ۋ �D��*wv������չs1�9�s��Q�����s�>��;	qquü����e�&3��G~�>�,r��G]{c
�Ņx���p�B��u ���B��.|l����7��ByY	�s�f2a���x��p��� !>�EA܈ ���p��31���2tx��jؼi#�{�y�UTD:눈�Q  ����]�*w���������];���t9M3��s��3�>��C��K ��f]O���z]�u�qI��g��o�e)�����.��8"�����ޚ��.@m$�q�L��Y�݋�99�3� �8�d���<1P(.*�K/����Bu"�#�D�5����EX�n^|�%���^��c�!�u�,������,7i.��bL�6-d������H��!!DBv3L�ڱK����[�0��<66�˵1l�!{LL $'&��+�D��0*�������?���9�te�:��}8��)R��ys$���~P`��f����+ ;v��']��(�O�<g�uVD��;f��8��S���/5M�����? /o+���m��������z�v���z f�6�V�f��v���G��4x?����|�=p{�����X,�Z��Y�0�L����zo��v��vCD`��`�X`�Xj�o��
��p������v�����������
Ku��6���������vC=��f��6��+_�Q�ן9p����z���`2�`�Xa�Ya�X`�~\���,=F�S�3: ������]�����f�ߚydMi��7"�^@��U�_�V�Z�S+1)_r1R����& 118k�x���QR\��H.5Kh8p� V�\�n�f��}{�b��X�n6oڄ�{������j�"..�ѣ����!''16[�>����rTVV6���dBJr2̍���/,Ě5k�d�lX��w�Fee%|>lV���е[W���#F�@�~����Т������k�d��[�{���鄈��p >>9�9:|��>�{#.6���T^Q�����u��vj����dX-���+*.����d�R�[�;w�Dee%�^o���ƢKv6r��b�0` R��[�6���k׮��ŋ�n�:�ڵ�������|��CVV6C�A߾}���|iN�M� (-+�֭[�v�Z�[�۷oGA~>\UU�z�0�͈�ۑ����]����4p z�쁄��v�ٯ��BIii��RHLH�#&&h^Wy<عs'V�\�իVa˖-�?�W�~�V�������Fnn.�����#==�6/Z���N���w�Ʉ��"��_]�QPX�������M�w8HHH`MBCR�C�r�ϡ+ e��OPU�Q�|���8��qM�Q�0t�|��(�!.>���ӷ/��!C�b�ر�r�]\R�_~]�O?�?��3�mۆ��2��kf�b��%;cǎ��iSq��ǣszzuN���:^y�U��ƛ��PA�Ν�ēO�wϞJ8�v��ǟ|�w�}�V�DaaQ��P0���ԩF�9
^x!N9eb��pj��{�|��gx�w�b�
VO��SV��;w±��/��=��9�Σw�}s^x���"���D<���Z�DFM��8����s���;X�t)
��k���43R��0b�\p��6m*R���-��������罍%K��� ��x;�iiiw�Ѹ���a' 1!�uU�G[�m���_�/���e�q����\}�j��l�Թ3����S�`ҤSЭk�6��*����#f�{����T�Z����o���hpL�UU���_���a���c�8++�)�dAJr2�)S�bƌ��ۧL��>��~̞�>��chZu�Q@iI	����$)�����nGBBB���u]�̙3q���T�� 6�M3�y)���7����DDV�Z%�{��~��i��Vy⩧#�?~]�9/�,g�s������g�Ɇ�����\��{Ӷ��p:�O>���8S��S덑�Ο��T����䤓O���������9�~�����������EV�ZU�Ϊ*y���O�-���XgBb�\vŕ�a㦠i�r{��O?�'�$�Vn'5-]���u�c��V��?�4_�R�����+���RN�<Ebbb[��������s�=_��\ix.y|>���2����kU�$&%˥�_!6mn���{��ǟ��#F��jk��^w�[m12�����?�)

DD�_�jm��x�z�.���9/6ȓ�k��5��t�Y/]-���"�ǞxR��燝��W.�����_8�9���Z<^o�cġ��������W�$&&�Đaß�L����y#�+R���_��ax�euɑ��GE���n�t��oi�t���߸Q�t�%%-�A<�">1I.��R� ~@��_��[��A�dw���V��H~a��q�ݒ�֩Z�~e�&�,�W�j��""%ee���K猬�������-r��dͺu�:���w�(ej���4��O?զ��G�̬�6c%���c�ʏ���$_*�Ny��$�k�6oGi&9a�I�h�v;�}~�|�ͷ2q�d�Z�m<v�C{L��v�Y���E��5�|s޼ꛮ���ify�ŗD�����s5zL�s�m�`���9�] �6l+�=^�\z��횏W]�'��}��|������?Q������UW�)DfBN>e�E]���b�����o����
���ߖ� �9J>��3���%��^�F��W]]�d�%��N�m;vH������n�#��n~�9���d߁�KG���Y�����n�Y���z��q�v���|)���{�%	���S&O����IgU��0�E�V�V.� ��<΁�,���x}�V�Y$t@����""��[�k���u��)S��漼f�π~hzBb��'���) ���X�|E��4�5
I���3\8�o+]�	���j����h�2�>�'PJ�j��j�C�����߭²%���k����~��#L{�R
%�������˯�����뽤�>5�9�K�����|�p&�y��g�tVɳ�o磏>ċ/�����������O<�gf?ge�i�k�O_Kҫ���O=�J�n��=�O<��#(+-#���?�v���k<��l���V���³�<�[n�۷�ե�����Vs�����f��>��Ar���5����Ǜo��nǲ�O?���|vl�Z�/�Ϥ���`�5T�����<���t����ԍe�7z�����c��
�Z.ս�Us1��d^}���طo���v���T����	۟17�p#�6oBM�4���cࠁ9r��� %%�����{����e˰r�J�߿��3X�sN��my����a��q�駵S/V�߇���:�x����n>�c��ХK6z��.�]�*W�����u�VT��:F*�~/��70}�t�\�
�̞�*���vLGl<r��W�^HOOG||<\.v�؉u��a���՝Ϥ�qW������8���o{GB����x�w�rU6�?&�YY��ݻr�� !!n�شi�l1�	@M�2����8��3P\\�G~�����=Ɓ��������HLH�����]��~�z�ܱ>��4źߋyo��̙31n�Q-��χ�^~�f݇Ғ"��:�q�ӧ/F��A�!5-q��p�\(,,D^^.\�u�֡���^fԧa��������O?��G�^�+��+V��9/4� p��!;�z�쉴�t$&&����@����!o�����=�7?�}�]L�>S&�2=�z���Q��i��z�oټ~_��ٌ�}� !>�i�8�ѣG�ꎀTK <d�ˡ�ܭ�yu�kQW�|�_""��J�R�� ��]��E�qy#"�l�
>rt3U=��N��?]#��^�
���Kc~]���b��_�o7��dee7S=	�?`����/-�[�*wM�[u�w���b���㏑'gϖ�+WIqI��=��|��z���R6m�,�ϙ#Æ�Y�e2Yd��iҳw�F���O��N?S�xk�lشY�+*l���T/]&��q���t�?&�U~��v�r�+P��0_Lf��5Z|�Y�t�KU��V�\��m�����2n�1�4S��*M�Lr�Ie����|Qu�㈓I������%kׯ�����RZ^.+V��Y�= �z�}�(��|�m���Z|ο�����_�?q����k�u��r�%��'���?�DN;��z�����������q��R&INN���uHjZ'9��d������������|�t�d�Ν��G˹�/�	I�^�:�).-5L�_MP����{���={e���7ߒ��� �TIrr�����o���g�����҈_'U��_­rOHZ��C��2�[��ʫs����楗_��fx"6\v��uD午HQq��w��m<�����O?�J���bj�""UOu��)�e����8M���v��
����j����Y��n�^�{<�>Էd�r9���͗���ӷ����\)*.iv;^�O���2h�Аy3ᤓ���(�1
���%1)E���FٴeK���˺d��[��$�kwyj�3�?���|��|���d̸�C�ˈQ�e���a狈���;��ԴN��{�!���m�\�����By��g�i�V2��0��)bЛSM4�E�?a�|��gRVQ��^RV&/��buڍ:�)霑)?���;��_~)���Azjj�|���I(��VFe@4x����^y��d`mF����;���I��������W_{Mb�/�J3ɔi�ʪ�k[��""�����s����Dd�G{\���N��E(K^z�U��x������V��s�ꐡ�F�7�~>��|�駒��E�j��v�!�W�{��z]�$����O>U{�nz��Xz����Ss���ǟ��脻��� =z�6؎�������~{��*�\w��B��Kv��2�5qU��[r�麼�����|�8y�ŗZ�
��,\��?ʖ�[�F���뺼��[ҩ�q����Ly��k�9�u>~u������8�����C-�˴��T]�;ŉ�����:nt��	�6�m��{�⥗^FeE�&��0�$<���n� �z����>���f���
��}6nl�����o���a�X��p���>}zXKgfu�=��N8����:e�D�v�ü)(����[�-W �l�⪫��UW���E�2b�p�}��P���>�)�����1c���Z0@� 8��8�����PRR�6��>�ſ�ݷ߁H��i�Ĥ�~���a�Z[tk�z1)�3�8<� :gd��5E���ܹs�s׮��Li�y�L�ݤQ�^����:�L\r�%PZ�c�������QYY����tPi����,p�W����LJr2,Cf����,]�zZ������v+���ݦ�5;��~+����k׮Ň~�E('�|.��RX�ՊI�&!>>�B���p�e�a�)���ՊSN����S�*T���eK{tcǍ��W�16[���I�p�ĉHMKCs=��=�\�}��V.��a�ē���t;^��7o�?���U�|�-�޽��wM3���/�%_sn<�	�g�v���
��֠��t�̟�em�ӑ��7�x:��55�%i�Z,8��sеk�n�桰��]RM��iF�]�H������^�Fb�#��eYE>��C��A߷Xm�����;���_#G��u�]�#�.c�ߋO>����k��� .>]t�SS[�@VV�/�:�v놙3ς�ln�vrs�"-=x��u?���ۜ#5�b����.@���V��O�>�޽[�|t��s�;���k �ٳ'��2�#(..��o�͛7�/�2X�����_	GLL���V��^z	�`�tw��~�	J��ڥ��4Κ9�n�q�>}0d�P��K��Q^V����@4MӚ-��,�+ >�����餶�>o޼K/1XBG߾}q�9g7���-���N��#G���5�VW����_�~?��6�%=-�YY!�9���ѿ�6m'%9ii��RQQVI4�|�ޣ;&L8�MkINJBN׮!�3f���)�@bB:w�l�LEE�z�!�����m��tn2Yp���!77�ݚ�@�=0��i�M���8�&��֩SgL�2fMk�Ͱ �����`�[e����+���n�t́et�������v�M�h�"�ݻ���5�<q"zT�õ�ѹ3N�~�aUdYY~���v	^�G�F�N��Plv;:g�يѣG���>�ݎ��$�������|�0�aÆ!��s`�X���a���0rԨ�Y�ZC!0�_rrJ�|q���1�� 2?��#��`������ĉk�@m/&MÄ	�����7������Ö�����>�+jJ�k׮0����|>����5���DS��b��9}��d��zz�`D�6�Jm�>�-[fp�$��`ʔɭjwn�0q����%���t,Y�eeem*i��V4���`2�[=�i��JHH@�v���b� 6�a����m��3�L8hP��6[B�4����h�a�Á�i�@����.��y�73���}��r�*���>}z�)�F��h���<X��o��xڼ�A�!11��n�SRS`���	H?����%���xU��HE�{ȥ������
@iY6n�h��]�tA�~�Z�w��}���m�6��o�1z����j�����$''#�Kv۷c���tٶ2��j��w�^mi�v�a����ѭ[ז��`;m팚��{��Q�����Ў��� �d�\ߴiS�o^�2�W�ۯ1..��fXD���F��@��r�4MCL��4�i��RXX��;w�߳WO����l����ܾF���cZ;w�j�V���;����iƗ۸��fn��N��:m�v:��m�-�)���X8���(_��~õ%/�e���f�w�.��c��{�n0��ٻg/���߆���vdfd�9��X���ۤ@��TbVJi!�H��J)$��#T�����6�5�G�����W��Ē����؃�̽�d�`2Yj'f���҉��m�F|\<�����q8���9 �)�@�MHH8��c�=D3V������m[�3���Lطw��vA�� JKK���ڪPR\��6m�j�"9%�]�n6��B��v�8m��T�w��)�.���Lf�����t�x��hTPPgee��Lf3����Ih�tɂ�b����$
~���-�;b�i�bs����j|��������l�Z�'���<��~ط��MK�^�O<�8fϞ��-Q�݆�U�ۍ�¶t����G����6��A%f���n ''6�.��N���p:�H	��pQVVVݩ��~
L��z ����d[Uմ)C�u������j6[`1�@��:%��c2���RZ��mP <^o�APD�(5M����P\ܶAZ4�`��5��2�B���9�+ ddd">DUdQQ
�x'-�n�a�f2��#�Q݋�)A��m�Ř�&�ڱ�Б�d2�|�^�V^OscL ����+8]U����J)��C7k��nGm��f�~�m� ������xRTT���o�]�K�1w�*@����]v����9�`>��M碦��E�p�iLGؘ
���>x=��E�"At�vxl�:i��;�q��;���O߾�FGZ�fmTݙn����+QT\]��(Tk���_�W����Y��Pe{�T�����zЎ���@�����G��e�h~������.���?�Ƞ���ʕ+�t���=�����SO>�?���r1l�0�9@NN`2��f����_�QYQ����r��	>8��4�cbjg�"j��M���x���;�<s�O6�f2�K�.�%:�����r��G:��� �>qqq�(����+�}�h���ښ�����_�k�v�ڵ�|���t��@��}0b��u֙8jԨ&�)���i@��������"�t�������QS�z���1��!+���s_������f�s�7� $�znC���#'�+֭]��]Î۱h�t X�~=���P����ʅ���}[�[���郣F�j�ل��m6Tx=h�Ș�������������mSi�Z?8P=�Պ�x�N�U.bc�پ��&�D-��U�!���`����wW�������rE�u֯��n�w().F「�1�2220|����OMI5|F���b���}�m;vT�����l6dtj��̨c3��HO7��N���E����$�/��f[:n@ v��'MBl\��f�-X�e˗G,�
��m��駟AĨ3�`��a�ݫW�w�;�W�����P�t���ׇ���A׃����S�N=/��g�n�6S���;w�t2�ZLucu,��ƌ9
��r��$�iؽk7��{��ko��9֭]���M�7[l�x�)HLH�SSS��c<�Hޖ-(*j�`F�Ôb��͆�$%%��8�D�޽z�f��������o���\�լ1��҉�&��Ն�1�_��.]0i�$(ͨ׫�?��.\tȿ�
���7�xOU]���G�8���1!!}g�Rؽk76���v۶m���[`ti�ѣRSSbNRGҳW/���� ��%%%��}�Y_޶mX�b�nۆ��b������ܩMj&
���a�4�}�L������ְs�v<��c؟�Ⱦ�
�����9/b�0�7�0u�T���ǰm�j6c��Q�XlA�TTT�/�����m��W_c�޽~:j>b���ٶH�{�n�e8߹���k�j��v�n�Tŷ�z�N��3N�g���/�7��x��G�漷QTT��N-"�hh�U�w�*w0h�@�y֙P���_|�^xa\n�!�2~��Wx��W��U������9g�k3�{�1�32��E�W_}��۶��) �������/t�}���aԨ����$
� HMI��1c�&X�����7o�m�/���|�}{�`������x��yx��'q��7�GCE���!Ҵc�:v��b"�Й���z���O���SO>��^zn���u���q���`�>��- e�̙ga��ͮ�o�>}�h�w5l\���|�8� ���ϰl�2�}���aÆ�ܤ�Ƥi8�	HI1�Y�g�~�%K����X��t����7
���!��W`KcƎAff��L&4��XE�9�zˉ&�t�:�s�u�(�_����fw x9�������栢��u��E���K/��=�����/���)^@B\�O�{L�q�=�*<������e����Vᩧ�Fee��{�2aڴi���>�/pth�5
�F�B���a�x��Ǳw��6������W_ᓏ?6\2>!	'Nl�6�H��Ï��5d��i�pJ�S �Ʉ�.��N��C��� ?���|˭؜��n]m�n���G��O�`ѯ��X� 6.��_0hР���ĉ'W_��ض5�� �mk�>) ���C=�իV!xէ��ݻaƌ�T��UM��y�Gl�:�}��'x�٨t�~������u������� F�Q����C�{q$�ڬ0�-���'����9�L��@zj*n����ۯ?�= �P^V���'.��b�2�5�;�ߪ�^���<�}�?p�����K~�6�L8��p޹���, ���p饗��Y澜?7�p#6l�ܪ���k��r�mx��wO0�ɂ/�C�a��iӦ�㏇ѹ��z�ܳ����BQ+{�+z��q�X��Q�UABb2.��rtJK��{�#6[�!x<-Z���΁-��7�_¶�z�����u'2�d�8�+躎_�	�^s-.�݅x~΋X�n=���-�����+1��q��s��#�"����8�N��[n����P�8�t̘1��}]��>�5�_/X �����Ѷj������E���ÿ_��M����
Ǝ�+.�V���$ux�SZ���/��2�.+����ч�M7݌�k�A�0�58�u]���~ß��>��Ð���S&c�ē#�-�L\|b�1�
�}�̛7e�+~]���g���>_�8?3�M)�}��pV:q�m�#��>�zd��t⛯��?���ݻ㨣�°�Cѯ_dee������NTVVb��}X�b%�/[��K�b��mգ�5׏Q0v�8<���գG��� HIN7ހ�k�b�eA�MAD��W_a��u8��p�93�۷/����҉-y[�чa�k�a떼�u5��[�����н{�QZ�șp≸��k0��Y�r9���T��rᕗ_������/�ӦMC�n]g0\���
y[����c�ܹؼqS��<t����IhR������aÆ`�*�ٳ��z����0` ���PU�B~~�?����Zx�_C 1�|�fo6}>�9��!��_|�Ep{<���b��=]j���x�i�zlڸo�a���@bR�6t�\.8�NT�������P�a��`�1������#Z}����1�Y����my0z�g��]x��G��o`���}�hdee!55&MCaQ��ۇ�K�b���عc'�~o�}ё��	����4q�8�ԁ	 �ł���
�v��K/�T�hӠ.��5�W��nǜ9s0|�p�1�3����Ʉ��r�ܹ+W��o�-�֭���y�|�;�#G�0�Y��=z��g�T���G���>� Ji���ǟp".���%%u�<�����}3j�\���
t��	��+VT�*�_l]�QQQ���2��j*��i�-VL;�T�{�=<p`���S�L���p�-�`[�u���;�g�N|�駰X,�X-PJ�������DGVv�����.�I��e��N �$%���^��z�MA�^/�lڈ-�6��wޅ�j��b�����v�ü��93w�uN�1#�W&ҙq��l;v,�5>�a�� O[ri��(,,DrRR�w#z����yUs����eO� j��̳��+�����<�����	��^��=	w������sϴ[0 M�0s�Y�={6F��y>�h�u.��ge%*+*��x�*ԅ-��!C��SO��/�����ړ �����܇��+���{\s><n*+*QYQ��*Wu�i�|��={��G��W\���!��I�N��aC�5 
�����H'?�h��;����Ç���O>�����b�"p��|\�q�2�T���+���;�����[Ӕ©S���W_��.��	�a�W��*���HLJ�e�_��_g�y&,&Z��[�P�+�j:��}�]x��'0t�(MC�`��@5�K�|���<�T�y�E��y��ͭ;އ��.L�s󭷠KvW�$�WTT`ǎ�ޅhn:zs@��4�����)���{������5kQ\T���Z�խ���̒�����1c������ɓjs9XGH <�<3�'O�+���E�����%ψ��GRr
�=�X\tх�4i��ڶ�n<�t�i��� ����4���vj�_�01�N��K]�������X�����¬�z��rI��o�V@lL.��b�;��}|��6o����=?Z�y��5�����_r1.��|dt�Ԧ�]D�=��ů��~=	<�l{��ߪ���f̀���+W���>_+ۨ�ra˖�����ݙux]g@oV�i�='���:\x��X�r%���{���ö��P\T��e0�w0
���I�ջƍ;�L:�F�DjJ2���
s�p��c�ē��w���>ǢE�k�.8t�N�̈��C�^�0��q�2e
�9f<��{���S
�9�2tX�1�u���ܾ0�ZYj����l2��HW�_G��}`j�H_�@�G��1x�Ph����޽{u	�y�6|x�s]ב��[��v���:lx��뺎~���j��b��(���9��_�ѫWO�Z]�S�f@n.f��\x���������`��U(�/���Fs%Jbbc��)Ç����N�	'��ݻäT����d6UUU. "���T8z�V||���Ғ��/8b㐐�ت�6�L�y֙0` ޚ����%��塬��6�( J�`�48bc�������sЩ:�2��w�ݳ;+��_r)^x�y�m6��@M��"(,,Į]��c�l޼�7oF~~>�N'\�@�v��M�`�ِ��Դ4dgg#77����ӻR��`�>�#u,j����Ǝ;�n�:�^�[�n���P^V��
����@\\,233�77���b�����̄�:��~�ʊ
8�Π�[,$&%Ak�ޝ��p��o�j�"!!�p���G���vv����\�W�t���"�{f�III��p�Dee%*&1�-HJJl�픗���r}/��I+_�Q����Rlٲ�ׯ�ڵ�k׮�w��n���!6.q��HLLD�޽1`�@���=�wG|\��;߫�n����=�4�II�߱���xQVVt\�a����M!P�p�@>��m�Ν�p����N@)���!11	����YY����n{}D�_�7<�ԓh�&4&&f����ڳo���P���]��^z1v;z+��]A���x<�z��z���|��|Д����
{LlVk��F��g���������J�l6�b�"�no�6~����/w{m�p����hَ�6u ^�.�^�70��R�X,�Z��Z�������<8X�>(��ߏd-�fa�! ��o�4���p���~���9�4>#�&���b�u����3�Ѳ�m* V�VKBȠ}0��<8�ېF?��z���ЯlCoo��k?�N^�)ԑ�|?��kᡦ��|	��:Q4-�����p�""��$ 4�ërg	���(J�Hӧ2�E9	���e�8""�(&�.͏3�6t""�������Q4-�����:�E�:�5_B�u�����(-�)�D�˝���;���0¿�h�DDD�>�.��V��0�E%DCm�::QTif��z2�E-�$�6tv�#""�Zv/wщ���VJ��DDDQIDD����Љ����ha������(���;#:Q4����3�E)��{�����(j�7�+{�E��&g�s�DDD�K­rg	���(��`�5��E��̶�Q0"��Љ��� ����ֈ���Z�Я�U���;Q��yl��`�XNDD�D��|l���(���Y�NDD�D���NDDtؓ�Oe('""�ja��V�E�0��Y�NDD���ǡ_����[���8�+Q���H�����Ba�;��#�8Rё ���,�E�p��YB'""�b��rg	����c,�j-X�����Vؽ�Չ���V���Y�NDD�X�NDDt`Fu""��ő∈���2s""�(��ʝ����NqDDD�?ζFDDt�p,w""�#B�m��DDD�,��eX�NDD�Z0�E+�GDDt��ќ��(J���;�Љ���Xx%t�r""��֒��։���T�c�3�E%�!"":"�߆.�r'""�V�V�3�E��*�棵��E��c��Z�)�����Yx%t�C'""�R�oF��Z5�ADDD�R-��>s8K�u���()-�����C�D:J!���h]ס (��4�]���������*�]�+@s�	���jE������U�HD�Q�y����>x<(M�b��d6!PFm�밴�����ػ{ws�U���J ��W�1J�DDD�C!�[�* W�߆v�'""�B���Eo""�Ù���G:%DDD�j���tJ�����t@y5�ie�N	�� ���v��H�����ZGӴ����2-%%�q�Ų������#�aK)����φ��F@Ff�q���wy<�" ���j�U�{N�p0:�%@��iͶ�����pD�g?��������9ETM)��R�V��}gm\�a�:����F�~�w��ի��2"V f��b���1&�ɪ�4��4��4�R�T��`B৪��R5WE�T��k�U�f�.�PX�v����RhxW����x9.����R�<\(T�]�R��ԀR����u�V���o5�k���^�=�:Z���Y�~Ԧ���������j��d}J��u�������4��Z��p�	��ʂޠ��^��u��c�o�5��b�x��/=��WD�H�����9��:{�~���������nHBi�{ͪ��R�4����k?���F��w���'��f�!��`geI��5�|M^�~�������4�	��t�cP��V�p��Vw\��n�f�'�z}���`����~i�'|�P������e��e��FK׻�68�W� ۯ9$���dݵ��p����u?t����������K�Y_��]�j�GR/���\�dX �5ikt\��*e�R�p��I�ɋz���ͯ?��ڹ};�~x�W��]��E��O�����FGT},�4��o
 �t]����߯ ݯ+]~�_��D �_W��t%"�~��s��oP՗]��^W�i� ՜ "�7H"XMŊ��>���]���>k��כ����}{��m�9��g���_y�7���4������]�78�J)���x���q�I'��^O���_��5oIݽj��O ��V��b��Ҡ���"5�RR�����R��$5W��;_���U_���BW_]�҅�r��ȁ?���M��r��7�R����d����/U�=}��Li��i
J��MдڿiJA�(/nKE�c}+M� Д��Ai�mk�Mi  ���;�ݨ�j�,��Q{JNIE~�<�쫇q1� ��)[�fʼ^�}>8u14��4��~�AY4(� ~?4ѠC�I5z�_�h�P ���\����k�R
���5��=�j���5�^[k�ª��5�)S��/uWߠ�cG��ɧLz������-���+��s�|6��0٘PRZ��n�/��r�������#F�87--}魷��ߏ�1���d�l����&��-W�ƥd�hT�Qu�T����7��n+�ꭣ�i�h=5�u ́�Oլ\I��������R��ڂQuU��K����[����_�D�N�	�ʹ�p`E���Hmy]�4����P��nOS
�i]��L�u@��lF �X`����*������t�	�v#..J)j|����Kv6X/�y	&�����D|B��v�G�7p9�� Æ��m;v���."�Ꟈ�����?"1�Xi����*���?�㳟�[��E�05�ک���L8�$�������M�Pغu֮] Hk�a꣏?�?���`��������'���Y看��6�sύtr����w��w��[o뒙���a���Lr�=�8"J�""�,\$	tMh��q�ۏ=q¸�YY�>,DD�XB��23�0c�i11��A?.\��Ҳút� l۱w�u֬^��_	������~�o����[o�S�<�$ŀNA���`��1n�ñ�d2]f͚�ض}[���j
@IY|�!|��Wh�p�RSS�>��c^�~��k�N\w�5�N6Q����[t꜉�cƞc�����ݭ�ye��ڎq������#�=.��xi��O�ظ���=�8�#.҇���Y,�SP����٫���7[,֢`�x�.��˯p{�	�>��3<��cpV��q��d6{323������7�Ήtr��Bb@���:�����:u�e�Z����l�2���V��
��U�qｳ�o�n4�(�����G5�I���6nğ��C��MDD�:�>����k猬7��t����N���?6��""���Η���ILL���#G���8"}���ڮ� ��={�]��A���d�'��}��*�G�w��l1A��M&�;;��"���.�sϽ�>DDaa�;��q���d6W[���b��%�r��j�O?��>�,�n����aC_7�Xٳg���H'��(,�d���>Đ��Щs�-��Ш}���8����T�n~߬�p`�^;��11�srr������G�?yB��MDD�>f�s..�������_�UQJRR���oDm���ȁ����f��٭[ϫ����/��F�����EXB��F�����,��>0�}c
%%%X�|y��j�������G|�}�)$%'�w������S&cǎ���D:�DDD�G����?`Ѝ&�E^�����rE])]D��>�N�A�i4��KX5���t���&"":8���[d�tØqGO���F}��a�u���	���`�|�J>r�a0�X�e}r�] ��}���NpDDt�:u��8�̳�&$&m1z=)9U��u������!�͕f����go����s��_o�!�YMD�jlC�f%�$#77woLL���K(���bٲe�Njuj �׋�_��?�F���0��~�j���x��"�t""���G���={?��I����9�|�p:#^Jy��s�vs��Q0hȰ �~c,X�l&"":�j:�6��f��g�"[�n�h@�����#Gs��������w?��r���]wϊt|_|���O�p��Wh�<zbb������v��ϛ����u�ge�?�x�4qR������й�Kq�Eg''��
�5Q�$�=�`Ăys���8�v�=�x(3���"�Ý9�	��CRb"����6
���˖.���D�ÁC*?��x���vW!�8�f�ٓ�����E��p�ݳP�*�R���DD�c/w
Kf�,\q٥����U�f|ڬ]���8�iS V�]������A�`��BrJ��G;��S�L����x��q.E�� �KF�;�j����GOLJ���y���ED
���/(�v󸸄���3<�s& ��>�t�z_|�N�p��:}P|B��P��<��#�$���x�^y��G�k�nn������� j6Q#�#��),�'O�裎����8�-'�K�.���:$����xꩧQ�D��vMӐ����i�Ϙw���`���8��#��DDD�ܜ� "Z�^}�`f�a������^3N���e���>o�IbRʢ�&��k��!����,$":hXB����J���V��f=�R
�v�Ė͛Z:4 %eex��G��/���4���]�u���W_nY�|n��o��B""���>j,N�xʉ�ظ�6kM3�#�=~�J�^�_�|z�8b���M&��[���������\�;�~O������s����GϞ���o����묬L��^ݎB��ޮϣ+ �}�=�x�	8+��txD��Qc�z殿�����>�L�����(z<�������]�u��xxUȰ�#dێ�ZJ�ۺUN8�$�vsh��m��㏱�c  o��v�����(��߸ 0pА�4�,Fϣ����7�k��."RVQ!�\�g1ޮ&��շ_������{���#�eDD�;�Q��ر		IHNN^n�Z���R(--��+�m�~��ƛ�׿^����oUӐ�)��S&M�{�Y3e�M����t�E��3N�̳�����ۨS ��K�UU��R���?�$��䆬jOLJYq�)����,"":�XB���������p�n�ܚ�kPPXئm) ;w��}�fa�0|D�n/�޽�_9͇}�����HgQt{� "澹�_2`FIZz'��ZUB�W��t����ILf�a�\3Y�n�{>�ҫsmW��Z<=��HgQ��UU �3�:�ŦZ��*��}��U�~y��Krr�W�k�����3g��3���0y�4�qNDD����
#G�i�Θ�P���+/UO�K�""�M�����=c�>�d �DDD-u�5��ڿ\ףS�����Qc�ɞ���.�׌Ӿg�>�q�!K��͓�o�-"��v�x���"�-DD�Nq�*��;��O��!�U۾}�n��z�*��>�>����S
��>�0�9g�9S߱s'�v�u��""���[�[3���&�%T)Z��R����󎤥wY:OLJ�8q�Q�9�  �/�t�~D=z���i��pĹC{՟�������V����G�l7����G��= |2�K����HgQ�qrj�-[�`��G#..n���(v:+;U��^���%蜞f8Q��_X��+�-�Qk��i�ҥ�[����7F��5�V�9-*Q�=��l�~{���[��qY]rdђ%!����̺���cBV�wꜱ����;�����@���������7ބ��G�>�ߡ&j��b���n�ED>������jW���P|܉���7��>�t����{ ��S��d�;ĸ]�u��M�>_�`�f�:9j̸����M<t�c?.��z�?f��g8�9Q��vƙ��UW����^���ēN�����t�������J偗R&�ֽ���xc��睏��^�]'"":r�����Y���G��ޣ׶P=�kwY�|E�������ǟ�G\�vs%)�i�Κy�$ p�uk�ϵQ��v~[�,��1�~0�r��~�?�Ou����_~%9]���jWb���{�	w��魷����|�]&"":򔔕AD���N�b��hG�t��]���{ٴe�{�	!{�k&�<􋧞y���7܈y$һKDDtd��変�\i��xC��%3N?CV�['��j1�X6;���k�������W����G��Y����}��l��\@��8d����h��<!1�s����$"�_~����#��DDDG�5k� �Sgddgǚ��OB�������Ymr�	'~4��S�}�y�:�_��M""�#ߥ� ���z�����u�׀���=����:�\ �眈��8q�46�;>#>!��s%�]���DD��nl޶-һGDD�q|�� ���g���[��f�L�>��=���~��7X�zu�w����c���7��~������̬�ו2�8��cbw�vƙ�fv���v""�����G{܈ظ��-
�J�9b���õ֦�:>�/һBDD�1=?w.�="��=z]g2[��	��"i靾0hp����b��a��""��������N8��8-)!1�悹R&;n�޻��Ǥc�;"ªv""�H[�`  ����{7[�뫫ԃt�-��w]|��h�N'�{��H���o��S�L �쎋�L%]w8�^�<uZ����GT:��N:���@$%�"%5�j����i�FU��j?5�Sv�,t��k6l�t�����1�dA�Ι8pprFf������Ė����LIM�ӳOߞv� p��wG:�DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDG���Nþ�C   xeXIfMM *                  J       R(       �i       Z       �      �    �      o�           ����   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��    IEND�B`�PK
     mdZ�����  �  /   images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.png�PNG

   IHDR   d   d   p�T   	pHYs  %  %IR$�   xeXIfII*            (           J       R   i�    Z       %     %      �    o  �           a���  �zTXtRaw profile type icc  x��S[n�0��)z^�8~$R��b;^eW�J�ё"�@`H�n-|DI�D��@ȴ�v=L�"�	�s,`�ۮ��z����"H����pz����3�ͬ,9&�h'�tN9#���(���d>CQ�h�|q�k��R�R����mOi�q�6�Z�ܶ=���C�>hrK$>���U`�͚t3�s;����%�S�T�c��\���~�y§b�_"%�G"a=}J�H����|)�Ni����2��yl�c���r�E��|�7$��8��s���.PJ����
��wq�8��P'��j����[ܞ�c2����g�+��|����RM�=�c2gҥl��ϞauTh���҈�\�z���줡㜥   %tEXtdate:create 2020-01-31T21:31:09+00:00��y{   %tEXtdate:modify 2020-01-31T21:31:00+00:00	�   tEXtexif:ExifOffset 90Y�ޛ   tEXtexif:PixelXDimension 1391c�   tEXtexif:PixelYDimension 800�요   (tEXticc:copyright Copyright Apple Inc., 2017���   tEXticc:description Display P3�y��  cIDATx��]	xLW~��d�(%�J"��}�%(�Z���B��_[y~R�R[u�E[[����J����ҿZ��j��B)��'s��;��Ĉ����>���=��s�s��-�37:�PTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��AW÷&��z\I���7�)I*�Ev�Z�:d;iJ�3mtRɲ�������V�$IY6��"a[�d��$}/����~�l���99��t.��$u0Z��d�M��(��5D��a�}0�*�
��?���h��dY~�`ȫq+��L��yY���@���[���������ƍ����0��`�Aк�C��"�|<B&�������r����t�PQ:�;w'N�{˧����a)y���3�t>���ʂ
E@fB\yyP� �f�3b�1�(p�3!�<ÃY=��䫄(�d���?0��&1A3vH�JIi�	�YCd��c,�p?��0���g�Ж���lqtws���%b�G��ɒ�2d'jaxR�v�Zl߈s��S�����_C���2Js;�i���8�f�ɒM>�Q.]�����С�x�g/�5J<����зO̚=�g����f6.:6lX�t]������B��5�D��;ѽ[7���s�p�0g�,�n�=_x��(���E��~/���u{���F�m�6�2�h��!����v����;����dX�i5�7�}�����ٿ�2~޳?��#n������1p�@xV�$��u˖�Ѳe��H�zi��|��u��,�Ν'�����ԩ3�/�5PP��7o���,�_���C�޽ѵK���ǚ5k�t�:>�,^|q 4�XȺ����7!&&�+{�_�~��d��ǎ	SԥkW�o؀������A��n��B�p2�7n����Na��>$3��ARLN�G��&����~�� �����QQ��wq�������Тe+xU�ºu_ lQ������͐�լ�K�.����ԙK�.��9����(�QN4|���X�p&M|�����5�OLLDu��x�"�.Y�9o��&�l7ww7�b�rD�c�)��?��޽E��jO����[���a�0�?B��ۿr6n����o�Y�}��E�E�:uh@lAZZ*�i`5]�ر�u�9Ǻ��<s�4�V���ի۽��1�Q�n�:AƢ����D�?O�F�g:b����a� i4puuÑ�#������W��u� ̜�iL8^<H�Ȏ��ʕ+Bui������®�v�u�zS����u>l�ФΝ�P�U�@.��+��������^M�5c�L�L��S��nW",�Y��e��'""#�|���'B�B�FMТœ8���	�R��ӓC��w��t�b�_G�R׿ƛG߭~=L�6U��?���קў��ݻ[��Z���\�rLd0�q�	��o@Ey.D<kI��
2^U��~�zB�!C^65V�E�6m�W���$!-^�j� ��溃��������͂�٤������m׮j׮����{��l"��e����G�fg�AQ�%{ΫbM�6��F�흚6m"�.\@�ƍD���]P��	��g�ΕG���e?h�V��\��ӊ�����ٳq"m���`1i.�[8c:fd��Y����<P��6���׻�2�sq�{dDG2kd'j	h�͛��)2;U�jW��%�=z|j���)�b~b����!JcӁ�L��+$3�i��ߪ[�Fc�8����2�F����~~���dG��?��%\�9���ɡ���3lw[wGDD���Ç�6�V�Z8AQ?��6U_"���YԢq�0��$��_M�i������W[P��@�nns+�F*Z��@'����!����ǤI��`�<a�CI�>��p������<*T�[�Cɩ�1K�,>�>}�/�h�M�vhD�*��89�-�aq�֭�M0m�t�jQt������5k?C��M�ۻ�Mk5���Z�e����ZSVY'�����L���������'����F����g(4�Ŷ��P�^G�>|<(��p������_�R�VUDK</`9rr��WhI�6��E^��9��~��΁�ʧ(��K�c��K�^���}Ѭis<���b�s���J�efp �e
���,���5��<�5o۶oD��h���%.�sab��F��%a�ȑ4I܍��u�Ȗ-�!00�==̤?�9@���������A��"���K�T����J��2
�������r�̋h���C�Шn+���\�t	�i~`�'t�dA�����Ӄ|�'���GEDCQ��z�5{zP�gA`�@��?�h����\�h*��5���]�r^^^pbb(��1��[ޒbo�ػ^8�s4�叽|�4�@����4}�#0(h�my
?A�#����Mg�<��7��?�il���_ �2Eto�����"����j�37-N^��4g��)�8����&��'�*JBCLQ�JH�C���=d��,���}X5D�2`�����0��g窆(&Q#,���!�.o���e�TF��[���9ʲIQ�[�<l�M�V��|/="D�xOR���vG�_G�3˚��7��aj�gE��s�6��ˋk�Q'I����܊�GBEiB���j���QCG�h4Z�D�$ݢY�-R��By%�V+i�T���I|3����4����ĉؙ}���2r����)���Om�fk\]�zH�|�R�iO�l�Mۗ�I6_dْϜf4G��Fk-匷�ݥe�k�\𛍶���V���_�3���X:�-�b(ڴ#ݾ���KĤ����h$�v!VI~}��+s�^����xg��p�h4"�E@�Ӈ$^N������1���	�����ǁ=j��������o��qbZW�?��i�1��wI�t�G��v��e��^3�x޹���k+�t�w��`-;q<3��rJ�r�##���Κr$55G��޶;�a�±c_�ٿΜ�V�{J9�Ԕd��=�(B���}�\�.1�7����׭w�^v�.\�[��"{x<����̣������{�"o���]�|ҵ�"#��[v��n�ٻoޚ>�Mۢ�̛;[�A���(Ks�#�����@�V�s��I������׸��������gn�fV��8\��@�*e	%F��#�n�����8v� �2�Ǎƙ3�2+yV{<6���ܜ����#d9�¡��ȏ ""�z�ז-_�M���^nzjJ�QNk��i�܇��#��~_�Z(_��?���&��2�G9��ɡ�=�gge|�yx�fY$�Q�/R~�'������ll���<����� ~�N�z�����t
s�PVQ��<^�q�s��mOrrJ@�=�t-���K		粲24x6�;�;�%JHJJ
*�|D��-KKMN!p5�olI�x��ݺ�Ge�F��kǏ�H�"A�ռ!i\�xzz�/_�<�R�u�7�u�����U�F��K0��N�rx����̬L�(B���^b���x:y9��}���E������k��%u����QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB��A%DaP	QTB����Blg���    IEND�B`�PK
     mdZ�L+.�N �N /   images/7139d0cb-a6f6-4338-81e1-1177b1f79563.png�PNG

   IHDR  �  �   ����   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x='adobe:ns:meta/'>
        <rdf:RDF xmlns:rdf='http://www.w3.org/1999/02/22-rdf-syntax-ns#'>

        <rdf:Description rdf:about=''
        xmlns:dc='http://purl.org/dc/elements/1.1/'>
        <dc:title>
        <rdf:Alt>
        <rdf:li xml:lang='x-default'>Untitled design - 1</rdf:li>
        </rdf:Alt>
        </dc:title>
        </rdf:Description>

        <rdf:Description rdf:about=''
        xmlns:Attrib='http://ns.attribution.com/ads/1.0/'>
        <Attrib:Ads>
        <rdf:Seq>
        <rdf:li rdf:parseType='Resource'>
        <Attrib:Created>2024-06-09</Attrib:Created>
        <Attrib:ExtId>a83a9794-4a4d-4c22-8a84-66c76feccbc8</Attrib:ExtId>
        <Attrib:FbId>525265914179580</Attrib:FbId>
        <Attrib:TouchType>2</Attrib:TouchType>
        </rdf:li>
        </rdf:Seq>
        </Attrib:Ads>
        </rdf:Description>

        <rdf:Description rdf:about=''
        xmlns:pdf='http://ns.adobe.com/pdf/1.3/'>
        <pdf:Author>Firman Abdillah</pdf:Author>
        </rdf:Description>

        <rdf:Description rdf:about=''
        xmlns:xmp='http://ns.adobe.com/xap/1.0/'>
        <xmp:CreatorTool>Canva (Renderer)</xmp:CreatorTool>
        </rdf:Description>
        
        </rdf:RDF>
        </x:xmpmeta>!��  ��IDATx����l�q'�U�޾��p� R !��D��h�#E����Y!�'����_�p������!j�9���DInC��vqq�o��,UεNuHJc��)�o�}�:YY�����*ahC�І6��mhC�І��l �І6��mhC�І6��h �І6��mhC�І6��}D� �6��mhC�І6���#�@8��mhC�І6��mh�6 ¡mhC�І6��mhC���mhC�І6��mhC�G��phC�І6��mhC��>�m �C�І6��mhC�І�m �І6��mhC�І6��h �І6��mhC�І6��}D� �6��mhC�І6���#�@8��mhC�І6��mh�6 ¡mhC�І6��mhC���mhC�І6��mhC�G��phC�І6��mhC��>�m �C�І6���#i1ƵϷ񵭯Ӛs�&�U��)F��W�W��������J�W���tL�p=A"�+�w��n�VZ��k|��W��|!#��ͮ�1��w�>Q��V�
Gt+�f >�4{p7�c�f����;���g�����=��#0�ʟk����z��Z����[>��t#����N�']��i�N�W�W���\_� ����5���;ft�qAzŶ&���5�~���&���7x�/���ޙ�,"9�c��DG�����0�^%"u|�l�ɣ�"���vc���>�;7(����h�Ƒ�C|��!$[�����w�E�/\ o��&���͛��L�����߼�&+��uQ8L&PL�$
���b�Q��U��x]�82Vq�ߏ��ϋI���s�Da2���s8����\X�&߄������Y!�^���~_[�u�30���DCYw��������=������U�^����@D���S�N|�Q
{W�w�#����_��1���2���p��ULJ�uc��x<f���F:�X��&��8�2������!�#
]��1�N���D�s.��^����%=�+�V%���1�_���s����!fAJ�;�Nb���e�t#ږD������BDƈ\W�u%�~��x��0O�2.H�Ȋ���^��8�kN�<���􌥎��L��)�fc��Sƹ�3���{R��v��iFL��m�U9C��8�Ç���������j�M����mM׺��`�5��wh���_���"�9K<��6ȫ0������b.�*d>x1��K��~�VE�h�F1w��xF���.n�*��/O$C�s�G`�4+}L4"	�xd仭Q�b$�&��$sb��p<�/���Bנ�n�Ȝ���a��H��w��Ώ�b9w���w<���Ǿ�~���#���H�I��i
-^1�s�_����\���sE�&�ۋ8��r�����ӄI�s��Qۓ2��2�Z�8�� �o-^��hC������`�u�H�*�4&~'�uĳas�[����Q1N�yz@��hX�`C�C:7oV�co��uo�Xw����|K�xL�u�n[���t�Gz��t숖�5�\Lʎ�=�'f�����iλ��H��&.�Ē����H'F���+��v�����s�G	���[��R���l�}L�O.+����,^��=�.^�'���P���p�T>@�N�V.ΊYc�8�g�7�Wu!�>��|�D�Z�η(�Z�[�E<�w!�ߑ��ֱ��	�dP�]dZ��"�I,�RU������v�e��D�M�5uJ9n#����c�@��ڪ,k�[��G}C>��W��,Eg�,�O�q��tׂy��5�L���(+���n8oH�Ƒ/��e�s��}���^ď-N'��At(�ǐΑ?�$p]l�i��4^�_�v�g�:27N�E�t;~��NJS��tMWU���3]W���9���{Ǆ��<���y�c��^pi5-���|e3Uu`����3�G@;!��.�(Eh���8�ɽ��&?�\�(����C�q4G۶&��H��99F�yy��m�D�cث��	CBz 7����q7v��R����n�fV��?��K���x��H�$ �y�W<��W��F9*h2j`�G�¦�-�d"�~
l�;�d���xK�����/��u�I�4�o�e���c�fx�B���d&~�q� 
�+d62���A%2�tN,Q��ќY��5Z'�|�D�����fS���ʳ�W���lV`{ﻅCТb5�P%��6/�k[�yWC3�ӱw�>�������p�������O�v+���^�}��y�r��O�V�@��t��"|���� ��(4�[�+G³�n�Ȭ�&���o�:��c�R���Y�V(���;~����_���(-
Q�t�3�-*Ӕ�S�_lܢ�F�M�&��C���;��zpD"S�.�-h%1(H�C5(�KXl:U~!fp��
8V=PN��ETⅿ�:fD�	W�{עjI�-*��CI��Ci��kI���(������� ��|ע�lZg��B��<0�<>w�);�HYGz>`�ER�{S,"���*�Yj�+�T�����_V�l8ɘ��*C� �;;�"�㿘�����_m�@k;U�dn�AD7����a:��\�5m 
�kj��N�����h��'��Y���b��?��s#�;��)��_��L;�u�jU���M�ё8�;V��`u���q�G5c��<�](�������h��<A$�����@�-�1�%NOd��;[��h��"���X�����A�n��:�޳��:u�C�����ғ�����t�2=�<^�3�9����\jڮ��U�c�F��O��7!Z� ���F�7�@}�A[!�
~�E2�\]�����_���x��T�S���=��q6�j��m�;F�X4Q;`��#2{z����L���3p����5O�wʅ����tH@�Ȯh�����.tN�>u�;1}:B_|#'�G�t̮���(Xh�!� ��J$$3HT���*����rR;��e� YP�`�Et脭y��Ņ�|Y,ձ��E��m����cy� ��w�_ԯ�;h�9Bö�4켆}��M��hc�ب7I��9���u�@vQ�P���x���z5#
��Ɵ�=2���1�� �	c`�	5��'O,�Y�D�m���=cӤϣ ���L�z�9!OD�L�AEMA�������V�����\T�#�,2����,>U5:���l�3uAB�B��|,�y��W�#��I����3�~��]Bs�& yQt�*3e��I���&d�ܮ-�B�웢�&�MΫ
�\5�������"�Q�3����������r����	w��쵈��x��=��2Π�!=�����S�LWQ=(�����s;�.�NL���l����}y$A�i,���7��.I��ϥk�g����TJ�o �P���P�dN�T�	�2��(G]\�Y2��N�^�h�wL�Y�V��ᚖtk��J:=���4 ��&jeF��N�,	s�:���m��ժ��fP~�T�Fn�_�������j��~3��q�����Q��mD�
#z����<Et7Q���C�ɤ��cng��펔*i�#�JI\���]T;_}�ۡ$Z��XP\�t:�m(X0�T�:�����0>���K�D8���ňC��L6�x�lbS,�CG��M�Ey3�1��"	Ӫ��;��t��=y��E6J��v��4��+2��#��'@��H�19"w3���%L�f٨������΋�%�!�"�ˁ�c�AR��'rh���B�����6������4�r��Sd+� ���q��(�Ѩ�B\!%Ve`�9�"��i�J�~�wx�D�ѳR8�|�j�qGʬ ��IZ?h��g����쇨�N�
#��ae�B�� �R��`�v���"x��2���� �W�P�I��8pI�F�Ύ%Z�%߂]�bp��
~�jL8{�1�t\�����7��q[�hj%;&ظ��}�p�!�n~�p�r��	����^iS�*�ɍ�Z����yg!�4nqF�b�9R��H�����>��ſ��dm�Ⓚ	�Sz.�&9ѽ<����W0�O�v+�D�$F�<1ru��T��9^��G�)ض�LH*(*M ��?
I=��2���E��y��6�M���1��`�7b.��tjy��K緝t��-yF�`��#l������(�;##!T5��䡴���L;(��0f��c[Jܔ !�� )r���&4�� �k�`�b(Z�E?{��A����[lO�Y,4�Q�Aǉn�i�4�J
2J�|����"�é���rǮeo7�xY�����n�iT]�xY2�"���z��S��s�X��Y�(QOPV��?�r!��ʢ3<E�͋D�(#l��,���x�`U�łJ$��/P�"��<~�19A��{|1��2�����oo�����c��B�2�^�	�ʪP����ayP��:��C�"�]��>��'����^\�م"��q��U S���$˦5IÃl���Q��4mV�bV;X�Xl�`�����J��&�QUY��3z8}V���ή�*�����.bۼӈC�KKQ�]T4�A��ι��J"�Yc&�W�X�F���	^T�@�C�Z��#hs�Y{¯�����e�s�r��e�!�ȓq�u,�1�^���i���/2 ��RJ���z�1'V�J�a��)�V�d>��E��$@�).*�9RQݩ��I�{ʽ=[��y�̚|ҿ�Yӷ;���2�������Iz�H��ߤ��j"��o�`��7���*D�A���d5/�^��b�l2%dIͫ�>F�	M���b�0��D�Y�RM�3��Q~��Cú�hc�Vq35kLXZ'��&�d��s۠ϗ�pq�����w�x��� V{%��cS�����kǮ[�?:j�\>���5η���t�XcS�^�Ɩ����RQ)�5�����#%�-�Eh$M�}|�	m�y��'�O��u�����𫮛��^QX-Z.����$��#!�"6���%����)<��hcQ� ,tE�F!��93�I�H(�'����j���u�Yl�mePEu+�Q\� ��U�Uśc�0��@6\�����7!/hE��Ml�:r�w2�vT /�� �)cB�Eva��t��@+J=�ˎ?Uا1+â&�ؠ�h|�(g!�%��B[� B�S �+�[J?|l���+@�&����kBGi�Y�1��ǵ�8��S<K����
�i�g�41W<� m4�����8E��
(T��@�E�8\W�d�m\[�z�A�J�:(�ߵbb���
 �n�=�қ%jc��x0e�Np1�jv�ĂsXDǉO���6��8$f3�;J�+F�Y������E"Kd`���6;�=A������zц;�z���^������;~�q��ZZ�2�I?��6q	^��h�cj�%h㊽�r�^jjC�&AA���D�Iߋ5���(�@��㉞o�3��F�\?�ʑ��V�d�-�(��w�}�0��>�"�靁�9ѝS!s���x1'����(��1�;�� }Hp��z�1K�б��Lʛ���Һ^�r��msU���OMcT��{2����F���}#���!-?}�FLL���4ݓB�?+7��a�)��4�Pv�|6?���k2;g�!9N���B�͠\�@��X�§WI�Q|��-|�$�co�	��Dc8��gך<碫����~���
�l�$>�k����q�,@��^P���`����]� N����K��p�:���r�A��K�G�fPq5.��ǚ���"�%��>�U�Tݚ�ۛ��}�keHZ u�Kg�����!�Pt�9qי['Y�}�T��b��N4Fzl6����"ʗ&���-~&����dgs�5��:7T�*QX��q6����g	)y"o�T��ɛS���Uߞ�D�F#�_�M-�p�y��Q���^��;G�μ������~^sY_6O�u�)?hK���c�s�>��c�^�_M|�)`����Z�$��ܡ�����*Y��6@o��~�O�7(��eZv ��>Sy	I�qw��k}������҃M@������ݍ��]/�����n=�xxQ�{���CTkw�}�pA���Z�;q�|�	��5Ȏ=o�"1��B�,Ib47��Q$�,@I�T��.9�{Qr��K`�rJ�sB���%l�5�M{�F�O=G�A}Қ��p�wb2���nY�gl�O�Z�žsO�V�Qm,UD�6`��,yvE2IB����hħHִ9�\Q��p��^�@!DJ!�V�j�t�oJI���v2Kͅ!N��(\M)1�/�Z�A�s�a7
�����&rP�q�$�$�YaR(_wf�G3l�S��x�j�Ā3%�V'՚��9Y�=�<��CR��P��|?';u�R$���\k�6\d���Z8��Ĭo���[�F�N��������2�=� h���yukt �~^��	O��ի�FNTP�lD(R<C��(-�!���à��q���k�1�or���s,B�<NQBg�Fg3e�L����,b"��h�P�BLB��֝����vh!�d�j��;S��/qK�)��f�h�]H��w"S�4�g�_��&c� "f�8�����<>��j�%��^�[G_q-$Ѫ��}�~QD��������+ѓB��(���iV:(q���@�@(��j~,]"�9P��% !}�̀��#�����
��aJ<�kNe����#>!�Kyi$7�3�r�:CS�0%ǂ�gr���"?;S���=��*���'���(�=�|߀@n��~�Ӫ���&8�j��Ypl�#��Ү�5+����睨pW�Rf����&$�I�LH#�]��I�e�S@�E�2�Ҩ�$��;Q���s��of�yu5���[�Tק5ێ�Ӭ.1��dJD6�M��SU���H�0��m�f�'�S���,1�"	�)Ţ�iņ^��e�jul'"�T�z�e��9uV(��O�q?�6�����y-l�?��rӔ�sM���9�K��lHR2��esfP�hz�������w�:��Wq]��N��2(а�����i7?D��=k摪Ӛ?�.I��}.d�|��{�)]0;a�B��u���ES����t��$�g%����۳(��Xg��yƋI��RDm]��2�	�klfs��Q{�@�X)�GwOg�wӑ?�ɢn�Q��G�Rz��0�Q�!(l`�:v���R�q��PS ��!=�u�s��r,���^��:�������>�Q��^M�36<�^��ɨ��z��X�x��Aن=Ӭ#u'�Ja����"��")&�X�1���e��0'g�}��4]��2]o$�|��el�c�
�<��f�q����f_��dlԂ,ʜ��ot���=��d*�2H:K�b�T�纊��Bǒ'<�1�z�}�T/z�6��!t�`�FW˯.c�#��	�.[&�)��[j�&��E��i29�"�#�*<K���ˏ�u�Z��hT�3e��7t��ms(��e�Q:�P))����<a:��P�Ͼ��1-��bDkx�եͭ KL@�1;�:�Ζ~��|��\�}����9�W�A��d`<{��K�7=����AoW=�3AJ���Qg�حk�Yqғe�j��2E�I��Ԯ�LΩ=�j��$�T�uz�39�ҕ����ǘ^�4o���ٌ��<�9�E�D�EN�5�:H���� �����9-	tq�BJ(�uT��R�Z��Ƒ3��J��I;"�[�bY�=�£[��l�&SؚN�}2�Pa�wU��)����%n����Z���tw�������`�@q\�d{
�l�������\�6�4E���h��S���5�ԺeaLi�L@.����Dr��)=YӃ$y�q$�G�ذٔ�'�(��3"�C�T�����s���0�+x��Exto�������.^�����C�cҢ��#@恍�*e��s�XTy�w�ƽA���x��bA'er�s����k�<���HQ�.(�r_K�Ս*��N�,j��d\��1UF�_�!Z�������L5R�,���W�e?���Z&.�����q��g1-� ���]��6݅���>��\�
d�R.�|�C���U���gYA�l���бs���\�H�)^�k^US(�=�౭	&�;���s:����9��B8����.�/<p^��s.�N��~?E��J����Y�횃I�Θ�����OmgEK���$��u�y���N�9I�x���F�M������jv.����F�\]����e�Z�!��k���lgV+'�K?�\��]�����\���ͼ��ȏ�A3j, ��̼@����eʢ��ּF���EU-�6BRh �h8�>��M!)4������
�_X�
#��c{238-��t+�]�l���:�N�x�Z�`�\Xj���
���g2�J��Ќ��)�7�̋�G~L�+j�d�4.�b��� 4�F�N.,�ѝ�ÊGj�%c+�0Li"  ��ɡ�|��9�t^Ei@��ܟBS���i.Fw3?��N=Yd�zaX�'6z Rz���Qe:6,C�r%tܴ�}�KF	��(�zŠ6�n��|zwRQ�B�a<�C�WkZ.��B�[3����p��>x:���/���1ją���¡��#��`ǋ6���xI�(=Gc�L�@��)2p��5�;L� �2�r��@r�X��@3ū���e�,]3����e����r��57כE�r�^���A"w��ڵN[Oѷ�� C[x��_~�t��>I�8R�ºf�ԫzM�1M�YT��+�L���1�mB)���@��%L�i���K�xk����U3IN�F��;;�d�W@T����*	���=���5�)e���������-Jح&p��ܺr�~�Mv`��t4�1��H#^�
�����N����  I@{���`5�,����wރw� ��p�������J�E	D�u8��N��J#�."��:1��J�0��ZEvZ�i�TښV6kX̗0�M8z�q�l}d�)p�@�����\N
�^w�l{�*"�j� �i�c0���j����O܀O߼�<S��
��r��F�|d����1�W��L���������Lʹ�ȕ�0���4�������j��EFqF��|Wn%Y�'m�� ^&濫J��V�ij<�^Q�K��i�*@!���~h��#�j8ҽ�I�`S�;7J6��$Y�'��+�Z�� k��;�}́nY%|���9��V�R ��u3x�
�5U.R׃,6P�c�&C����_�1j�Y��8�@�,��z_
�p�8��G�X�=iNd��P���swfe*P���^�m�R������X$���"�ϋg�]ܧǤo�W�u)�rp-Jwrk�#'����|���o�y٨k��W?�睜��K�K�����+��c��qfW��Y-O5ͣz�t/��O:U��
ˢH@4�/:�A� A�#�(*�.S������R�<���(Ҏ��wA�T��{rBR��)�Bӳ�cS���$�y���o���+y��>S�GY-�@!�4f�ٯv#�	*ڤN����0�Jqr¦��i��e^7��*�K��`�������%!���b	���]U�_��h!{��ҧM�k��cgO�ف,��N�C�OY��51N�����jĵ�غ_�M)��� �c�W�� p}��]9��,u�ue�L�+M����k���^�Uo��������̬xHX�Q���&���s`�o��uti�d=[�W��#z8�A_�z*�̆l���u�)�˃�gDR�Yǌ'��ȟ٭)�4O�\�<�'@�\S�Tp�`2�b�����	��s9Q�cARLe~��I�~���,:�"�^�������QjܨrT��֐�p��U10�R%���>�6p'��z�̣�- r���1���s�'d�@o~�i0J��uGH&RQ>�%����{d��=�#��N��s-�� �)g�@9�B𷃆��"�GK����,�Q���`��"Zʜ��|c"l�Cm�%�5R
���9��{S�'"��.�B�7�N�<�و��\�l�����ūpu�\����d����-�#2�J$R'�>R��	&�.� �� ���3*��h
׶��84	������EP�ν;A<\�a�\q��G.\�����h+�RD'���%E�KǞߒ��O�إ��~#pZ,j��b��Q���j�Es�h?g��Ak��/sP^"2�ɣ19[�)��5�g�p�����L��p�hᅫ7�zx��}�u���@(��H�y��rd�e�@2ƴ���R�H?��<ց��֬ls�I��AJ�Ɯ	�
A�֪��<"�m1aFG(�A�8���(��h�tB��j�E.5/�F�v���I�~�S<��kӆ�lӢ|[i�����w���������n*B�pq�x��e$����WIIV�:U���`QE��l�c�}�}LF��-�`�"
ʜ{�F�r��AKRI��l����hQ1.�7�auJYd/�;]H�|S�<v�^\�N'����rZ7%}8����l6;NjsXjQ��A�[��������yG3 !Ϟ9�xq���Hi�\���O�?�
����;�|鍔�m�9� ҩ�H;׿
»Q��n��y�y�O�=�\�B�k��9�s^�uf�Tй��{@ˍp�;�}l ���9q��]�b�8SƁզ�O�C������t�imH��R�f�����t3-� }@�ޭ:�v������_H�C�V -��M41k]'��%���C2 ��dx٭�na�\1��,<\"
���e���B�Ѓ@���,�����E u��.F��C2V���*�}ZM��$�O�蟵(��yN��%e�Y�ERS�����-�����H��9�1�P��%�Ɛ%r]ud@1�K*�X����CIj��d8id f4(ś�Ɛf+	f�#���xC������:Y��q�
�4�	�S�@��� �{�}�'.���:{�Ұ�т��h�Ǿ��_��ڿD�Y���̐�C��DV]�i���F&��!��Z0 @�:s��X���w���5����N��ʍ��$��b��8�4�N�"��?R�Ai����)���9�l��ӝ}�YO��,B�Xܨe6��ĸq��麧��}d���Y�A<�[�����ާ�:}&Y\��Q8���I��`�a�'7�L����&��i�1���)N��<�q�:�C~������bd���'�UhASরB4#��u�^�C���Ĕ�&�3�f3hV5-x������^�ޅ��?�0�F0)G���,���N�cY��ڰShf�("��q���!����hVJ����mx��pD`����T6�&��Q.�;�-e������R�2��OD������W��~K4j��6r��%�����F�z��K2����5���2��Ob&اQ��{ua�6\u��[��w?�)؅ă{'%�;S4N��,VT�^�"t^��z��'���XS�@� ���ʛ���ֺ�����x�ʤ���y�J���4���{�N��d�_|JS勨/J��Q��,���I�tg0ym�C�Hv0?&�K����2����o	d��j��RT�C�`���#�(]ۍm'�մ�<f3���N��Du;X5�� ��D�#�ÅX����76�(��u��6(�q>Q:2�Q��d�D�����1�K�Ń�@Fr�I��iݬS��^ұe��M3�噃�/ͤ�؏铌��Mc)���tg�1s2�"��:�����v�ܙ�ikD��m:>/er-o��J���t蔖�S̞�e_���3����u�y64 �j�އSz������ Co_��(�do���+h��2�xgU�w��/��
���?�𾋨sKq"$�O���Wt�K!;O�5��G�B6��l�j=�����t�G��K���r���+m�t����z��4xI3g�dҲ�I��I^2ʩ��*o[�ܱ')J\�NX�䚁�KA�.-�Ak���q����A��Ժ�$1�D�u�y�:1��l�N`��%����3DX����2��كD��1J�RA����C��@��Ku�R�yQ����?�>#�����.��j)��d��^�բfe@^h���x��lk�����+T���1��O��d�pik/�XZ���T8�Z֍����9~�M"��Y��14LF*���W8	
�`�")�/�vCFP��Y2
ST1z�Ԙx���d|e�]r���S?7��	`��y�&5��>�����Y��%#"ym�d!�c&������Z%3�� QK��N<�u���$�7���6��JL/�W�vШ ���F�w����J�*�QL���X$�I9���^H����A�� �����My��>��6�چ%�s]�<�'G��%��,.%:�^�X�)*�T�U�jW5��9���EI��*ɠ@P^���-�u��7�����:�������8�F��U���H�H{�r)b��9�f)�f�A4E�8���T}���(��)}q{kF�+Q�(K(%sw�;�-��z>�e���R�"�N�?�r�{oT���J�e�küx��Q1�������ʮҩs�i��
Ǵ#q���̩��є#�xk���o�Y1�o�l�@�d��o|�6m}��7�� �Kt�梙+�N��lHzҷJN;+�a|�<��c�n�9��C��.�KϾ ���0:<��X�s����/�^_Z��xyn�·�`��8����������";�I�˷�p�\��3��]f��L۹�"M_��$Y8r���7}UJ�]� ��I�"$k��#W�59�?<za��^���,jό�{'�:�,����q* ��*�
�����ӑ_�8׍=���/��r�T#���N�]�#�Qx3���r�84����Ra�Vu*ˆS���Ti�V����zZ��v�����ه��!���׫�m��0�:�D�ڔh�F�oRp �*o����t~��Z\ո�8���HII�6g��mK3֍o9M6,`���ɩ����>���@��G��D�Х� D�:m2�K�\��`�RF8w�Y_h�u��!;���ζ H����޶��iS�������Ri��Cu\�
S-����v�;{�~ܵ�(�.y
+�d�ƶ"���� e��-NuF�[ڪ��4G3_ޛBy0+���rt����q�u��0-/��v{Y�v����y7kL���-}��P�K8�MQG�Q��I���u)��#r損�:Br.\ �B3A�
��D\��n�
�NZ{����xdO1�CiF�)�}蝀���QF���A!�$Ȇ2�(��:o�X� l��
��	�qe��bQ#$f[��>0���T�k�v�F�:��G�%vj��2�{���C���"�!C�roe�,d$����Ȼ�i�s�$��sK�,�x��vYs���s�DU�ʵ�H"aL�i$�K�_���;���6�7;J�[�ͅDq\im����]�u�2�i]����b)���B�x�c�ٸP�g�n%�^� n�=n��r������4�L�X�嬃��`��k�ƊÄ�����_8��6�m���l.���H+o�>���. �ײ4��)�g�ǌ��n/*|�(*���UAR�.�n���McK��ߩ:�������Psu�T����lF3,�s����q�%0��03�x�cr2�ב�6�7_eB���-���g��T�k?�q���,}�߇��:x�>N�P���i��򂥺��_����R�(�~Fs���'�|~����{o�	��BT�@F�p%��T�FӁM�J�\H�'z!�H����]���v���������|�q>owg{W� ��`G�M��P'�lr���� �+�Sł�v�I�{ٓ���`��G2�*b�U�9�Ci��|���λ��Ç�D@����+�̻t�2�x��F1�]Ј�l*O^���>������[N��؀��h�02a��M��
��9�N��G��x/�B7�?��t�*\�*T���&�[4L(Ż�!=���-4=1�bt������{��ޜ{�YF@�,����u����}m�D��~|����!���{�݈.�ߤ[K=G�̎�~A�`#��U�:Ɍ!:�UP��e����K�����m$t�M��̥2Q�NezF)�i +�Kf��uL{Ǉ2�;C���b?_�9�@' �G��RB{~�U��{�8��g����MG���V�)ёV�u��g`�0��H{*v��(��$� ���R��hKIW���4�-�n��To)�R����J�� ����	��O���(���r�r��0oO�Pw�ୃ}x�|���l�r$�v+8��f�>�W�� �S���09X�Y��K/U��}6�y��әS0������[�s���-{�k��#�k��3������\7�G[���K�Tlj���"~�,�h�8�0m5��-�}�zk7������э��k;���V�`�Ϸ}�Ѧ�LUʶ���Z_�E{���6ƛ��~�8�O�Csc����۶��5,�=;�Z���uqH�O�~�A�kZj�B��?+�T�+L8�Te@fU]Y\ T(��%H�CT0H閴qy�G��C�%v+�w��)M�����	mƾ\��44��KQq6.�QH��Q���͋A�(�h:1���nz�cH��a �Ǆ�*"��T��X:�h�`A|��[P-��OAJtS�SM)F(0��.�5u��u����V��%k������΋A
ﰧ��>�0S?��J�h[���̃��Bks(=��)ؐ��R��y�I �+�T���9���?*3�V��El���<ѵ^u��O�wN�r�hjY�� �� �z���p��1��Y8}^�P��lPf��Y��H���i7� �)-�8����Z��*B,����Uh��k�V#`J����3*Hx�q��ӪJ<���'��R���İ����7jDss�X���bu�<G��
�����0�]0=΋ԁ
�4�/KC��9ɣ'��w��)'�y��eǱ)�ߌQ3���
��T�h�A�����G�SS=�	iqz���lͲF3S�0E'b�����t7���}pj0��7��A7��
.��h�������p絟�s�;�"o�ľ����V�Dg`ۢ2�Xiћ��72��v���K����/��iY�� �2fT-��r+�(�dHF��b����$fB�H{�<u>Br<�^m�{�V�i�rX�C�{�p�9�F(/	�Á�>��/��>@ <�����ǟz�.^�b3��B5���\�v.^�S��O^�GG���������WN !&)J^XZ�����v�ɶ�yd������ܛ����k��_|�|��6��Q�09)\�౞ ��0����o�k�L�_Ȗ>|�&��k����T�* J��N��fe�7Is!�ϰv��(��{R��}�S<8�6��K �>K�:K8ɇ��
�G%�85C�t�81d�b�@1��ۣSz�}uVe1������^�L�����J���I���19k������`�Q4�s�/�i�v?�$�~6j�f଒ ŀ�N�Q�Q�]4P��	�z�"�����j�2̢��U[�!9����9���J�MriF�7G����0�\!�8)&���1�3���s�x8D����#8B>䵏DL��9�9c��j�)�J���qy�vd7D>�u�r� �ѹ��s�3�Bv�T<2f R_�\�dm{_K���S4?��r��nYz�/�X��-��@J�y�E͘ơ��V=�6�����j��\������}��K��~�⥣��^=�i�ӓ.��d���AS��g���G����ݢ�,N�&��㖻��Vh��F�'��:���"�2��iC�q�|i���;���Z�V�iV.��y�dy����������E��:8��Fo���ޤ}0�F��x����e�\Yu��<4>]�}�:w���9F�_"(�u��ܣx�$M����� ��JQ>+� -�=@L������lD[���+�DX�&�ֿeo�E�F�x+[�X���y�W�0��
^D��W�){� �ų�{a��(����E�#�"T�Z��iiyŌ��y���,��� )��x!U�
Y[H�b�1�6pE72���biO���h!+�c�j�hZ^�E/J�-�\.��j:�@냮5�BQ������E"#���P�ӭ/2.B�7vO�2�jTg6 �����U�J���[��.}�I��b8��5c#p�����xU���=@J�Nt�u@����	��1D�r:J�ц؎S�K�iy�T�4M�����<��~����~����P$��;�c	{h�����EA�p&Hzm��X鞈jBn�� Gn�m�a�4A��T���'wB��S��"�#)cw:��g�F�r���^ƩCM�j��K�m���&��~�!��@�(̼����	d-9v�E��;��! �51l852���1���	c�^idP
�H����B$�:JE��j�]�������W��
�����S�x�'���~�ix��-e+�dp-�K~~Ym�F�}������y�G��t]�y�y=�ꆂ3\�!e����_ez���D@^S4��)ۃ�C)��\@Pw��ex����;��.���k���88:����?���M��)�˫���<��|��\�+�6|�砝7��n��Aqu��!�8�N`5?�Y9���7(!]��~+���H��>v�
��/V���{��nBy� V�!�$ZP��ܜ��Q�h������
܈(��G��U��s����_[�n$��\I|���4���͏��N�'K�Gun��w�V\r��t'f�̇�O*���sk��7����2�.l6B�!$o�7kO��&�����:sj;���\�'��e�.;�H�2<|G��Da��(K*J���%gk2��Q5*bc�N�<���1�Cl�I�
�vZ�L�b�5
�����\�k��ǈ3�����kp��~���"�1�qT����m�aǣ1tE!�K�4H{���L8�t���M^̫�s�u;Eo)C%*�K�-Y~�Lk}<;E��R��U2} \���>ڜ�ɁxZ���y�x�W��~ȕX���c����N�Aaks$jJ�7��?��W�[�x�ڣ�~����9|�]n~�.���u�[������>x��9��As��Ӯ|�
c�k[��~7.���rR���v��6�����#�D����a�J�$�a�K&.s�#�C��`�q��$Oy;����K~�ꎯ~0��˓�w�|0v���t|��q5a��bMY�][u��1n#��;X��}���{��_����8��=���_����;Iw�T�4Q��f�*7zPښ�zOz�@׭I�ސ?c$��r!@ʞ}rSQj�*BI�lR�!P�v����1T��d�к>2N��9E�&��b
]��v�r�0 �\�,�)(�7"����e7+�&���'
'��yN��qɌ\���+*t�����"��IAi s��*.9B3�1H����C�)jSW��|��	D�%����y��o��ܘ�g�����.�#�RS>�]��(K�qkC��¹-�yZ.l�wRT���xƷ�TFZ��g
�߅O��w�V��x�����VF�>��h��Iΐ�� M��DlOEa�6ݤ�� ܩ����c���Ri�W
��e%\ܾ��|�&38����1��8���{��K�W<}�.�f8���HX�(�#Ox����u��[�x��[M��4�dtd�[���pS�>l�wg�c�St's*j4֪ͤ.u� gj ������:Y]�H^tJ�J@IЁ	�@H�0��" x����`Q+(�yLm��l"�4���#�Aky�Q��Q�}��!A��l��ܯ<���%|�dz~��
��><�K.��=
KR�aA`��ʂf�Jv,�N/����B�9]��֒ma��B���;e�9��Q��Z�! ��S�V]:���-���&�1bTd<���^�4<��#�ګ?�|������̏����N���0B�xxp����>�z.Ov��}�+���e�sp崀%��b��Q�1��Zʕ�6x[�)ZF�� Q2F��c��AP:���]��;PF������l�8+�է���Q��9� �pZ�t-M���۹"�mdi��jT�?�f/:�;�w�yy}-��:N<S\���������:zR��߸��O��1'6�=��Ȋʹ�?D Ɣ&k�/deK��4qϵ�t�2�i�X�5Ʉ�����\�^*S�\�߹d�Y��d�H���]:Ea:�:k}p��i{N��:����[݅�E[��J��m��e|��B�-wK*�s�Э�����KAӬ��]
�le��@Y
inݒņ*f`1�;-���Y��R%C�ZN3����pn�����/�ΰ�RF�lgL���ĲH��� �A����B���`�u�\m�?��_���Gv������#g{�>��\A��GG���ꁟ��l�f�������b��EWm�A�z?*���~&�5�d�y,#d�n�_Pv��,8Y�ýw��U���l���B�n��B,_�RL��j������ǈ��\�'[[�8�xugWp%>
R8� ���Q���.��|����w1�/���ޙ����P?���eW�R�hCd�bj�rT�@^jݡI��4��#+q-�˄Jk�(#�ĉ)�!�52�E�I�72Z�G�*�M<N�N�"�-{�p���h�<w��5(\u��h�� ET����.!(,8p�
����r���FC�h{~��y��19U�
dTpH�6�x������D.+�9�C��U5C Y�[�<�{n�-��Q5��L�zJ�vs4*��
^y�ܣ��+�Z�W�\/���x�������>@ax��8.Ż�#eEy����}�Q��;�wN��F;!&��f��SO��ך��y�k��'�R1)z[�[�~_K��*BZ?h<�B/�i?BN���t�."��M���4ͣ�Xa��e���So�-'wi=1olN'�uƼ��\�����/�ŭ]8><�7��7����P�~hT�H�He]-���(�~��š��i[K[��\?~Q���ϩ;T��*�j��H3(֊����jx���uT��v�5��"�6����H�W��0�2�[#�}.M�pڷ�� ��F�\Յ\W#[����w�b��9����+�U1�����#챗"TG��j��a���x,ŝ0`�깝� QA2�岁QK`� U��M��ZL�&U!��d���O���tT\��$�����������p��-x�W�[�]x�ݷy�!���s�Nrr� ��(V�8	H��5m��F��	Q_:-ʐ�d��C ��lQ:|[�s��2��4��#+[�@i�{[;�䣷`ow��k�޿w��%�f�VjF����+�E>�pa�rs������|����W��)Σ�(GG�Bk!��
b��ے�v�׭�b���Iv��HOl�lRR51N���Ŝ�ү�'�f޳�IYe�^�٪�sQY>EO6��?gۼ�;卑PK̎����o���5�.��N�9���w�}r9����q'�9��4u�����R&ɚN���Y�B��4�,�ЛC}�֪�ȩl�U3�VA�d:[�9aM&�^p�d��Qx6z]��W��z��.����$�z��Z	���)T4K	J�*|��pZ-eS�� �1�9�.�����?���G%�N=a���ȝ�֤�u�����3�P�Ȉ�N���D���jG���ӆɆ.��5��B�ZU�d?�v���k-�HC����[p������j�Y�g3ьR�Z���x������{y��_}����S�W��ϯ=�����L�Y~���߿XįW��3[�wfm�m(�r�"�Zq-s��Y$-�ƀ��h�;��lMWr!�ďQ���'a@�N��f���������׮�[���h���r���r�xl�R�9���/�o�m�w>7��������[�_~��uѶ�"XN��X���� ���2�(���{�z 6��~�D�����MF7��Ѡ�2��c��A[7����p�FU�Z4��2khѲ�H{{�|��������?��_�{
G�h{к����}�)x��-�<�fO�������������A� �߁/?�\,���M��`<t-�h�}���7aޮ`TG�5ށg�ނ]<���Qp�9��<����'��[�}�ۺ�(�fxm���3����^����}�><�<�s�����������������]^�[Bj�y�R	�s��gx&S}�R_���շN׫�2���i'����!�K�i�)�����z��&��1��y���&�7V\���길�����jp9�x5_����A��4R�n�B����c�G
��sF�JG�R/�Q�	@Ѓ�'Q�p\���Ǯ?�}�s�6qu4�5�~���:+�.3�޽(� \��H�
͌�j����?�>H����UH4���,;bL�c&�x��=�C��P>��Pԍ�1 Zè��Vۅ8٨�R!krh��t:���p��N�c�Iվ��z�@��`�^��~�9��s�+|R��|��Ν��?�6K�q�}�*Ĵ_$[vpV���p�_����������%+�L���>
$�L�-�k���"'8���d�gk�_�������#,�v�
�~����r���7o�o��o�W���|�2|��_�o~�p�r�B��n܃������_��`#�����	�o�� (okB�������} \ՐƊ��uoK�M:�"�y�ZKD��9" ����6��|���ƍ����mo�W���[���T�H�~��4N�!�_~�ǰ��/>�<��v�	|������7^�>O`w��[aPķ�d�uf�ڋ1��-Be%���!��5��s!��k%r1�EϑU�!Q�D`��E��pzs�d���\-f�9s,�}|�&|����.ά�;�(~J�Nv�/fԞ��@�~v���ϛ4����u�)��լ�J��?�ֽ�]g6��2�S�&�f��N�N�N*���t�R���!�(��5m�[#�5P�l��F�������i2h���5!D�����I�a� ��6��3@��_��whx��]��إ1H^Z���R�K׃�ta���1򟤖 �C��߷�1��%��;�4�����3�Ar���]v������u�Y"�-Ɵ���n�L�hbu���OF���-BK���k{a�Ǘ���/?��?��/���µ�?���v5��v8<�և�v���2tG[o#v�#�;Ա�z$*�F.?��cx� {n-3�f�q��Ҩy�������
RIu��J@�E{]q�ӕ{	�r���k���v���ix���{=��d������*_���>x�/^��+�燿�_tO7�b������e.{Ԑ�T�`Uՠ��1&@�Y�k/3&0��=/�ǅ�3�
��A�T�_x����.[���}x���Du�4�+��P�?�,|��/���n�_�/���!� e#�����ͧ�O}m|K�j�'�=
c�ڏ��r��h�0چO?�\�SX�8F�Cuwu���ဲj���q����O��y��hy�����8F�s�����?�#�^�����}xw�`��;t[��N���k��0>n`�����^ܻ�}�9**�zŠ�B5��_{�h�
4rk��is��=/��m4���rdD ��5�}p��"�&M���p����6�ϙ�2�?��L��,{����H�&i��tE1x��
���D]���%���A�CUi	�Q"����r*'��U|�hc���(%� �ϧ�I�� m�
�ʵ���P��hQ3���nZNwcϣ�E@�	yG%�5��ŭ=��}���@�&���`�!�h<�gp剫p��ux��c�T+.r��Y�b���(	�y�������x��1��12�wJ9�kO p��t��4G*�Û$�0��a���.��o�+?�`Y�K=Y �h�,�x<�bYqj�ߍ���y��Wෞ�|�_�K;{hɚM.z��y��7��~�o�{w�B:�x��Қ^��W�����.<����3��g?�g	�����[w� h'Ќs���I�A�s�А�-�_��".Z���@kX@e�k��+�MG}Y�yD�ɰ��O<�Q�����c`�����~��Q�M�Eo��6<��'RT�@�is�yC���m(�i��|�_�3Z��s)�h��2Ky)�å����ǒB���Y���"ix��%��K����=�����Go�aR�p<�ZU�%^�ջoC������1w�p~�/���w�'w߅��=X�5ϵ$#TN��=�?�i�<4*im/~��'��Sk\JP�Gџ!Jj[�	R��Ƹ$���q�,lqZs�ӛE���&<�Y(�~��S�C?�o�z��drH���e`6n���q�}�vPMt���Ɏe�����zc>S��P�[ � 6�Z)�M��d��7)��>1��?��]kYA�su8�,͆�^vӏ��TA3O�_�~a���דI�O�v���{�k�+��ߦ.�
��˴�n����A����T��H�-��ǜg㩀�n7=:�_�����UC�Z�C*�r�>a���15;��lH���>L�'��'#�e���Q�4��~@�V�(���^�7���W��������0'�ڶq���=@���HpNSe��u�tm�G�'��4�\��/?����֞��<� .ּ�Ӣq�g�8�Rw���l��[Yh]^��\ZSji�)eT*lJ,S�n5�DAS6�*|�Vi_{�ݹ���`���u�������+����A�?`x����E���ݻ�����+?}�y����u$$jk�$�U\&*8BV�"�Y��{�8���L�tY�����^S���(�UL��7�=|��-��Տ�4fv�ԩ9)�E�w|���;7��~��ǟ�%
4���h]ÂR:@Qy���y�W����}x�w!�K��ށ+.�K�>>���;@�3�hn���շ�޺�.�[�
9`�����m���\(F����DU�n��F�m8X-�ѭ���S��o=��x�;������߅o�q�Er�<��%|rr~��#H�-��1�1<�{���������a�Cz����>��o�n ��a�"^'k,,�rZI�M�~� ��A��yr#B
�Cn�i�mSD�}{;(�]k���9�`�n!�ׯy��t�u~�)`�K��D��j=<�w~��g�C~�U��b�[DH�TIM"~���ӈ���Ndp�2��QH��Q��i����#��(顠k��Zw��"EH	f;�n�B�
ڐ誑���} ��������>�|����a9�>�	5IW��@v���}y2��(Q#B8Y3"[�h!�R�?�S��ʗ63�-uh̨��R垕�b��]���n<���_�	����Ea�S^7�Dc�Ns,J�E�A�eNGQQ4$���g��Ͻ�<�}�x�u�nmqⅭx�����r���kѺ������{�I���>O^.�v������w
?}�N]Eɕ���&Lr_J��@�d��/m��iM6X����)BQ5��]��9_�^�?��?�/~���{����ë��
W�\���#<�>��%�!s�U��t%��0i���\rl��ڜLNs&d��=��'T��&N��ŕ9`�2�z�F��P#�!g����E�6m�Q�c i@��(��X{��O�į�ٟ����0���˩������n�v�;��-x��M�����|铟�{q���aNUyՈ�����ER��M�� ^�-��"�m���gǋ�,V���F��E �0K�S�;�:py8�E�鋍��)fϟud���}�
� �%�Z�h��&r=U����p6���oLSzFO���5|�oR�~�x�Y��V�>��4GNEN:N�>=S!3z7�H�ӈ��ݒ�+ć���Ӿhn�;vl�c��g��}w��l�6K����ie;Ǜ�*��Ps��z��8�PW��v`o2�=�o����wG�[3����x���g�s����e,d�nҍ��'�c5��jYލ���4�8+�lT*�����3�'g)8-B���
�A�2��v%�H�C��)d�;���TV�\TerF�2����=?�?�+���c'�脪��[M��sWo��{ORd��
���5�ߝ;wV���tu����-��U1�\�9IrE �#9/k$�5�uE�ޱ�<�>com@���!9�ٙ� ���/NA���u�p�������p}k��[���z��?� ���^��������o?��?<,�/@�����q�׹�>S�f� �G̓��N�\��iߛt��NVVwʯ�_�/�нVV�t�ꕤ�iǳ%Y�EI�ę ��ԙz?�}�SU H�Vd�su(���Sgx�;�g�SD-<�Hc�E�F=Aǲ��b�8������Q!�� �=e�} �Ϲ�ssM:���Ck�wt9��2-�L
�����4�jlP�dǳe�V39:<�N>���}y���MA�����}�4Q������-�q���҇���/�^d�����{�y���J4�W��A��l5x��h��9��4Z���if|���yj4t��m��󐍋��o����ON�Lu�Vkm����ش6)�ti$_������:GM;�O�H� �����w6����]���CV��l�����q;'R%}�H��,Rs�~ޠdϫ���C��9�В�Dc#���)3������8V��|�"R`��4�~-����RI�D:2�C�Y1vi�)�8P�֮ 0�u�V$�qQ6�P�J]�-`PEt�<��i6�2�d���a.쵶"�ju���R`I�1�|zYL���Zrsl�=��"@b�Y�f��H>�^�\�L[�m��[4	�y
3E;/�����j���N�%������=�pk�4�"�H	���7K?-a�&��J+u���$Q��X��DL;!�:[����\R����R.C��v�-5"������RԦ�;�/��/����v�y:r`�>�r�>�u�>Y�*�PՑy_�u�M��O�ky����?x��|�Z������to�>��	�Y_��<n;�4Þ�"�uT�`d"�:��F���	�P�|e�(��dOR�E?�F	j ��K/�D��.��7�����;T��ittT��FWV7(@F?�\�,߃��9�mC��:fH��9v��o�FMJ�����ÏD�HRj��͘tmOb��._�\.Q�A��#��R�Y�ۥ��!�9�@dz,YS*ժ6�2�9�JļX.��/�CY���x�ےo��y�Cn]���?:�:͌�Q1S��N��_�;�~D��@�a[IWپ��m��tQ3t���^�0 �]�|�a�N�LCR�@V���|�d`M}��/�0��`a�c��tD���)�gO�[,zڱ�����ՠ� �Agr1�=�ys���q�<�� �̏�^�~��g%|ܖ$��Hz��&������Cm����C	��>��5ٰq`[�{4}øU�0�tl�Ǔ��|�DT�Y�-c�h��U.f�U���Ls.��/J����S���`�c�� �A�Q$%_i��9�$>�k�t�m-׃��-�yaAA���PJ�$"Yf�����?JT6�Y�݁;���Lݚ�P�O�I�����Ƽ��-�Ԭ��ꆬ��4��d&���q��C�ƴ���N��~���s]�=oSSSI���
�����i�G�V����F�#��D"	������29l2���XfUt���4y����_j�����՚t�o�U��ٱ�s��V����y�//����^}����r�����Cg��D{
�+Ru�XI{��5(Q�H�BA:A��L�Y��$2�c����t�t�hq�|F�cI{�����p�D%^?�<��Z�Օ6z�e ��E�\y���u*t-:}�Zd18!�����CcSt`|�W��+�
"cj�q�:A�%6hK<�A��� o� }i��+uG��:m1����6������:����ᶹ߭ѧ��4àpa� ]��I*W����!���^Z�a0�`�ȉ������`w�F��,U����2��5������(d���PA�k&�~�sOr6�d`.�l����½ª�������3M�b���AJ�Ҕ^t��b��k��d�Bs��_P��"���hu�":�a�c���0A��n�-�[��v'2\P�ۡF�IM#���w[-�0�/EvOy���	�=��W�#��O�V�D����RP�R&�U�<;-n=�K��)S�R;�
��^$uY�v�v �m!j;e��m�8
	���Dj
{J�&  � Z���6#`��cB�m?��1T5o���r�Js�Z�p�.S�-H����!aJ�)��niB@��(��z�.���ߢF΢mh{2��m�A�R�y������[W��oc(��v�K7?]������ڕ~��F4F9z��s�湗i�4J������\���-����g�`����?�p�h4�CA"�z��L���H�����&�ۘ��	$���m����^ژB�"2hR=��^x���~@�ϟ�۷oӯ�kS����ܤ�w�R�V�6��(R)� �;;;���& ?[[[)��%%��713F��͡\�I�4)�f��f���	b������u�^'.^�HW�\�{Q̉'����|#--$q[���i�h#�?㡆(�{@����>L�����ߠ_��2�|cs��o���.S6���~����@��[��I�ѽT�
�(Y�9?����88�4��"&#�YnO"-��?&**��ѐ�k�Q�S"5C�2=Q8�~��i�aO��OUk����?����:�,7���҂t�2�Y�t�+�>q��������63�>n�)yD�ݰ�!!���gy<G�bI�L@���=ҟS׫e����c1�Y����[���n&Q|��6u���L�N���b=�,�	��j�˧D�d�k8Df����K$d>S���l@��A�i�(�9V_��t`-8�:n��K��pC`��<C�������$O��'e�1�P���1<���B��i�Q�?���p�x�`c�.������~�}I[�8�L��N�j_)'��#��\MBB��R�`����J��!�tB3�nm���3<��⒲T�l��|@A9�o��J�pzb��bݮ�Q=�{o�㧿�]�����Y?ȗ[����MHC,�(�p��c�*`����样Y��;��cD��J2H�f�}%���[p�tbvA
9�-/���MOM�A6bH�d����]�������8$�iQqW���ݞD�F&��+P�Ӣ��K͂C(���o�ާ���	c H9���Th���7����J�Ny�х�t��"l�*$�~��lR-�R+���r?`r��k�TF�by�2���w�~�.u�m�l;���SlĎ�'kw�AP�nVy�@x�s]_�P	MF2(�����B�A%�/�(Y��.�6`+nI�U � X���!��5����"��χO��Ƒ�S��:�5L|��_����u����X�Q%F����8"a
L��mх۟҃�.um0������m���L�x��lp7ZMG!����1W�Q$mD"=!
����#U�(iJ�i3�����(�7[���Q<�+K����a��[��:��z<���6ջm�|L;�z����'l����R#ʞ���++�_/hz�2LyX
��͚|�H�L��0T��6��� �v��<�����y�Uhn|���{�=��| ���i�t��az���496&�E;߸J�����JcՂ���Y�h�Bƃ�\�>�]7;Q�� �裇w�I]n+��9����v�,͏NRm{G2d�Y*�iCO���@3쩈��moIm��W&2�gίHs���D��/ҵjQE�j��AD\��2���`kaa�������ӧ��?���{O΅���EZZZ��C 7�M�v�6,��ڮ&�2� �L�N�'�DS��T�; ;����Zj�c3̹������3;v�XZKPz��u�8 *Hp��:77G���*9rD�hw/�0�|��ԛ� �N&��i#�������%��@t��Mn�*9�9E�@X�>����S�Z�?8�
Y�m��q������Z����\�U=!ȇ�erR��~�'m�(k�кTp�e�vl��$�E(��f�>��.>U,ۘ�j���Ο��HZ{�x���"J��퐤 A愤���5qo���3z?7����c�U����'����쥫D⬁O���
�[���n����F9�eT�H� S�On%�=�ٿ2s=J"v4[�N�kM��O�<�ǒʯb�JWV�3R@��󑩁�Q���	�����6k~���9$k���<��Q�G2�1pE[��CA( �f��|�0>�a�rd�`w�͆�R�m[��n�H]��7�BF�!q�,Cl����>�M��4��Ir~rc�Z����زeY_ڀ�����dn�N��j7<1n�M��(�ү"U
*rs"K���d�!�-)�F�]�qG(�׫1�g(��ّ��rv���u�?]__Yo���;�w�?��d�rmKx^�Q�gC��D)"L��T��gZ�9i�g
�%WZG�aM�b\S,v� ��V'��R����bhу�ezȆ�xu����ѽ�U^`wiێ���W���)p�0Jű*u��C[�)W�R�	�<U%I�C�i-�P��f����kl8��UrEW?O6���[+��FKk�&���B��N�16<���4}�o�P9vL��j�i �T6� !=�>��J1�0(|���e�?o)����$�t���}t�:� -4g���+��#;�=>�/ͷ�K����:�y%29F��{�ġ�#,����c��)��S ����>����Ut���`�X��+�#�P��:��^�p-$� .jXxTd�[�����yW��n,R���:I�@X8[�,���JU�Cx$�8�@���D1�"�u�Џ�Ro�5�p ��Z"���(CH����$X$�6h�4J�J���B���b��E�b��+Ԣ� "����n/�#'�SK����iY ��+�H��0l�#�q�>��:d�}��ۻ��m[��dԄ)J�ꙅ��Q����w��NȼP`P��W�0R�(<Ƥ̀�C%���A���f@��6�����tom���!QG���L�6ʀ��a��������4k̀m�J=m�vH#��^�#�sFz2��<�M��%c���1�^Z$�ӣ2��N/�RwA�"�^�%�R��P?
�9�
��1�0��
�x6Д(H^��Ђ�RO��6S�z�����$�`�� �_���� � M�!��a���= FI-F�6jd�y�wW�OX��%�{���� v�ԩ��"���ŏ>�H�0���D���J�"��p0w��}�0�> ���<��e��?�vH/�uY�t9"���"���&��m�ԯC��������H7���kH�c������'�G~/�?|�u��.���������i���c��1�-�D���Y�JEYH�2H �!'���y^ �L�KdmKj�T
���X�btj��������'m_�5��]���ދRR�Nl���� &�ELC�_0 ~Zt�J�y�i���z�t�!�@2��~��;�n�G?ѫ鰍�W�U;��?�ba�Z2�����~��p��u��Ud9�
�&l���	�;��;V��0-R!E��VJj&:�X�%%�]g�Q���	�C��*�\����3x��Y�h]aK�>�꘡�������b�rd���☄3�����?[ v$|����v�m�~8���{��`��o���}�>���{��Sαo�P��C)�ǉ�Ƙ���@�r3iE��Tѽ�}wwq'�u/V���h�jZq��o�!��o+�*q��Ƒe��=j8A���0N��I{&���Df�_����K޾55��w.\�����4O�v����^�X�^��ڄ���&�~V�ʏN4(V�Ix3��}@h%Z{�5HU做a �
73�]^P�v�i{{�
l<`��9ʆ�>kM�e����ͪt�-t�,ˈ4Ā�[�0����Y�'�5���٨C��x�*7���xn7j��iI�*�|;GlT;��8x�j3�u]�A��d�Ih��~A"�]+�d�;G��P���k���ߤzЦ,�3?�x@�>�	F�����``.��#5J�ِg����g��8���R�e��opq�K���|��m��N�}j����\����H�!�.��>zU�GH��ƨ/E?�(T�ϖ"G������@�˗W�T"��QE>T��
���� ]�e0�°G�������B�Hu�$�Yd%�V���\ @�?d���7`���@N��ԃ�h9�#5
T���I�I�~���D���B�	R�'�R򅜒-�yG"�H��` �1�et��16��bGv�2�1�a)y��Ks�u�˽{�徴��S���h�s!�b�ٌ\�+� � 8���hq�� �Q�Sc��a@�
 	 \KK
�R�"Mߟ#X���Vde$��c,���x-���!��ERyT�J��ҹC�����<�\�m7)�9��cr�����U\M+t��eZY����Z���Ŏ6|me����G��]q�Ta��;���n�Z� ~%������)2dJ�?f�<��_��<yR"k׮]S��� ���@�J=(T���f��|-H��63?J�"_+<k�]a)����BJ��At�E���8>j��Æ����m�{{wGҔ�����k��xO�{ ��'�k��� w��{�}�>�xH/]�ó���(��e32O�"�Ck�4�h=�����7�ƛ��G�^}���w���t�L![�n� �,�߼BG�ґ�<�=:�$��5>�WZ�4�=�Si����jO�E-����"�X�""ay�8A<%#�H���ĮH���I�g��3�~yN�}7CD5�ޞ}�I����g�	�l�F�k��n�5���_x�1m������}�m�z�ۯ~Qg���I��� �B�Y4(SA)X�u PQX2����s�� u�K�tJ����0_F��[!�a=��� &*�[�7b�)��8Nᘃs��ps˒��^�X��5	5��a��2��nF��B�p�܃WS�ֵz4vr��f]�9������:j�|�]�gg��j�&R�k�'u�ź�3u���rO|�'Uܲ��>9v��2^��b0�lp��cw���y�ۜ*�����Z]�u[w��w�����q�[6J~ ��u��a��&��~�ĖTq�^d�Of
?>92v����'������������;n��?����8��3|碧1�/��T���\"1��O�ƒЩ'�����h�T����qp@W�w ̴�Ɏ@r��!<w�����GF)ǆ���Y���$BϨ�˰ѝ�\J� n����6��0��U��~`�Wf 5���В��2_k��� l�q��ԶS��:?D��g�'��J�:w6iec�N>*�o�Æ	 ��(b�І��ʌ�)�AS�}j /�ϑ�P'�962ϰ�>��҇�	gI�'
�7lX����Kt9��\��D����M��F�P�ֆ���c�2���A�D%�� �s��iߒ~b���PI��N.*(oI����&����մ��!Jѣ�4ơ���Z���}VR�Ba�,���7�)ҡ�ǅ����Cyge!���MC]W�H "�F�%D��.*i!�zTrø�E���XHÃ���Ǹ���껲�78��f���� 1\�X�Z[��+-j�f �c�s���t��0��\��@D�X(�H�JkVxL���G��Q���\��h��	�Y��_9�"}�?��VCꄈ<��X!�T��g�M��k�rx�⼱<G�-b���C[�00{��F���T.�%�duc�6k[J"��$m���@r��0�i�(p �fD�Ezau�T.*Ra�"�����4��~D�ז�veN@
�7�������i��[��.�_D�`�+���G�XxЎ�#��������:��cɄ�$B��eq�RX�~
Y���\F"�`}��W�]�pA"j�=����&�WDiO�+�0TpR�1 k�AVe��?��G��!��ZD���w 6D�iD�<��2�.c� AJ+��O�S�TFzL��}��"mHe��z�.�:���q�˫�������ᩣG���3ZQ��}��NM5s<��q&I�b�셓��^y�~��/hw�N�T��c � ��w?z�r/~��u������]���\���-j[����28ā2'˥C�g����'d;|=%6���%a���'G4���j+���zR5G�HO'@�
�X���o}��}��Q� E�j��#1�n��~P�y7������?�ͼW�m��jՌ�xzܕX:�ё��T�t?�h�����X�;�n1��G:�v�r�Xi|ƶ�v#�k�a�V̭��9Z:F��HiK���G���#C�+�����TD�I�ҵ�y^���.= ���"Gd��Cq��M�zoe���;B.�[�m��L��:z�NO.�:ӕ50�t8-���&��6姛���Cќƚ�n�#��%����z��m�A��>��>f��ౌ����i������W�n,�x�{�{�b`w�)D�<Y�{`d����)z6�I+i����j˿�;��-+����a�Á$3�Yl����B�Dw"��iJ
h��A�L`����|��W&N��3�͕���{�o�nw����^�rA�Zr2���4c%b=X�l<}�;E�c��5�0�HRԛĩG(��v�&K:55Oc��DD��FG���3�N�啻���ŀ�')�#H�DYg����!���� ��A����&�_�9Gy��-�q'a@udr���(�u�*r_�����#��b�Z|�� @t�Difsy:<=O�l<tD<6��H&/)���b`�$����L� �d�t��-��y��#$W̆�����ڵ|��Y*�<� ��K3^��O�����ZJ?"Ҫ�S$���{�����JM[� |�ϖ�=A|߀B��	��jC:R
S��oa�=U�-S�G)`�>f����IOJ��!)�n*�k��� "��R��(�PR�-D�zTr�*P�x�w�� c�4��I��
�.%E��@���e�S���F/d!��Q���i'�-��xF/�[���{��Q��`@S�1q
��A�3�SjL�ܷч�S��
�zd"��A���(�A�\O@,��-�("C%6�ᩰ�_,�$���W�(Qn��nS��0�ǫS412-@�%���Vug2�I2Ru��&h�l�Af�J�R�v� �<�顭v���D���c�M��8�=�#��}z��BwvWh7iS�$ڎ�k��F L��<~� �l�F������N(L~�BIE�@���r[����=��t�:Y��P�y��Y��|�������=#2[HO�#i��D�\ICU��܎�z�M�v����~��[]��}�|�R$� ' )�9� p�����g�g�WP{�tM���֭[������� �q% �2���5#��Ы'C@�֭����i���~Gd�ϐ̀��7��^p+�|"M2T�lH�}7�U��$�k��>=3#�������q�>���&�%E�G:(�d��J=��qWd8�<��T�K5��z��Y���w�ux����h���"&�x��~���S)�S���'Β��Hp�-���. �x�ej�I������u�e:6{P�K8��<u�i�Ѩ���P@�D�C�Y���d�--� ��Ʃ:8�>���d�1I���7���f�����9MMJ�4����e{�#�A��7%�K�1]aX�m�C�N���NC=����-��{`2��wr�m���c�����j˥��0�#�͑�x�o��d�m��&-r��-U������D����׏����feEݯKs�掸9z��5����J�eC�O���gh�2F��Bjn���
��4�(ztfz�^�X�c�T�C��c�-�㣇x�����HE%%��U��Ī����R,�	����&�3[��)݁*��֨���lV<(�2���ne0��+%�t$��I�ю#��{q�3P��v������>������>�f2&Y�"��;���H�'��t�L/ބ���QjG��̈́���L�����_f��~۷f�����ܾ�p���^r��r��w�5�1��������N�bc�!����A�Q+��"��l;�	7O�1�b��6L���QȆ-����N������[<X���e�J%J�H���S)b����]^�C/?Ecl�(�R�H���FˑT�T���Cm��_:zZҶ>d�`��^N"�� �1pn�1x��c+��YL.� mn5�S�P����	����i�]'?��0�,�'���Z�ޠkK���D%u�;S;���0��������{�d�R��Fa���A�a�pwl�}>5p��"J�E �4	�8>���~ۓ �a�5G��I�G}�ͩoK�H����@JK� �0x�d$R����j!�O�9� ��f�uB���V��1M�"��|e�#�u�0JE8i�(V�c���6���D.J�W:ܧ:���x�����틄I&�mvئ�%��hj%b[�U�!��a���/Qʀ�X,BꁥW$-5�����F�R��� =�@�m��NC��j��� غ�nh{%���JE@���0$�����"����r1O��π+��W�"�������=֊ ;tD���}�$�NH�k���nW���4�<�}��|���ab@���o�4�Q��߸[�I�@Iޣ���}l�!H'�H��W�r{wi��M��K9���&�R���?��x��><C3��}!7���#�2��r`�FdP�ba�E���eu}��s��;Z�C�aW%��c���xY�g���[R�������O�9 d}���?R?�4N������fd#����D�@s��ʹ_�M�b���s��M�  ����&�ZM�����[��*�ׇ�K�!�HÜ�{ �,�!��s��w�����<�.j�J�c �0ǀ?�mg����������-Z�ݠ��\���������M�_��&����3/P��;��ҹ����ءU�i@ð��G��iB��S�
m0�Ƹ�sMx&��x�8��F�_��F�,J�4�á��'��������\��w��r��Y�^08���苻�'�����Z�y?���1�}�"��|7�����jG�~�0��q\�	c�#o�6���7'Q-�-����I��vU�X�xs����ߎ�9Z��ذ�G���Ht��G'G�鵃�i�����h�U�l��R��L��KG�Pv�@+2��o�}��O���{n�翜Md��|�g���X�?�y�m�⨄�]������H�ܿö� �pa`hi�n����5v���GZ�i���G�}��Ϻ�^���p���>zN�� ���C3����l�B>wӱ����)<DH��62�^���lэ@��E�v��:�0��D�	z��J;#V���*��X=�Rd��N|c,c_�L_�ꓶ���N��^�&���jH|4�p?uK;�6���.��x�A�����h�uZ>U�St��)6F[�靛�ުSYr�CY���f"���4 +cdȕ��a�`D۝�	E.���h��jG�<F�?w�2�oP���������<\�$��2��>$��^'�k+��f�\�n��s�t��I�����J��[t��]:21Go�x��
U��Apr����}�[�6H{ܦ)ϰ�0=A�c3t�����L��#��(�F�J������-:T�o=/@��a<12%�$k=n';ґ�DS��q�"��y^&�&��d�b�E�`FG��LB���'v�'-������D����lN;����*d�����v� <�c�8l$N����a�9�`"Q��ф�;����3l��b0�i�1�	!��@�O�U�H���!*l�J�].'6cCM�u^��\����H'��rq�S�:Ŧ�`�ry��~��Y�LD��#��p�z><s�?͸)�vv"�q�8��`3��HK�U �`��׌4@Dr Qc1>9I�l��:��ౝ�{���u4��u���p�lmm����%�x��٥��:�YkD��l��4��6Ȕe���O5�5�rd�]����D����%��%���!
�I=���,�,���1:|� ��]���]n>M�^��o����<��Hk�-oo��<��.,���U��{��S��S����<As�vy�)�	O5��B��s���@$�T�����_Q{��*C�G�3d0� �#�/T�������u:q��á����~�3I�D��� -�N��2lϪ~ږ�fqV� e��T���YY]a0xC����4 K �&�A?�~�7| @�0 v�s��������$��t�lV�ý��M-[��`��rI�2���Kd��S4oE��Ta0�I���\��q473C���������S繷LvΕ�my��4}x��̾p���l��K#4�@�=�Eh!�Y)�	�<�A,�#�V�?��=����|��>W�㸊�s9ڰ,���6i�Հa>��J�7�����'�4;S�vp���'��$�#���/l{R��On�'?��Vʱߦ�a?��o���?9r�ed&ّ��tH$:s r]�"�I��dI�����z���t��1)�����t��]Z��BPX�9�Pm�^9�c���ڝF�*^�LL�yCYca ���
��� j�ᘽƀ���]��؎�9��k. E��(��u!�.�U-^�ȒLBǀ�4�R�V����� �2�^ي}	eRT�P?���#�����Y�y��M�g
���;͵:�+��� tt���AY��H�0|"�!���l�*&���'�=�[֫6'��˫~}էd�'�-���3����'b�*4`��!�()6!�э[��X��B��щq�?�@��ѭ�ej���@a�����m0HD��<��o��|1�Bn�@�H!���W�&�˺T�zyu��&��܉�4^�H�yut��<9\]�MKl�Zl��[ts�6-�}���ԋtxꀀ��|�f���g�х��8M�7���
�st��M�MIG>���ߥ�wo�RkG���[1�`�����;�a�x��SBq]n����ŕ�������g�����S��u�>�]n�Ov�V������%�ݳ���`�,'e����R7��ޥt��\�Fk�Z�='�桯!��LJ�p�T� ~I��Yԫb0[����2~�K��uї���T�R�L�BI"���O��m�e��(3�H�7�B��o�R���J/��43sP�!��4�6n��"�ು����A�O�&��f���Mx�_�R-�A�"R�_�	"b��	��ٹB��9$���{*x�17s`F � )
,z8_�؆�-��B��"��:���35���x<��kB}NDF�#e��Dt,�5S���B[lq�l��VKEΤ��R)��v#Z���; ���Y��a�x˺P-6�޾�!�2���?@��.��{�W"D�P�7�����{��ñ��C>��3����-�S�����gQ�爻�!�rvԦ
�,x�]�3H.���p��.��A[�]�mR�Rw�!t�0@A.ڴܪH{Em�H0�i2�����B����$���/Kd颸�*��P�0g��3ԟ�0S�Dq|��k�t��� l����w�a�� $q~��KE���L�J�H��#G��n" !"����s现ɢ>rm�!9t�*HY��,���H����8]�֫������ee�B�f�N=B�x�U��_�+���*�6k���Pv�B��/�l�J�S�2��@�4Q:��(���5X�j<N�;E�}h"k)M68N���2�����<�u����Q������@01�����_�Y�y�)��OG�ݬ�6��j�r�$��_Q��>���Q$GQ2U'ҵ�p�����l�������Z��V�6ن�6m񺻼v��]������!�H���;����):{��2���E�� )�\�рW���<���.��
]΢+���] I	Ef�~��Z��52�r߆�J�9�$�	��dII�����.��?�o?����HR[A1yf��uK��|�vk��9���V{|�57�:�9���9��g'K�O�Q@po��f���HD6�v�*�LLm�3�Ź�?[�sseݎ���ߑ|c�a �C�p  8 ����|P�����{��BXƜ���.�����^�L��]j���@E��� �;;+�����tA5�^d�����I��]��H<e!�d��a�򣥛�:3}�f� ����-��r�>}x�V{5
��DY.�ݑz���D��H�`��.��<AܺB�Q��Q6�{���"����F���	��OV����Y�J[<q�r6��X��\��Ѽr�>Mj�]���L��|�s������}6�p���l��r}�>Y�E�mܣ��E>� ���1Y���n
��<����,z�C:y��s��fشQp�x���T�I��>��F;��ko��o��NW�>Rd˫(�K�ƺ�������A��9s�光�����$U�#���Ԗ���4<5~�5
�"f�L�Uw����)I��|6@u�n�{=���mu�z1�%���j�,Ԋ���O��lU3����3����Aӻ�M��[������m*V*���Td�����߁2��FQ��b�מ�G�aJ��$d:H��T*ż����f�x1*ߎj����p�]��DD(hb���t7�1��
��(���F��	�SQ'KR#U��E�O�ՐwE�������̱S4=9M6һ�w{mI�����z�NI�@�~��僷�a 2ύW(��	�[Z��M�oR�	ȏ;T���5�
��J(���]���)����GHF'}Wڀ����4�W�@=��D���k���~��\NR�PS���	 B�a��}"@9b��&Y�U�R!�%R}��/��7>����E�)����
0h�C�L���F��I����x��	�W�\<^�61~-�<�i4%%�US�MDa��Y)�����;�h�D ����QI{Fo��hԧ�X)�<������dK���Q/��Ͽ@��ܠ�w�K*W��!H�Z�Xc���>��y5J�ep����&��	U�54,=�f���#m� ?��$P�$L��U%NFƘ�p� �Ta������tu�s'���~r`��x�j�j���fiT�j�?o���GԀĎ��L���I���i胺������d� *��Fz]2��g���؎.
�AեO��&���Ͼ,�� ���� O�<�9D��������!��#����f�x�x{��	e
Yj�ʑ�@.��L�L�� {��4'��o{��l��=q��i�^P�h�?y{��R5����@��r�M�3Q��͖�Zl�]��\K�����V��AB���I�h4��B������Y=X9ءgt{���G����V��^��'2�O�&�e �������:�S1���:������L��;����`С���^�!ך�w�]�+˴��%���8�R-x�wV釗~MMa�d#b��JSj"Z����H��ܡC�4;9I;;��إm�i����t+�:m]� ��^^�7�vw��m�OP���%n�omS���lwi*W��:O6;����.�Hqs�@j\��uy�]Y_�vP�� ��	�#Z��60?�������|�*�.u�ν�6mZ�o)'����<� �M_:�@&	1��9�	�S��t������]��L����>�ܫ9دwT���~j_Cp�h62�RR��1�ɖ	�f��+���ow{��/�먇Cqw�AV�,i�#Պ�T
�FM`��4qz @a���Bj��h��^ML����ɳ���<������A�ӓ�;q��+w��M�ųƢ�"�Q�ʍm�tH �R7��<�D���#;�ȵ
Xp�U�A�_���������������޷�nIm%���$vFi��,��M���
�?e��Km�0X��/�� 걸M~]�/�|T)� � �w8�T��Y��
Ѯ"@B���{��n�~y��>����;�L�l�jm[h�m+#5�w6���G�֖���K�y=�֛�w����-� ���cf�:I�.
G��8�Q�V�hek��u�������%�C$�oPs[�C%��H|/]�IS</��ߧj�Du����J�(���)��@���,�"�pi�tت�%6hőCfee�~�ӟӽ{���{��/�@?���\�%�p���= ?�b����[NKL�T�0�m�4ƈ1P�����t$�T.˫�?���s�&*j�=��� 9[E�]�� f3�}���him�6wjT�?@[�� ���}�Q���He؎>�����F�<U=�?1�Ge����ϯJ���F�ܗv�0��^O�_`p�����&�FBD͐v��x�ݡ�+Hڸ�U�z$NL1�-ap��|��I1�Iݺ��o'T��"2���O=]8FKY�k�a�����b."����bN��CV��������v�FԑS�ȌL�����r�˴���-����ʶ$��:�A�i�ԑ⩁�i`K��i-�~}r���� ���)GR�ɺҤp	H�¤%+y&!<�!«�`�շ5Ƴt�e�T[�
��-m�D�%��w-;p]�c����FKծcYm[	W�\��2B(���ű�X4�bR6>=�y0�y�u�k�pv�y�"֬�4�9�ԭ�}_HՉ���P���Vء���DC]�	�����$~`��h��6�a ���&�!rGtmP���(������ �ց�'���
aM�Ѥ/�  i��UK�I�O;|�ݬMݼ-�p��9����ȇ�"o�W-p,�QDd���}��	�d�:��"�;5�#�9��}f�D:��ҖS��+��x|,=�+Ҁ�L&C��>`��n���N������)cp?���jI��F�ŗniP�Fn�<��"@p &`��.d b)FԐ�]�����k��D��G)��6��S9����U�:�EN��I/P�~"Bz��&t�Ds�>5�noR�שZ̳a\�c�S�ߡ۫�(σa��P��o��l5�P��o�C��/���eF���aNFRV���L��-���l���s�j�;�^�j?ז6�z�t�mUe+)�vb�ɦX���a)��T:��?98>�Z���sh���4�\���7K�����/�p.Wf ����U��HoԵg�f�,�=R,��D8@WiŪ��#��gІk����J��WE��Ց-��b �R����N�ݢOn_W ���f�T��6�Y��6�k�������4��ߧ����Kw��k���ƚ���(��8~ ��W � ��n��+���`���/��@�A���J��"3�R��d�:T�8�D!��\�V��4�*
�OD�Pz�.���qQ#�h!O@ь9��)���[ �� ���|��I���������= O�׀P���M}b�%�L�R�	$\�@"��K}(ҟ]h}1(e@}��Y�q�y����RToIT5k�A���z95^�w��"a D-J.��<�������+R+��p��5��?#uȘ�ͺ�:�~���t�5_m_m_m�n�ɶ��?�R������:�)]sI�� a�c�V�.�y���yЖl�<�ɪY9r�PQ� G���Q`�E���5O5uta��WB��6ݨ�I����
]�q�jAWJ�=��x�ez套i���2���(�s�m��6�o`�|�~������M4`�e��c���|	�|�v0�CS��;?�}�E�H9�u�����b�ɖ�߳��p/a�y��,���Q2 ��𣨛�E I4P�oG��>����[&�1 t��D��E��>>*9�[@��!p1�-�0[�Zl�I� (ʋ>o0����0��2��2��8IS�ж�q9H �ږ���x+
�j�`!Zf���ь�+}��KU;K��img[�h��q��&:r���Gin�*хQ���&�����8+^�l��"�-�<�
��Y�T���E�D�H����FD��g��C%`�(�Dx�!"���"	��o�H["a��an#�n)SL��<��{������Ha��,��#ex�^l�;d�����5u���=̞��n�X�3���@RX
�x�,G�E
���6_�c�������q�װ�չ�5�9�(�a]5�}��*ѿDR�,�nCH>�}l���,E=h�yrܮ���Vx�N�UګTۂÂa?�n����=R:�%B�oƇ�XQuŪ=+#}�'/B�0�Ӧl�G��"=��Es
�ld.�-Z.��$�f�+@졸c�B؁+9�諎�VDjG�����ԃ�{}�n_ؔ�n�-�b�����P����(��L�� �g!�h�Y�V�D�"��L�b��V��✥�"�.Or/P5�yA�P>�P�����	9@�%.a�t�<�}���p��j�����al��Q��A5V��8╅S��Y��:=US*�%WiT�ظʸ��D��jBDJ �V� �a h�ܤ=��1_K�բ��S4=5��F�:�UGhav��o�Җ�!�[IM����T]�VӐ�H�+_�����-�Y�� Q�@
2_�x��P�h����P�,$g�?�H����	�P���#G�Hݢ9�a.E��\fQ��� jQ?�BԤD	������'���HE��IM54�9�0�F&M� ��dX�Ǜ-`)��Zm�ɹ-��W^�������6e0!s��dMH˗�����^�s���J�p8C�P�6ޮ����*�']���\�Y����V��k ���KZ0���Һ������F7���HGEhl����e�P?�%�Fb�+�aR�10�������:9<�[��|�l
��Éf�6�5���j��M��K>��/�1������lҏ���v@^ӐֵC^�x��Y�X���Z�uB�N���2� �j0��:�vtj[F�qp��:���T��m)��(�s���o�؆���_�E>r𽛎dZ��'�ƪ���^�%1׍�$ӡƿAH�؊� ��b�BKE�� wB��J�{�6�����Q���> �r�g�]6*bWj�$E-F�3h���&iɀ�`L�^�S�9�l��yWX�"	۫�v�ˉD��YX�{��Ʈ%�� h�Ź�8�z�,9�,��;��v�D2��v��;	����7�{��<,�N�����}Zln�jgW�m �lݧS�1:91G/�:G3�2��6������Zv�D��Oxe:��;_�#a2L��n���{�����m�\��2�a;)GHgĤ� �X �1����=zb��J�$P4�����.�C��ؼ)�NS/Ӱ��\�T"LM����!	���#�j��&���{����7�~���F���x���������<�k" @w�)�<��l�e��Rs��H��F��L���0�u;b�!��M�mp԰9�0lw��ב4_�� '��ݦLo����})�9���3D�m�d,}sq�g�Kk��~jl$���{J6�M��� �Y���q庤N:NH'���C6|��Z��0���D��VX��O+Qb�1��l$G~�����%�uju�l@��jxr��I�4�d@�&�@d@mi]ʔ,�Hu�>�pT}[ �]�i��*��R�?��TI��n��u[�l"R��^~Nn�W��Q:up�
��xtmq�B!���R�C��+ 3��	����sѶ�2 ^e:��
��*Ti �����yܼǋG��p�P�k�Q�����^��-�{�7)�}���N�~	g<���� ذ5�o�'�?��o�¡C"ar��]$H�!�2����<#�N���Rm+����GyQ�i�����0#����O�EA��s!*y��E:|��� �a�&���B\����}w���$R�4,� ��>����.�h�H_��Q�B!��o�Ai�h���|��P�m  v`�7!��ó����T���z!�&����������/Q��z��:��#mL�����?��-���Uz (���=:pj��L%�S�G>��{�e3i������y�ھ���n�x�� K��c]��!�DA�&�k�����&�;�G$�zp*!�It1�i�8<���<>�lWX�������ȹs�Y�e܌d� ���r�ۨZ��ow�eÞ�yƍ�� ����n�&u	i�N"���a����sms$��9H,q§���p/(TQ�G3�랉6J\���I'�f<�$cP~��c�����Tg��أ���3V6L������-۵�8��@ RX$��jS��Hʨi2���H���V
��؆���o�Ž�崊n�����tZZP��ʻm봾>���W��i6)P4��J0�uw�s�$�-e��hҰ�M�D���=<P����?8v��ù��]���o�GmЀɳQ9����O�w^~��Ƨy�WuQs�^�珝���oѻ�/�=�u��?=�&�x�Dֶ�-�l"U�����l���;?�.#�*��џ��5h0F4��з����wW��*&$x�u�'ڇ#6B�s��� h�C��A��4���8�IS���C��o�s�i �|�+���p�����n2�-:�^D�F@gG�[��б�9�.$�aH�M�?D��W4��w�����bRS'�m�э@� "�V��	�~��.5�@�e������ZM�T�'q���$��6�u�NN�g�ؖT�G�M�q��/k��,�+�l�#E{G2������0P�	��-z���r݄�l����]J��b�e�9be�[����R'!�2r�ɠ��~���B��9��8O�"����|�|F-�5����Ṙ�me�JKzaQ�BE�#��$쳞:��yn@vPc ���w����Tn����=� ��z�$t��,��׿'BĞ��%q���U�0��IG�$*���M���B!mi�J��=G���\	✞p���^���O�}D�<'���J=��C����L��w������3�۩o���C�!��ϒ�iID�dHȢl"���u�G{���]C���%M��	4�A#1H"cƘy_����[�AK�Kܵ��p���ۿ�t���y� � b�F=�M�)����/_�h"@��.è�.\��S�Rdi� jM�����=�F�L�8�a�SdA
�e�v���2)����AXfe���W�a�/R/ߡ��Y}@76We�Cn���樇Ep#) �}�Cʆ�D��G�I?�0���"%T���,�����^�%@*K�"�-�:˿ڞ�-�%	�mŌU�M(��!GإmY��>E�c�&�}ɾr�I��Q蠔̮r�A�αm�־�-�WU���J&,h��"'�1��Q�G��@n��Ih'��1���hlc�<��f�#W1T�|"Edm��PlTm�$z-M]c��S>]k88u����t�a_7P��|I�I�ژi:�ӟLz�Wu]8c�$��J��+YVi�ہ��3��~������b�%R���d ���u�	�ca
Q�b늀X!��(����(N� 
�X1ʤ�vK�Cq����6ME:��g:�:�����Aƀ�����S/�KsGi�2&Ž���`Kx��x��v������oЉ����uz����˯���);HW{W)[�i�����8ͳ��bc��W>��w�P,�ك���ϓ���V����?p��u�E��!���E�i����������,����M��C�ظG4�K���I�D�t�l
��1��iu˴��?�4(���%�*�����&Ŋ�O��?��M����o��xv{.� Y�r��܆G����T�(L`�^[<\6�H,8J:C��L<���j"=D<��N��q�A�(�b�S�����YJ}�ʽ���z�g�)��Ve^�����.�+c�����Ce<Zi�ҿ={��U��`(�\qU1��D]bq&�����#*�"b�1�P�����~�T60("m%�����
L��n=K4Q����B�ԞZ�Rdo91����U��AS���Jڥ%�����Y:�+�K��4j�3 �(h��Q����!2�됇T�v���E�FW����۵̀��}cWR}c��Mf+Rp�qu_�>���I�d� ��m,�W,%�у�ZS(Q�5������ �K��r���ْ�3����Ր�w��dy��Z�������*�Ta��h�ҍ;7i�]�&?�6���"�I쁴�DK����7���K4;7G�SS���o������?���%ݯ�T��h�����(}�)��LI�˷������������I� ���ݡ)��2�'��|�9�S S�c�P�3���ϟ��M�C J��h#��{�rvvV^A�SUoX��Q�/�Ѻ�ѐ4��>	�z���obW�=0n3ٜ�G�;H�ZklQ� j�Yk�_9V$9��
k[� ��C��vlOӫ琖�ZM�p����N@���W��ٱ�A�i`�{��Y����I��W*�Z�"�:���Y�_ؖ�ډl�u�׃a�@$E�"n�Z�,��RsH����6��������TEMy�����ɉi��׿A�j�~���R�)�����+u�bODTD*<�f�&���W����K�F�F9'O�ߣ�v-��0/׃.5��_t$� � 
���Wc�a���m��O���yk��&ă�5l�A�ߢ�=����H�Sa����z��7�a�3��;�&VՏ�r7�����yQXFc�TQ�'�YzƷ0�8l���Z=(}%��}�%���������GD�|{~�{ p6Ly�V�ը9�5� _e|��u�wc"�2˛�a��E��#tb��^�C?~���,��R��G4��izrJ��7�6$u��cω����ޥ�ܻFMHl�?xH�"�� ���������'�*������������I�i:[���-� u�R����:j����p����#��?����qKi艉����!����}/N�Ş�R9��j@���X�z��`U7Gn<��bC��DZ}I�l�a�b�h�;P!m��B�v���+j1i���Qt�mJ��@�$�W<4;/���q# �2��H�ep����^h�Z,��x�b
ҖIҩY�pD0$ ��u��D���FOO����]�'4�qؓ:X��f���R���!�#6���\� `��H�E=<�	�J ���H�����W	���d�B��p,�JݶJϱ�I�H��f��{W���ڔ z$�P�*B��ً�@G�0?`*x%�ۈB ��-����w��x���ȕK��������}q�x��Hr�.r-q���!GG�	⿂�1��k��:%,�b��֬��xtt�^}������k��A�h� ��n ����ʃ�t�ڧ\�N�P�Uֹ��.t��+��,�n+�L�]�y���MLL�ϠoiyIH^ ��#b�eU��ߑb	Pb� �*&9%��P��{n�JT�!�s�7C.\P����4��!2x��9.RK����қo�) ͤ�mB�b@(��x���ƀ5 B�-��/���>���!��T�Ͱ���e%u2!4E���q�� i�e�&ԣ,�V�Y:�0OזoJ�^�?�HŐ [ԋ��>��~�(�q||9D1�5�_@Թ��-Z���K�8w�6�@��͉�g��[F�Fi�1��]��-R�D������ϺŊ�Q@ƍ��*@(�0)�U
i)G�vf����d�u&v�{�3+�vW��=��C��r�Z)�X� ��C!�
i`(B&�+�
K�K`f�q�i諸�˧�|��|����UuuO�HD�����|��{�=�1�������d��+o��� p�n������"]d��d;��͏���#"�8�Ϝ�s�'��}afV���Qg�+�0��i�%Iq��)�a����#}��DX�[���k����Q��ce�V�.�#-�}l[���oEΝ������wV���[��걟������� �2�ڴH����#C��f��d0�=z�L�?��ע�o�o2<1I��q�� :�hWS*g�ޗ!̌?��=s)���uߐs�rXe��s�I\�Y~m�������� (f`��|60���ƽF�k�"����JY���h����o^~�^�i㛧���M	��х%v�*t��=z��A�\K�G�z{4��|��#��'����l���C�Ng+��n1l.Q�A'8��P�`A'm�U�.eD=���T�
�%ze\H��2K"'�������I�gn���䥤��U�3�n�a��I��H��Z���z��'�ؤ����J��|�T5��U�Tg㾾�.��>��鑔GB�c�N#2��G��T��Pe�0�Wi�\��@��Q���0��c(�c1�˴�j�O��-�Pi��[�z������B_e~V �An�]?��Lx6����ȳ�����օ�m�o'՝�D|Q���q�a��x��e$��R�&}�._G��_��F6~*� OߤT��Q�r�� ϑ����ls'C���F���(i�C�:�h攼��5׶��\=A�&��2ζ/�������B�DlS�?H�>�D��������{*} /D{+%�
�@Q*��i���AW��nT�;��Ugp	W 
��)$I`�D�?�V��q��;�{��`B�!��%; gs�]>�^�u)�1���FOY�sCzB�v�1#��?$"��A� ,�����1X4�R[�S.��X ��^{�.�3�fg���dޚ�&���;�;��� ~\���1ɤE�\�H6�4K�W
��7� �+��׿n�]�b@_ ���KY'��{���!S���y��BV��� X]o#�>��-�7J`�mt`Pzy_���(IŹo�eY�G��-#C.�c�Nzt�1Q�ǬU�t��Y:uw�n�l�N���G��Kӌ��ڦB>�c���`��Ʃs����[i�)u�ҽK��}�±0Fk!���Z`-�Ə���f����}sAe��Ǚ��43^�i��LѸgH�TbX~�Ļ\��"�w�ߤ:�Cs_�m��<�=�Q������w�w~L���F�^��}�7i�����b��ʋW�{3��k;�L_oԅQ����#.D�����K��<����n�OoD��ŭM�	J�d0�bMӘ�r�'��� `�2IOI���߽��I��C s�f��`�xlm��v���l_����#���hry��9�0l�K�#�����9�Ό�hf�� aly p��ţ��H�j=-���i�W��j��gv'}������:U�\$Z���-��P��]��a����)�D�
�`�K@�9�t!��>;�ww6�1J���eu���	�:tb�]����#�y�ZS�i� �=v���Ԏ�Zx��A�F�/2U ��E�V�6vw�7L"�[!��ɡ�������q^i-�L�!Q&8�c�7�J{��U�H�RDu�����q����t�)h�oq���spt�@A\�'t(�I�P��̾~¬8?�)�{��Ff%D���ut@�2�@)�$ҋ�>v�k�T����E	�-B
~� o�B~!R��,��@�����d� +}Jd!3D��M��O��+ ��h��D��©БI������s��4��y�,\5e��ĈR�2)H,��� �1��(��	���w�R�g(Z�DA6S�Y�ʒ��B:A�^$�atG=�l�)�A�8'�H�!�@ƔX2��z]�e�� S�XY<AdS���c3����<'5�����H�yëS�c0�?��J!hR��<E��h+�b
�:Ҽ/��a�u#�So�y �RJ�F) ;�]��·⻫rp>�F�J�^��*�q>&�}�(��)�z�j10����Wx�U�>�4e��,|^��z��Xʇ��ބ�X��Q��2D!h�~=#a��.�MRJ�?�b����s��Xl�ؖ,2ĕ�!b��\���x8�$�
�����#��2r�I n�3�%g��Q*z��i���� iž@�s�y�-;���U9��e*u�π��3�SD}�x�Y^^0��f,�K8�U��i�*�tf�]XA%�I��Qo���蹋����0� �}��2\[iǷae[14rDY�]�pD�^'�>���!��j8�
��ꢔT+ߖ�fy5@$; _u�e��_i�o��M�[S��m��z&��f�#�f��p�J����y/�,�͟H�<���m>�������Y^k;�>�f={�ݥ1*:�;��{wi��Q5�Rn��r$6&}){(�'<�o�/:y'��k�RF�*����N�C��[�g�: ;*��~��^II"�H������`�x���~��t?,YPx3�ީ?���ϒ!T�p_٨N\���d���^�ȶ�=����>G�p2)�a��I�a}��'2� �'nl�/��X>cA��(d�8��Je04FYtjw�����9������zvB�B�N�N�.]}`�L�	������>�������E��6�&�g(|=;Ĕ��DHjD䛝�l8&�+<!�AJܾN_@��+_�z���6�>]8�^�xY�!����&tdv�f �{� 7�����_��G;���?_���G)�0���]�!�]�����)_{i�,-5�2ڳ��(���:�F���z*����I��Ơ�_8p���=f�cQ�"��גq|0xX������:�y��8Ӛ�M�%5�T��Qd'ʢ�n�#L�H"(�4N`���Ȏ�h�%R:1pșd �a'�]H���o �8|�cЧ�x�XH("?��2�G�G�Q!�rZ�x��k������Oa���҉G�4W$N2'����B�ĳ=o�|��/>([�s�@@w��p�$��_Ni�煊��`��!5S���g��-%�VR�O1E�n���@�f0K�_u�"�{��b=�:��C^���	�� #�~��=���{xn�ʘGi̒�L�l�Q��hb�FI�QQꋒ�%�Ѐb �R!a}�c���'��%~}��` _�B�A��4[-�G*�j�������M.2��N�zR�	P(=�d@O�̫�C���d(��tCj����g8J��5:���j�j�2Jh��n+��ع�gD�o�AQ�@u��}������5eȰ�,�YNf�;])�����<���l��������Z�YGH� +-Ad�(=��̢�~ D���p������6 T|����9�菄��Edч鶢V��d��}9��0s�=�g%�?{^�{��F`cyq��В�̳� A+9�-Z��׉��<eG���A����~�F�w���3�:-����r��_0L%�nd�1��!9�A��1�ϼ=����7ۯ��d�|�3b�Ò�	�@��!i˴�,^$�A��\�4Li���ݍ5�'"��&�\�)�Y�^��jH���I�I�^�3kh-Ң!�J�x̶e|����v��ܙ�fO���ּց���^fɥlV�X��=ɯ��D��UY�d�!}~dZ��ǲ~^v�(O{&�A��G����7MY)��h8��������_mޙ����υH�fo��ς;:��(�k;�8��w	s���B�A�)�L&`��|�y5�`'��mQ��n8~mw�}N�C���ۧ�Ipr�'�X�r�!�C֛<HQ!����2��1���j�x�{@�L�g�6@�b�}o�.��M�&��J�^&v�L��ݠޣG��W^�;��oV�n�a<�H�e�dl\t;3F���Ov,a�$;��h7�е�w���ͯ~�.�l��k�PV���r60\	��� ��{h��;S���cp����
���Q�2:�-"V-�we�هx)Hg�|gy���o���0�g��c7����]�wF�Y,en5�D+��g���]d����y�����hz���)�C��Z����CC�V��BU	�dDAҍ�1�����d��ܞhz�T@"{d%�<�o, B�b{� Џ����j�I�J����Ch �KRB�,\,��'`(Q�H�̒hL��Z���:�TE�A�^�Y�qd�f츏G
K>�(��fy�KԬ#sVQ#����W����˪.�d>��[IY@l٫��_�Ta@��XD�ڌ������甮�{ĮG5�1!�-(���{�L���"~~P}��dV��K f����g�E���p �{�ՠ���W.�DG�,1�lR�������ۣ�΄����7�h��FIo(A��T�}l"����L ��A !�@S�EM2Q�X�H��k�H�ТG�F�`el��<# )��|��i:�|��V�v�v�\�ÿw�L9☜\�(wN`��`<ȅ��d3���6f��쬓�pY�Բl:��˗/K��� �@(���o U �o��y��b��e]�O��l-�K��v��V�Dʙ�����u�9�g�v!˃��HK�G�^�r(s�:���o�5�RN˼B�YH��l$�3Wg!AF�@��M4�R�^��jJ�&�Ӆ��TY��`ԅ����qE�pN&�����&��~e��;K|�����6���=�C(�a{ʐƘN&���1A;�B�X�VS�<t�KR��6hak�Փ�q`([�g�e�^�n0��/�	A�m^�S��@?�d4wc/��W�� �LQ��`hO����2s��륊��Tk�ר
��J"�M�8JX� $}����Fx6(f�X���P[�Q�}��ښ�>_G�j���#� k��S�"u�,��1�#\�l�7�|��?
	T(y.��Ŵ�W�L2"CH�y��Uh����ޘt~zz������걽���w���q�2L��a���* ��f|�%���9�:ϡ�&I�Yw��;���Q�mVj	}ζ��ns;]��ʸ��bm�}�����<
����.[��l���u��؊��A��Rifz��ij�����I�f�\���wzR�;�er%<��ͱ!�D�����^�^<~�^�L��Ξ�w_:*�ab^�C�<��8�<�+�@�l��h��4�io8�G�.y����w���u*g +e�w��^�SQw>t��\c;�v���s�\�|�fk~�3�����	����w���ɛ�������FO#X�D��M��ꓑ�`�
[Yp�Sɪ�-���Im��ܣ�/5�8�Yv��lhN/�6.j-;��(��AF�|�N� %h.�TgF`Y(���.�ă.],N`�`��Љ�&�[f��?�� �&S���j�$}\!J��=�~�z�2e�KH3 n����5Ϸ 0
���1#}q����p�� N�	EI��R���|;����I��@��Գi�)���ɬ����І�%+ ���'�],Kɶ��ȿ���dt�e����Kk�զ��t&��!�h�Mvd3�R���Jv)>�h�C��$[�x96�@W^x^�"�-�P�:C�0�?�:�_,@1� �Y5�7�P�Ѣ�/\�K�Oҵ۷����b#P�,����T��l�TF��X �]Ęwe� ����Y�`��"��hP9N� 	Y(���}��1�2�� � >���ͭ�LF�Nb�[$(�P����z�n�z���3��������E�@���M3npD�� PW
����+=� "^s6cZʆ�;E2B k���5d��D�Hҹ ��f���9����c�	�y�{��t@�/��0�Vhav��;Fk�(�]�����kmI_����$)�����|��p��弟�8�E�/S�� ��jkk?����?�gqn������_Φ>�߇�U�����������t��3�Ă6M(i4�J�Eq	�Tط��[Ox1z���e�J(��/�@.� 8X�� U<���ԫ���v�!2E�Ð�����	tw�wi����2��sdC��AK�q��hE�E���L)*���G?  �t�8�L$,���̉��b3a�Q}���A�O�vKl:ز�˲PZ���@�W���T)��4PB��ɄIє���98q\��ĜU���Ʒ��T5Y��)��pTJ��8��u��p��v�^��ʰ��Z�Yo�F��;���x�4�1"�,���]X#Y !L��`%�TYjs��=����2O��{:�j�za#}uu����n�>G���^��}��l6�E]�<u���>��<�v�:���,�ɮ��5]:	_�[��P_S(H5�qD)z��U� FT-�$bFJv����U��M�>����I�!?�����0Mx�'-���-4j��Q��Z��)�Bv����F�6G=R�������В��k�.=I�o.JI@�c�s�s'=!�S�F��[t �s���庅7�LB�7��eq?�O"�p�Lz%�~��4��#)�ZG
.����?FK|7�G@\�g�3�l�M�
����u
`ע~g�zۛ���]�v� m�F�goj5�l
a���IfNk<��Pu�>�1y�i4�^���Q�~^��Ɍ��(�"kc�eA$�6c��p�E��3�i�&�P��H�J�0|bH���֮���j^�P�D���'(��Hd0b{
V]����������1�/G�ɹ�dA,�	�����ȷJf��՞a�<�<��~�D#��q䱎dP��&����8 -|I
te�U�Ɗ
=�A���DJ���i�X|�9�����<��E����f�3R��>�!��hc[�HH�Rj/-0ЪҙS'E�����4מ��x@7��aa������y����^�u r�\_����a��*�K������9z��i���wi4�H�a$�E����1:uꔔZ®����L�,��޺#�D.$�-�1�W��S[�sWD� �_(!ņ���)�'�8 ������Φ@�db��i���4%�fYIq ̃`��+>?�km�3�~8 &6'R_&�yd�+�L��!g<�Rd�y�5ʦ����
�JQ���	�diI�.l&�E��T�����?4�c�G� F���b.���������瞆)y2���,��<(��=m�PN�5��G� �Xxf�����}��{�Wܲ����m����#;�����x�3����?ַ*�c���ޓ�\ v�^�{�;pu��O�٢w���ٖV������Q��s�kG��c�* �o�ⵇ���]gW�)
^GK��f���t���j-$l�ȳ�W�j��5J��x�j�_r��磱S1���$PVFN�@ c��u���O烪�=��a�E@�� ��[bK�;�b 8�>0Z#��-T�h	LVf�4 �WU729�y�B��At�"k�������=IT/��蔠��|�v�=Js�$mB�!�gAE/n�����n�^�띷���>�+)}���׉������;��|7�1ߧH�}y~9��}ӂ���Ǚ��Ȕ���d+S�&:[���Kz+�9�߿���ݽ��cJ�KJ�Kl\��:��DƋQ�#�)�s�6�>+q���
��)��2�y��#�����7�[mj7�S����^���v������H�3����NG9.�8-��ѐ~�v�6�	���Vg���x�.���ݭ-�{���,6�i�٦a��pOh�'^B�Μ�lgLWw֨C3�����<�<qǗ'A"�$)9�G�A8�%{�9��n��͖����\������/*�>�b٪{�|��A��i9�0T�=aK E�м�����B� ��;}�j;p%��=�{1�����OǗ�hif��DA]����9�������0J�ʓ<H�pv$2	Q�v���Z�l��D��x��x��PBȨ�cl0���dM$����R��'i�.%.�����0x+�-0B��w$��^l`��;�%�&�`�x���0�"���%M��߷�W��oH�i����$�`���.��[?��r��'/�K$�'Q�=��\��������m�/V���8HD�|!��by�oq_^���Al�A�)����{M�K�O C�$��õ4����X�۠͠K�LU1�EeA,�e���08񽊔�H���?��* ��6�/ �q�W�s�y.B �ϣQc�ߖg��Wf��d���+��Wy?����Q��L�bQ��	�6��+s��^�R�A�(�z!Kw�M<�ql� ��{\�w_�?2Z;h�/ь+�4�oU�;���R�}�.��W]� `�߇ߎ��m��M�;�* Q��P�\����@"���Ν�cǎ�+{ue�8��?��k�G�`��=̆�Ke���Z���%�����@-�2�2hUjl�GF�,��h�a}@���T|3�V �<��xڙ�	�ᾗ��|�"�~%�C-}M8a[���L����}ί�c�CvF�r�a�!�_r�BDW?_,U�f�}�ɵ�k�w���x"�w��\_Sj�tzl���ϿC�g�������*��S4��~�=��ϼd?)��q@�0>�x�_�?/6�3���j�;,��~���=���Qo�6z;ԍC�2¼�J1@��|���b�I��U��:�V�I��]ȲJF��Sצ}@��h����2�JY��b��f��@��@:�ңI��3�{X=��OA�d.2#%��h3B_=�*��T ��š5���2YP��)��HJ̧61��oU@^<J�SadK�!�P��*ϭ	7�ScG*8b��[� ��D[��YJ����P��͘*�] ��j8b�S�8<����O׽ڽ�GpU��^P�PP�k�G��~4��N2�F'�ا��b��s,��SR�_֧i����:F�^Ij���f2zi-|�~��?���lo�����Z~0�|�ݤ��C묹~(�KA�uj���6BO_8�����)W�l�����A��A�F1��@�;�p�'=��@ۥ�������G��Oh�oҿ����$�����K�/ѥs��;7���#b�'=�ܺN��N�.�D�(��^�K�.\�Dǎ,�&��;�y��7_��Mz룟Qo�#�T/_x^�?�X�G�"vn�2�.Jj�]��¿*�Ѧs3A��+�a�,�6[�f;N���w�^�������ϲ7�����t��.�p ���c �Ad7�U��\��dzA"!x8`s�������w�^m���'�ԉ�F'���xNF�[��\�S!1�����8�<�z&Q@Ô�N:����mڽy�N%�>א2����s��;+<�Q�Vf�>�$�h{�K�bR�nJ�]S>Wl����C*7�T�6*f�7�6ʀ�,�%���I�%,��pBo�>MFc)�e里P��GZ�ܠ���-��w�xr��,���c�vc��my�	S�/��K���"��2��{RN�EZ���ZUJ^�Ͱ
�g�5��"�M�O�l�7v��No�z|ܐ�]n6����%���Ȝ��9����˗���/���e~�uq���Ai^�Z�T�A�4�0c�M�oP���P~,�����Μ�����m$s�TI�LblK��|�l9���e2ٙh&�xU���'�?�h`�o,��7�?�A|3�� ` "B!�T"���l��w,���e�2�Y\l��k�)hnm&�e�,�(}�������FC�9�s���(��*�ƈ��[���[�����#�C����@����"5q��5��w�#�2�\�2����0�N��~���#e�Ua��Y�c#+��l".EF�C���K��_���ȫ�؜�Fm��jz��yښ�P����pG�*O���j��?汃�f�f�(�$k!�?��x=��J5C��)�ڡg(��d22�N��Ӏ�b���v@ͮ��\?���}��Pv�g8��b��<��)�p[�����ό��n�~|�Os����c?	,z�i7`�v��E��L��Q��ЋGOә��B��h��C�mz������y����s�A��?J3`�S�C����v��o*��	B4 �$H�V*�͘��)Q��f�\� �=�n%4��2�3��h@_y2�P��Q�?ɥ]���v���G!5���Y�Sˋ҇I�����0���� �H��&��%[:FՐ��i��GնO���Ī3b+�>-���!|�G�:�a������ʁ^SI�SSk:�g�������'��Ca�Q�� 5l����0�W�:y��뿬=���ؿ�����U��ƃ�����A�6���{�C�# f�̺)��S�#כeJ��L9�	��c.�U���C��N29sw��ݥG���~N����jX�?쾼O��/�KPLJ�io�]z%�^ �b��Vާ�3���}p�o�������"qQg��r�F؋x�A;�0X
b���Z�{�����+������1;��6����O�@��<�U^�'�w������_�7��%���D�y4أ��ߤ�hHq˓t?z������_�!;P�H�u���=z��G� �Ѹ�@�qa'9&��2�KHS��Lq����M���}vy��k���۞?3�~��0�jzj p��T�':d��l���Z{r�s��)Z��%�W5���;ʾ-7�[:F�NWj����x!E����GT�}3K	��!c���0��~N��+Ԭ�ӈ�7褗q�2�y�͊͋�,u��{%�d�Ǫ𘩰C8
H���n��)�Q���Zj� F���#�:R��PEJB4�5Keq^S`�������������V<��$���h4$`����=OJOe��祦��fS4I�4pB���i�E����ɴC(!���H���̜<�$L�e,6%ߔ�Y�B���B(������
����X<�@��J?ʀ������>���ȉt��q��[0%{|��L[�FW���7d'�5�m����K��u�zr/�d[�F�����8��qG�"�ۘ�{7��I�Hj#�4)!n1e�Ij�PN,�}Ψ���&�������h~v�N_�/�H ���͢��czo4��a�� d!�Wd�+�\�L!�p]�&����˂���Ҵ|�1W:
����}�N���闿�%�5�i֥�3�X��
�1����ޡ���n�o$Jl ���wߕc�}�H D W�[[BZ#�	�����xf��q�]~�ya�{��眑VZQgS�j ��k�r�)YEe"��4̡����|��4;I��d�����'�E1?�r�3��2��	6
��/�@�+�dTdA����SU���8�<ݪ����s��l�;��O���'�I����OM��
 p(�`� ��l�W�ݟz;�L�e�0\���v|��>=(�â�s.���'1ݿ�F��v4G���4�n҅�#t��
����`L�{۴�ݢ��#>���j@��0J����0|�l����P�J|�Fb������M��;%��"��l�O�6�ђ7��L������|����y���ߐJ�Q8�����T�u��K�6}��k����E	0�,���:�s�]_�/���#����ڥ�Dc9 /�&���}������)j���]>A/��D������z��#ie6u��#�6�TZX�d/���Jd�e�~{ M����C2L�]�mw�a�JZ��&��K6W�Z�U��y}<^���{�׶�Q<W�ﾲ��W[q�kzRߣ�z�)Ȧ-�j�s������W�ͨi��l2s��*dmٻ�7�|����~�[[��O�\������n�w>��(�~�K���K?Uj�Q�^����1���\���&W.���<C�p�Dl�����ザ�@&�o#�<���]�Vig<���B�FJ̴��~�g?�Ms/\�,�Bp\w����5�p{��J	M���V���~�v]��/��Z�6x���{����Cw��h�C %H�{�E��Kt�'���Q�p��n�G�ѝ��+��,�d���F[�eF^A.�f�f�����۟!<���f9/!��g���>U̵g�]�݁� �q�����E6 ��G��IvL��#c)3�%�6�ӚY�>2dw D�>���'D;f�z�����#�4�}��� �r�	IJ�xg8#��B�@\�ق{c3iWR==dyz;��"s 2ɒ��j{�"54���dc7b��(S�.��u��{�ɆJ��2ef���5�`M��B�!��l?��{0�3�M�{؁���� 3���0,�g��-W	bB�r�h�I�EƁd�*U^�ȶ�x�j�3 �D�U���V]����ו�3q2(h��[����R�s/	h�F8�0��O��j�Xf�	���e|��_�����+��+�m|jsU�0VFYD�7oKƫ���|F�'B��Ǳq��&���K�b�m���Y"ur���F⮺�Wa)�L�jbfz�E#�,�蔉�JE�7'2'l�?���rVQ������d�\O�c�,�V������j�:�Ȁ"d�A����\O��������t��E �[��uZ�{��1�}�d&�ܾM����D ��s�iyeE�5�`��x����З���}C�D�����Ŀ�5={�l����fs�z�،*eY�L�n&l?�qI=S^�lɱ��f��E4�()UiD�؋�;�9$i���,�,��}�@�'��)��gf�Dy4@2t_��òA&% �3�0��~��3�$�&l?xޏ-�Tg��9f���0��fx����p��;����O�ƛ�f]��l����4���Z]�"��������T�����f��1��4���=|D��65ff�>7K�:5�hڮ��y^#P��6�,��\�v���"3L� �=����q%���+ޔ�@a�������Yar�5��v0�zVOM[%$c�s�NK����_���]۸E�3��|�ʉ"^����苧/�hc���Q^�m�ʩ_�:�0�uz��s�K������pg�T���0���\�7._��ݢ���U���cg�ϿBG؇���ŦT5��z��㱩��}K�AW�H�L�'�Iع���0ǻ
��}��d�!j���4��_)��"Va���[޹Q�@��x������ZG����6�q<l��\����b;~c#�R!��+�).��n�(���-U�Ӟ6d���u�I���6��-
����w�����T[��5�_�����_}po����m|{�gGt�e��V1�<3X� ��y�Ծ^ܟ�������3�h�����[�LJ�
&�NcaD�����wi�FI膑9�c���޹C�l<~x��Q�^�>;�k���A�N6�	��x����tc{�Zڗ2�{�����Hŷ���r���عGJ�TٺKG��Hdh�������4ã��)Y�]{&� �,;��>I��X��&sV���LG,��}[� ̄x~��{�~O��ŧ��_�$D�yJJ��Cw/���O��q/����Y�V�%ٮ12<�_��m6a���y>��د��C������<��u�]��ߢ�A�zM�z*�@�b�)mvv������ߙh���l�y1U�:?/6f5%%���:��߯J˧E����8�(5Tu�n�:Z��H�:��LJ$��z�FY"QGd�t�)�x_��3x�*�MX����S�Dc��Z�� �
M%� �TM�`�Ă*��~9�Ӝ�r�:������ӱ�c���AG�Y�A�(�AϠt���G{��lm�<':�ȹ(Ì��~�<6h�. �*Z0*t2�[���e"2�_�1������_�l�
�S�O�b�l Y2�l�ݿO�����>���Z3:}��$�GrBG�Hvഐ�O��f6���03����<�Jӧ�} TP�\�=���-W�t��q�a'v��L���Fy$@�^�Ǡl����~;�K�X:�<�=�א	s�� T��ZX�-���8Ο�ɟHy'@���Z%s���3�issSX�`��._����@wE���$����#��@�-JG�[{��=�����`?����@���\���ÿ���Ɣ��K�B<3̇&3��X����u��a��qF[ۏ�7�Q�hA^�'����C��]-#0/dC(��-���(<K!��̏0�*#Ar���:�Y�࡛+?����`Y�>'���8�!���%�v�)���\��0�����	�~�m_��qmE�W������ˇ��Ձ�-�_q�� 
?홚��W2�i%���D�Z��(�Y�=��56��6���� ��F�Ӑ}B0sC[�@t�mG�l�<����y�a���F�TWǴ����Vd؛Q��>z�V`eV�d�(cG�{��9�Z@u�"v>�,���Dc��Vg�������}��������S��ߠ.�9�F�I�k��A�����+/�L�HS;���K����/�|m��\�J����<w��t������Uj���\���Fl�k��ȯ��9�TVw�m��H��6�<"ӂ�F��(�C��؏`0��b�'4ď��h�=��������ն&�W_>{�ϼj�-��GI����m�1�~0ZY�o��x�?�J�_�h@p�3$wR�%��8���̵�� ������j�I���4N._>;3u���k���uSyk���z�q�tE���޺�`���ïlŽ����G*���J�D+�ll΁<:N������2��r�S\'��5Dv�n:X�'@��ϓ�?�6Ɋ/����D�tdg6�1u:#��n�WiTJe��/θ�vcz?����#��3�C��9B�?6��O��`&���{d'���vKi�g�d���H��K2c$�sdj
�l *��y����.K�"���r������9V�a�B�����������K��2(�[W�<OU���^7��_���` �c���]�}��{�ZX9Jv	��d�
�!;�&67��ݟ���R�
��}D�^H�U�"�q�ݗr>Ld�#Zh�{jJ��m�x��y��> T���@��0�&@�0�,��PN�!���|��PդLtȆ�9��4��D!$C(��P�!�ŗ�h$ȟ���ƃԫ�d|�� fp㗪R�P)�FS��S�*ɂ����0 ��e;�hZJ��	?d�t(����T��{{����1\1�0N���O�	�GʠfvnV�u�^��%yfR&���%�����'��G�L�(�����4�QL�&���W�iO!.���90��<���}_�^�������햑|��|����Ls<t'`.ՙɈaΦn��'�� W~IʁEZ!5l�c(�]
�I&Yd�p ���e�,��Z��d���<OY)�,��9�'��z�yH~�?'�I	gI����Wb� #��1��c) �dbb� ��/�`<�����a���đ\����sE�1�K�����+SE6�ȑ#��w�}�S��V��te����4�ǘQ�$��"#J�ֱ��!��I)B�A0a�z���^� ��w<� M��ԯ
�m�5��>�4��,!��̤���!0���`�\�ěy�:<E��"4?S&���n���v�{�i}̊���~����XD91�A`Q��`�r%?��/�_��i��i�'�w0�����Iš�hlϤ������=B/�A������!��@Xm�C2���MRÊ��l��L�*�oJ�e�M%X/�� �b@�f���ØiO�]�G�V��4��АZ�lE�X�m����0���J�����ӷ�?����rkV�eO��5K#kڞ��lkHLx�g�Z�x-d��47G;��w�u�����Gwo��/�"�O^��Փ�\�9  ��IDAT�d{��ܿK�kkR�&���Kta�(�f��t{����ˢ�=i����"��t��·���H(���$�7��R^���W����;"�v��:��H��\�:{��?z�^y�%����߽���v����͵�{��S�Ƕ����ߺ���%��O3~p�W�;j�ocog�LN?����f�����+%�{iH}h`7*9�3��4����2���Dv��:�/�?j�F�^tЪu
���P�|s��VRj��Y{��??�����O���[����åk��7L�r/�>.�5�}4��i���g֙�R�2}����.d
?p�@1�@2�ʮ�DrK���l� ���p��]��BF���+J>�Z@�l�Fk�)��y�x�d��x�P��d5�Ȉ���I慍A�,	�F�2];������>� ͸U�+���fD4���)���b��A��	]��>������pmՄ�jh��,Y�'8���ez�ږ>x�������s0����-Ot��̕T(Y�*>�gd#�ݧ�W�r���a���Cҫ���o��H"���ҽ�tk�G��c������7 �_��� 1�:�����W����B%C��4=�+����"9��Q�0��I�A k�!�T&�Y��E>g�-D��g���2L��*6�(�Ŝ)�1�̪TFW}�S�aa��A�R��w��8�T�T�g����D<kF�#]pfT���8�q�R)�k�3{ Zx�T�rǶ����#p���)�3sQJ\Q�++�`J�	�*F���9��8/�Ɍ��{�,,�l��N pC��L�)�pЧ�� !|/���('���۞i���:M�)�Ĺ���f\��5�4Ԯ5hoҷ��7v ׈�O3���ɸ[�e�C�%��T0������lp4 �a��pTF[��]�E1C� ����t�Ϯ\1e�]fЁ7�o��c�3��������}x�#����!KX��X<P���%���B��#����ӫ��&젆I�*�N����ׯ�g1�Я��Q���5����#�	�C�i�]�ȴJ��l��B����6��������Jh��fMPGk�#���m$,�e�!h"%�1�'��	B���ʶ��� �͔{%C�dN절��Wr�_����e4��ǲ�v�K����s$.�o�m�-������������3��=U�PNh�,�?����m�~�'�oo���q
� J9��-�D�fo˯�fL�D��J��Ϲ����c+��n���l�m�
��=��(a�fj��x����<|+�� ��Ч%�g<'!�BX��B�8��˒�)#��+*Ez�"�@��p�P��c��)ms����Svj��`M��ۣG;�� �6�C�.-����	��<�ϐ�f�XJ`��`ЦJ	~C��H��V�Y6r)�Dk�	�b觯�ƶ�"����,�f��������{U:�>ɑJ�N�,ʱQy:�xL<���\�I�[7Ae>'��tl�M6�m�B����c'i�,�ŭ��tla��k-�}�����x�EZY>F77�)Oh�%��KO$�:2~t����҉���p������>�GW���#����
ߍ#�7{�>�v��|�����n�Vg2�����n6:7*S#��	V�	��d������y`y����2��ͽM�w��b�!�C�� ���&���%���,�{��R��Th�f��_d�����������]	�P��ͼ�`������|gg��ο�y�qٟ����63h1"W�h~�b*�@Q.��aW8�r���@�};<����-˘��.���)�d ��?���=�;���3vY]e��� ��b"˾�}S��Bd��������V{<����S̥�%��!��U�pS�9�!]8��Bpѧط�)�$��m�L$L��q] �%����L>."z���xE���6וQ��� �8؉%�i�/���<�,����9�d�Js�'jv�AGWfics����&�?ڢ9�@S��0<�Rq=)1F)X�Z�/�;e*gsj{��=�F�ΰEF(ϋd�����4�f%4���ec��fE*b0��{����*�VBi�U��:�Jأ1��D<}�ٱ!�䗵T��!mW�����%��N|6&�(�$�dN�P'[�x=�0���AO� �ɋF�;8�(!���J&�*���%/. �y�'�c�!��0e����ӆtE�����@0�<�_mؼL3����≞��P�Z*Θ�O�ùS���ϰ�hYJo@��W��A�I��(����#������ջwp�C���l�p���^�5�,nD�E�@yyP �尛(��yx��c�d��`�kD�C�c��	��>S�2���,�^�4V�C"b�������p��x/��>C�/�Y��d�\��pZgP��H������k ��P�y��9���I
��>|XE�L ���?��?���������ߥ�_]��� �{d�Ć�q�/
���� ��w�Qw}n|:�}vJ�'���uJ�]���.	 B4\�Pȫ{ �vJ���R��_�#��JC�gQ���A�k�]S��KvPK�Ы��n�%K/��mX���Fo��NR�P�`�zf�ɷB��2�k�;�o.`H��XM ]hAxZO��K9Yt^ |d3�N_Аvh���-?�n-t~�W�*1A꼽DJ�܊�NDO�}
8R�ǃ���}X�үՖ9)�2(gmU�y��ٚ@�8-]�ҏ��%�'�?s���K�͍i�mA��r�ۅ���"�!�Ȍ� ��&�
)�Z�"�d%�A��� B�� X�W���	��i�H��'ԨՅ]��h�	�M�W�w���Ѷ���+�~&j����������� l`2�h?@�-�8(�z�v�Gv�B�"c����ϗZ���̀��oCU��3����X߯2�m^����u����T�WE�L���Vؖ�\�����.�����ٺ��|�A���E���/�Gwo�.��fyMb_���;ԃ�У;З_~�N��n\��k��$����h��s^�����Uz��U��>���[�^�	�˝۽��X�}}�ּ���^�����j�Tߋ'Y\����7�I�B��_NUZ�H�'Y���'�����dpe/�0Q�������DاS��+Q���������t���b�� zS�Sdi,dI}+ߤ�K`-U�ο�°��ti<~������fOR�����Q8l\�Z=����'k��ww��~6;�4��2Q���F��`���k�>�5em=��t�G��@���g�3��|�4�: �bN��t �ک�|i�r ��" ı� ���W&k��ϑ�2��RҦ\���v��x�\C>B��*q�.sM���#���g���?'�^a�*���qsvG-�Pb�@(���_����Q�Oo�>0���[�����ת�ĉ�@$����\�.^�Dg�K��F��K��+�.�MB��l�Z5:vr���9Ez�*��H@��@�Ͱ��5O�1���DY#KF���'��}<w�p�1��(AIMFz>�<����;��R]�ɡ�� ��si8t���h�G"��=r�A�S)��P�
C}��~Jm~��3"������)�xu�b��3�?�8��?�,M!2�ʑ�C����0mia��.�$��DR2a��2�%�G9 �r�f+�[z}^���Z@�"R ����hU�]ی���R�	0ȋ0�8!^~��>Ea ��f`?.�e�\�q�'�8�ϝ���6��ۨ��`�H�`�*/��.��77��͋a�C�D�	����r�fAbP�HO�[�>��X���#+Bҳ�7��!���d%�J���R�/W��s=���6c("���^Ȳ���� <�c�߮���#"Ӌ�%4�%��+o!� -�@Us��두̠��?�9}�ߤ7�|��޽+���RS�7�����������H�R�H��#���Wp���,�S�P�
� �Ȃx6���H�����ҫt�7I3 ��3�S�\��5�IJnG}~�#�whg{��<F�>ʎ1vc����6�b*mLzA�ˬ%�$���Ȯ���쳲��+��M�����<3�����}֌-%���s0�fm��|
2ʁ�޿{��r���F��`�'2;y�HME�E6yf��=ΧݞT��k	�&?p8t��8�?��>�g�[�0X�o�aO��$_E��PH[G�}�'@2.�̫R�f�����
_�8���R?h7�S�X+�R-z�r��/�A����n����u���1�Ղ��I��s.-,H�tb�`���ҳFC����%��V	2kJ��('\��Kx�� �:Z�m�;�i�"�7��7q��T�
�~�b�CQ&�G�Y��&�C䒐�B���[T�E��� �{u�!�}���	Q��WO_��LKh)BVo�����6�=qJ�� �|�=OM���J�޸�E�� y4�{P��	Y����޻G�IJ/��Hͅ�~�J?��=�+�ݓ����f�(�g��v�Ag�Bg�s�G[�iVj�M���P�ݹz�Ӭ�Gl�*Q�����$�'��D'�J�c��M(��T�x����>dک�)�����XGUl��?;�����[�?��}Sf��c��Bn���.��
P�ws3�����?P��H��� �͟���W��/-^�L��!��(��n�8���y�~g�������*�4*Ss��j�<V�L+��&3�.�E�\�N �6wjK���)�>�� ����`d4%��Ss���o���K�����v祖��DyS���;�s�N���3��f1���z�̐�h��.�6D!D)t����ltJdG����/W���{B����I7����5`p[[�z�[�ۂZ���L� r�g� �͓���}p_7�d�dy���畁��7DB
ƪ57#3�a�4a�c!� ��A t��0��}��P�8KG�c:ɛo	��gSa#l0���͆33�@��J��R2����n��i̷g�!o�ӈ�6��J CJBM�F��5^l�Cd�"��Dzt�!����5ؚ�R4�f���i>�*JK:�r����ߦ��m���/�]_�J}^��A?Rq��(��BWƋ烲�b����yRV�V$�
��>/
eD�^h�$���[sGiĶ�=���|'�\"vP����ͷ�f��s����}:J��Z'�h�d�΄�e��D#���A@��M����g*%%� .z0be�>t��� I����o�ZYY��<��F����Egs�a2�LI&��ۛVh~��G=���ݼ��K1m�K2�����L԰�lL�4�T��*:	SVY�ٹ��E�g�`z�d�,5Mr!x�SG���I�?���s����	���ۊ̰�lf�c�:x?D���9��"�������џ�{��^0��F9)��8/d�� L2�� �Ȩ��,�&RnS�X��9	�T/�y,��B��eȸ�HB��m�َ�_{����LY� ����v?�;���|�v�y����⿗�|7��x������fț�ɘg����ևOۤc?�[*����1�RQ�e6
,�(��sl�3�D�n��"9���b��Fk���V� p!�(�$���S4)�#��?q���`P�O~ϮU��ˁ��>�|.7q<
|?�r"�b�M���O�-E@3_���ߔ&�������eh�Ґ;5��P֯����������A@u�@�r(���4gx�B��n2"5˸G�� 0��4��ue�����3!��Y�����1� �;� \��MU93!�!	��ۡa��f���/���+s��{^�kTA�J��R�ʡ��]�!� ��l_��X<G	/���_��RM�h �y��MZh�h��D^C ʎ�=�-+�4��Zu�Y_���\��]�
8��^8q��W�y(��2�Hli�d.�̘�:JuEM�+����/�k����T��~�->�m
�����iva^�g����%������]a�o�ׯ�?���-��C	�bl�56βٞ7ѝ$�Ǯ�zZI*����(ϏJ~���2�t��x�^D�+*����LB> �kQ5R����3��IO��.�Z c�	�3`�]T�ɼ�D�AB�1��	{��4�g���������^|�j?�����_�]ZX�j,FJ=��k�v�o�pҙ����>�ۺ|;���8K^�f���*����h��8��4�yf��-���MA����}L�4}�Q8[���eA�_�����D{��D�,�ؙ�Y@�K�"�中��]��]O� �HJ��4{�c�v����ep:z��0�eC�=/�<h>��MR�T�i��[��O���e�jj�����U�4��oZ�l��k�L�Y̠ŗZU��a��f	���}m�c>������-��(р�No���kg �@'�aJ�W$�����ف����C����@&o*Y&�4*�ҧ��šq8\�P[�Tm�s͏G�H(-�(�f	5�(ɠ�d4B�Hz}��W�X��1�� �ῷ6@l�j�M6�sT�F��qt�:`Ј�kW*�۱�hO1N�KF����K_�*�[�߫�#���o���6R��oid QFSmP��A0����~��y��g�U`Md� �PL��J���S?�N)댩?��	Q?���Hgv@�DB���:Gd�p�H���b �����A�'@>��L���k$�5D��:���<�����Mvz2F����D��?�c|(��B$�닧N��+�����;��ع����:�p�族QUJ�|l��T���ܦ��_�����b<�S|L�?�������:�/�����16;�@lpLt�xM�ܫ�)�L�<Sv�-8J�� �>�O����jG���9';��c���Q�b�Y�>s����o��G�?�!]�zU�=BG~�� ��Q�AdAD ���c�ҥK��s��w�<�N�Ź9��[�f,�T���}�[�m�utL�ʢĉ�{ʇ1�ELF�`o���$C���� v��MG�(e���ӡ }�<�bv�tZ��a�,�4���|&g�6]<�]ð��d{O�8��{2��2�%��dOz�4��0c���>�����'���T%�=P�i�q�3�]�̳�s0/��9�̮����_�ݲ�}Ƚ7��ޛ���S�i%�m�Ml	y�P-u  ͗�["$Z�'���+������g������*Jxt�
�Շ��������ě�q��y5�/62O�z�cL�aO]qM&�V0mN覎$s�g�4�u^_���tf��0P�����TfD֪=�9�"�,��Y0�f��n�DH3�!`�@�WM$'pu��I@G�Q�F���Q)���6J���+'%؍������y�3���6iE�Х#'��lkңZ�N/?� 3���ǻ�5*�FO|i�A!�P	$�t*A]>��,rYh��9BF�&�G+�DV���z~�4���{�n�jw���-���Tj7��=�6���Kt��9��ۥ��ma��W)�΀ ���������<Zn�ɹ%�_{�����_JY��j�:���e�t�:����
�%4}�w )���P�>�*^Zf6hm<ce3{𙽂��9 �K�\���v1�\�"�����a!���l^O��5����~F+�4�J��Ѱ���Voݛ��~��G;�r5l7q�ZOZ�F�0D���]�{�~�ޣ�����/.�/��2��;*|-PYc�����*�t�懟IOL�:��}>�tQOr��ڗ1�l�D��{ r4���)R,�7� �M0�{����e�\�&�]��GMk����-1��Q�S�����9[+�`JY�DC0�w~6r����wj;>\i�s��[M�
��埢��ޝ�gA!�m���Ӆ0���H�/��HIl�LŴpk|>S���:�BDY�hp�-T8�.;���.�M=�'l�Q�� ��b�@���ȴ��tdzw�������ɨHJC�g�dی�P��v��63̧e�@ی@���=l�����@�*d �&�PJ7�l�]�&C6NlL��d#4�@m�CYPx]�LQ��]C�}�Q&��:����8���)[��!�F�?E->�f��`2�ȕ޴���R���B$YYO��H�Q�2�#;�iC�� %���L1[�Hi�Ǹ�!-6d�'m"U�(�qJlOi���[��51xg�V9ar�B!F��|H�zl�dS�M���ސ	�d��ύ��`ɒēPX����l�$BޯZ5�O�����ٳ�0VQ҈������{�&K�#M�#⮹g֎
A $R$�[���e$k��~�O����d�-2�~���$�L��-kɺ)�9l�lp'P�
U�5���7�ȿ��#"Ev�#ꒉ�ʼ7��������CfU�g��UP�8���zK~���%�1��+\ R1�!��?�砅ΦϲV�-	�� � P�3��@�{�ǯ3y���4�Y��ǫLU�(��x�z����������
��[z�s]�Cn�#]wh��� �����1��c��s�E��͛7y~���`����l�TE[ �1����
�$)lq���eSY�����T��d�¬�Pm(�^�(���+�~N�~x,G�w����U��O��x��Q�
�\)���ܯC����,oE�Z_�_��<�$�}�j¢V��5��}^T�d�NH`n*�I��  ��؍��5�Ҳ�\��@��ǿ-�C���W璲kg��s�`����ت�}☜�i{�~;�k�$���{�Xf�4j�G��^F�~���;�VI�)��(� ��y �:;��_Ufl���M,!�-X�6}����㑼�w(��)�7��4[��yF��z���`_��hwP����1��C|���hzJ��kǙ�*�Q[�
\Ύ�u����+���tN���V�We4�}H��S�ݐ�{2�=�����������Llr�.Wլ!���D�T��>�W^}�"p�%_z�u���/�|A����*�z���+�d�\�j'�Wzt���;���Y��z��
�.ȩ�c����r��m
��k�>��v�����Y��g�,��7�n ��oO���3��Ί ��fu9t��X۹"�|���U`�����We}{K��1�!2��g��w߻)?�������fy��W�Ͼ��r����m�/�i.������E�C�7亂���H~���r{��V<��a�-e�Ed��1W~=ߗ���8hϼ%�6|Ah(��38��S�Z������HBLK�!�~ �:S�?�Ba����O��=���a����Rn��bSA�G����*Н��}�l�~G�q7+&�}��[�B��х������Y�g��h9}���?3+ʭE7��R�t��O+��z���Fա�_p@��f�����W�D�64R�?�45(@��[��e8�e��o3��q�\h՗tNl�����⺲�yBѴt���g�p�:�ɨ�8 K�p�����YK���� �P���5vY����f��( i��֓�9�p���=Er:N9��jn=��)�F��1;.�_���c��35�p<o�\q��C���k�*�^1��|���-'
�N���e��@��+`ʦ:��!4G����675��@S����3���+.M�L׊�\Ǣ`��ӿ�A�`���j��� ֓�Id�X�1���[d}m��+*7��t�=ecu[�IHu�~�Ѝem��`�@�g� ]�^��$o��G��>B\�z�w��Y�J��<[v�q�~p����WĠ��:�!��6��������ԩ�� ���Ŧ
` P������ Hjލ5��iab$&^ٙ��m���YZ��tS��fF�9=>a}&��t<�g�3��{���{�a�s����e-�	0��"4�bf����/_R ����=�'� �B��� ��)���B��g_d�<�n��{D𲹿%׮^��*O(��5����{�PSC�MU\�O�&We݇�pQ%kS�6�N|c#��{xZz� 0�Zfv��|�O���������6`CV���o�l��(h�����9vv.�"
z*���ܗ/~��A�1 N��ϰOD�g�|��������<Er<����f�f���|������2�o�g6Խ�qF��t:X�kv$��L���<�m}����5�����C�Ƿޔ������ly��l�*�%�����
k>��J0� �?�@�}Qu$0�̎��S�-��! �S-&q��+2}߳2몁�J��<�����7��~6�zL�L���d`�̬��Ѥ:��A�Kp��:-��-.�[UM�������(m�s;�Pa8n����7cMi���<�{�����S �vۘ�V�ݰ��y�Us>���?=h̦gm�	��':�.��woɯN�A��X����� ��'9�T���j� /���a�B4��@��(�*�>@�d�4z���zo��Yȣ�{�hoSv���]X��٩l^ؑ����|�7���T>��#2T�Nʝ����81�
? 4n�X��7�Vç��tuo�܂O�!��9�=�駮��繬��{z����w~.�W^�-��%�c��'���w�Cݓ�r���W��ɪ|����)��N�o������ʤ�Iҁy��Ó�2_�91��2�C��Ὗ�;�ޓû���9=�1�������,��p����x��r&{w?a��GO]�;;���?����=ɏ�]�P#�wz$����C)���������ܭ꽣���`H�9?�����r���'ܒ�\�����}�B���d!�Y��������J����w§�g�d��A�j�#������,J��_�g.v�2ꞹsԶ�Aq�zB���"�]���zN"8(3�ibBN�zN�jkTf��<����:�3uK��K����}����2/�92�i*�Ӭ�-�;˪�aP�S��7�g�\8�q��:�>�Q(b�[�d���j�"MMa���C橺���c���Bģ*9�@�
�	FV� -��N�ҜϬ[X/:�8gp�X����gF������2�Jj6gW����DǢ�`.	�r㯶���57�63f��P����|����'(@��+*�q�tL̎7���Iv��
�t����Q��c,��θ���=  ���r���,����u����S����5V��	��Auė�.�S�ϸ�
� ;�`�݅�Ϊ7�Nu~j���-0�*��q�c0� ��ܠad ����@;j�lJ��x���f=��:�tr �x/P�������?��C]���
oW��5.����Ž8�߯Rf���
,D��,z���RAj*�J,���r*�~��܍g�/�� z&?|��׳RrR��
|�w���(u�"��Be3 �����YDn� �Ȏ�}!�Q8ʐ,٫��?������w���]�|XgPV�vp��4��/=�\�uL�����s��.������&����9@H�Ɲۥ~6�7rN@�����#ރ,ha�O�R������C�;/��Y��m��D����˖�顖u�z����q������6���
��� �6�)�b����v����ye]�VS�˒E-a�ʤȸ4�g aa��XC#��ãC:p��8>K���zA}��X�BV�>��=�W̤��~�=x��u�/�����o|����D�0�/d�8@F���`�$�M]R\���X�`�I�v�U'�yT��^p�.��y���G�J�N�9���a�iU��֮ړw�6�_G�##�w��V�\N)�~zv̟s�8i������}e�֬��6�&q�Z������|?�-2(�1�"�t�+g�;��������7�ǿ�Zh]h�h"&n�� 
�)���yy�0��̢xc���Z�!q����O~����.?X"�����O~Y0����f����q�/�� 
qb��[�;�M�9�uF�r��S�+{�Ҟ��|<S�� ��Q�z�.�a��[���X�����é<,Wd^􅝳���o�>O��������/��G��l���T(s�Sӹ�9��j�uO��m����͹��I9)�ڕ}�x�ܿ�P^{�s\�{�d�ѡ|�s�K�����w��ɥǖO��>d��rn}O7H}�������h_�;��_Qۆ��^�_������5gIM���tF�ڣ_������eck�|S���L���X}b�k��������dzxB_��j����=P(�@���������&=�K��+?8�ʨ;���%xL�V��11�l���ԭ�d�+���Σ���`Ogc��#�������ݙ��3۷��=���=��䤛��t�)4�d���x!'�eM��v1�kDw*9V0;A��o�V·	�zf~�����z�9����r�`ㄥ��a�eբ�J-*�Kx�zM��|!�XT�5��dŹx7U�Y��zf�M���E����\�K��bP4�lR�Kߐ�d2�aր�YPWIZ�
�#�w�*�7�0ؽp����oUJ�� ����\S���k)}��c�H���+�L��~�2m86x�A��|�c�40H�Uz(<X�K�1:����<:c8D�gg��l�-5�M����V���XX��Ec�����cT؁P�:���\<�C��<�-z͡'�N�Ei�E� ���5��s-,����|n�%�z��ܣ�0�Q@��l�?�.#��~�c�U���X���m5(�� �0���:�+���U@qPǝ���"8i��*+E�'-,x���Be�8q�aA�|\.��COL��2&&r�}w�̡��K�� �j��\���w��t�Xa=$;.���F�T2�A(�U�qxPG�P	��3x`C,@q�\��T�`�ߑ�~�#���\�:��?���d,3��9��J/vG�}�"7%7B���.��Ce���C	�\1
���yQ���æر�-e�������w232ұ�L,�_��{���m6�=��K��W��!��G
Ѭ~��
�n��J��"8���,l�{?R`s��]fU�K�d��f��C9W7�deu�TJuC�&I�;;T,��
�� UEN�������MYӝ��![��z>PS	����3}��UP�RWԌ���I�t �{O�8f���2��g���}o+��E��~ ��W_��,��P� �
��9A�ܻ�@�����yD���P3���)��4�hb�i/<�d�i��s6&5�?�dTSt����rg�X�N@97��J�#�v��f�@������K�֭�ܻs[�\�3}/�NԆ�	)\���Zq��aA�N��o����U�	/�Mf��ഭ�%3���^�j����Y��6���o��fw(=Sk���'2�dG�(2
���Fk�`U�~Xf�@o�]�<���UU�˚����9�O������@�+�+	��aY��˚��s�a�׃��$%�{�0�"�ֳ��(�Ld�"�l��GBn�k��d=]���z\q���c�Ǒ�ˆ�\e��߻H�.�~Ǡ7�]��P�s�����G
j�����c��{LN�b�tB�u����%jŒ*�_3��k� ��$���CP�1]�i:���SY<���o�ˆ~��n��������g���^{M��]�݅��k�q��K(*�M�0Iźͅ��D��ɱ��~.���z_}ҹ�1�?@�pw"��Q�/m_�g��!�6wd��5T 
-kn�z/_�q�Y���s|��/c��ǰ>��������7V.�g��~Tn5�xu
+�h�qgɄ�໱�% �.�h�Hrt�p�Z���9�����������E�㸶ڕ�5yQ6Z���ͦ��S��ރ@�f���ŞO���eA�`���Bh2������xV�0�΢�V��<Ӡ�e�d��˅���2_�/��/֟�<��!���$��gf.�	fkn�ϙ)(��U�n��dtP��z�	��~޺�v���W�|�����}�'%��C}�0!�H�\v�2�t�N�b�.3�R�̗Vԋ>P�&����L����X�'�30q����*ǋ1efYH������8ųA�-3�rf�RLk���OR��S
"K	೨tlp �pZ�Ԙ�`cD��E�q㳠J�a����Ft�T��z���牵��8'���M�~n����I�O���[��s������D�������	Z����g��M��/r׸W�C�IH�j$3|Kf��jz�8�� �3uB�O$���~f�%�D`4���6,ʰQ;JE3��]��e%��Evgi�Փ	Dc:��aLs��ٹ��sT��vl��K:3��f*�	�<6J$��\T��ݕwn�,m �x޸��l�N`hwP;�n�H�3�W�A囌FnL��l �P���rV�|���76([M����v<K�:��^Xso�  ��0hE�A+Mrtp �ݣ���J_���ν���g���0d�WIiu���Y�4΂���$ ���]�=)�ݮ��3�����<�}[ ��@�'��C�A� 2���X�`@zW��8GG#���r�V�zU8 ��b��=ww�	�u���P
@H�-Y�|j�4�
���#�J�*��~�@���]dc�3�_f����Q&  ~|�NM��ıA)��(2�x߅juP|T~�3�a�c�9��0x��O?M�q�Z��c ��� �!*À�S�D꽸��Vv"S����{9������dL\U3�p���IF���hc2S'�T�E	��i�<C�
{V򬺭)��)�p��?����ד�Dz��V�^�aVA!_�O����F7��=�듼�4s���V��p��H�e(K^��7~.��}UAa%��B *�j��=���^;�C���Y�,�'T��Q������w
_��@-3V�7�]�4+o-/l@�e�zvLX�����Y=�Z��1�]���/S|�s�MF���( ���7s�� ��;D}2��c�lw��y��ֹ�xr��K�hp�ase�&��������]�?��=���X���CE��4u�,5��T8�"�rw�R�V�dp�dȶ�kf�Ȱ-�'2��z��V���b(?��!(���N���-��b�6~�g���P@?)���#�P7V�D���\NG�$}�Zޣ2|Omʵ�W��g_��.]�MI��l��m�2�þ�	���b+3� �O����q��\/q�,���asa�21��fp��L���� z2��z�� 8�K���:��@���:�Aw�G� �2��exJ��Thż�=�mAr��u(����xYb,UM�,�Z�l�f��g���2�fMM�|fŭi|�X���LͰm;M��&Hm��	8��j����z䯦}�}�WU]�3��9n�N�(=�`���/;Na�\���HL����Z��r ��g�ƣ�,c_�@BOC�s��U������-Çh�p S��r]@�}�P��#ӲH��t�Q�::��on `��$?�z��ǧ���������Wz2X�P�0c����Y��@��:����{3��X9���T�ij�,6�o�%��(���@���a� 7g!/�7�����r4��`��9"��Z)�(;��`��tDC�����rwz"{Մ���pzZ��Ԙ>l?��3?�z,�Q�FG���|$ˑܚ��ɱ�u�����!#��z������y��0+�$}m擊"��LTjɍ�h9�}�+����ف�{F���%A勨��������;;�g="@ފn^0f�Y�9�����1�q����`�P���Ơ��>f�3�MԒ���"'�/����"3��h;.�t<#��!�[��&c�ٴd�����Q����Ɏ6&�������#��3�?PRA��Y �8�Xݠ�@�x`,�����-�����%D��3��~aA Fma�zt�|��ߕ[}$�5������a}4q�{C�2w�rˌB����������EiklΙg?({��Mٻ�|��g	��l�QB`��N��Qt��"�|��d�����{	4�m��'�Dg�䒙���,��S���:��ҹ��39�j��r��2��{�fu ���+���zD��n�`_�z�-6��� ���+��@����	��UYW����!#����?0K���/�>�=��,2�낙?������-j)��J����K/����}�U�˪�L��i�� #ʦ��Ԧ�\�����0�C(M���r.�с���W�X�{�my�C݋ ���L�![7��4���NҲr����k$�e�Jo�l��ݿ��:�(Ѡw���Iu&���ln��"�#=3����^k������m���g�Z���O����o"�d�+��<q�pF@��V�{����>PeBg9ix����g+p�w:�y��]ќ;EV�k�s��:i��� e��JR���q�'(�Gf:D��p_�]ښ��^1�qaj�&��@�&	�ŝ�|���ƥ��q��>�3k�7yb����p��}���gw�ɝӉ�u�j�sGMp��Bf�k��NI�ճr� �u1ԑ�G�^�x�VM��S������&;�U��10w�:�y`� ��g?���S�7F#��V�������� �=���˹���ʀk��?��Q�|��ߎ����_4�_��Ѧ�C
w	�9�߻�@��������������<���d�oB��2(v	0��˥���M�<H��s�㲴�'�Ȓ��L�u|͔��e���2\��df�
� ���h��O���ʮ�ˠ�@���ϽO}z�{F��@����+"-��s�Z}M�-��ؚeV0�j6J8&���/D,{�۳�u�7�l"�q����r�N�N3�F���^���4n����A1��X1DG3��:�D\09�r�d��֭jZ�5�Lu�(,(�Qʘ�G7�Q�P+�E�w������-�&+ �I���f���r��&/>uC�Թ\�cu|v*Cd���'g����:q���t�糥�)�ۄ*]���RuA���$�8ׅ|9ȷ>��|�_��v����Y������[o������`N-��P'�-�����ވN��ܟ[BI��Y<H7�b�jܜ������{Cy���r�;�2������y�N�����.FF�C��l&O����=+�_�!����N���O�'�n�;{�(����ċ��o�F9��9�� �0��T~x�=�=ؓ��e�/����+�����i��mO��ۜ�����!���2z|<7@ˑ:k��8��a��dұ��<Y�CZ����{�H���m9;�`�:�
\Q3Ț���5�uQSУ�W6���SSa\��҅-�X�pdz��̅�%��Ll$�8P���33��k2����hd�&�Y���-,CX����f�[f.q�Ϣ�W�l"�XU�3���p;]��'/�rcS6��^���s��EF�2R��#���G�2��tc��g��Eo���>�&u�� �>T����X~��?�4��F~*t _|�3|N�Y�M��j���Xc��2�Q[ޫ�O���)�oB ����Q%;
p�� � �tZ�u��y�n � 4B�6�m���L'S���c �	�L(����;9<�&7G a�H;)�zށ��t4a&6�@d�j`�Z��Ҩ9����:sl��Dϧ��c�24������U�����z�G�wek}�qd��þǫrI����L��u�@������@5���!�00._�җx��Z�~d/]��s�`>��z��69�O#�3���%�z>n��^G��>7�4�d���.����JF�q}3Ԫ�x0�ĕG�A)+���z�^�R'����}������c���3G��S��!S>m�f��'�������-V���k39�M�'�EIhK2��Y�--'^�� i}�����fN0��ˎ��Ҹu�n���H�����~�/-��V^x`��ѕkj5Բ*Y>'�ϓ�LO��d���A�� ��$��c 7�t���3����
�Y IԈ���Xf�����>U���n�w 9L:�j���?յ����>=�Qї
1dudl��G!�gjEq,��tL�����g�'����bkj��.���(U#@�~�`u��p�@c&�<���r��YU?���@�w�'.��y�����]��b��׊�+��,![��R���s�Q]4Ͱ޺І@%L�\������\W?b�`v�ˤCpIa.�%p*�`�?��}�����c���y ~X,.���3�¶�	�:l��v�~����9�=q�Ĺpd�F5mYZW�����=�	��TA��������}v
+�Z�'��y�G�9pnη^��]N�?y�ߋ�'��`8 �U>o����4��@��&[T�2�e�,i=�jL�~Yf`0պ.���:��K�j@�8����t(�c.�j���8�����q���R&���Y�X�UDך{j+y>n&�@0��>��98���%���r��e����m��&��������|����G��H��|���`S��_�������>��~�{r�<�&�5k�FcEʿ�ҷ�/���	1��j!�{q�&��ț?��뀞d��O`�n֗���Hr�h�F�h����/o�)�2���A��E�4�q��yN����s_���.�0ce�TXe��H~���O>���c���ˁ|��/�!��r6=���nsuC�:��_��w?��f'2.RC��]_Oz�W�=I�E��5R�~r�C����ta����S���1j��Y�}�B,Ef�fX�i{O��v�H!�
W��r(2�j4:Su��b@2w�K[������>���9���{���dF�@�*7=<����#���^u=F��
�.n���_(�;�L�j�n>���,0�U��Y��N�c�$�[n��'��v畉.!�X��@4���x43u�`8��Z�tuEJ1�l�0�Fk�X+h�q"�^�f���� 
�x����~��$�� hr_�^Y撽�;6t��8
���R����L7�5}.
�{����:�{^I��� ����b؆�ș䜰6$s��ĞK��	DKz�\��GdY�}�g4m?>���� |Bmm�#oL?��lDeHUGb���ʣ^jMs>�����������SR)��&�$���;�#b����� �q��8 �融��D�3��TF�v�U�m_@ټ��%��ݏ�)�ǁP ��xឹ��|����P�z�)y���Q,\�&�-z�38��8gP�ۦ������U4�>g�2R��Z,$kA�4ў���e��kA��jIY㉾f�h�2�[�im�P6��<SYz͠���ߞ�B��~��� '��_O��B���%�	�����������F��H���m́Dlt��3,fǪ�����6E66�j͊�r
��vǂ!�$uW�p*��W�byG�{��3 �DDƇ�:����&%sfC�!���c?��������L���Y?R����IT�n(u���2�k{� H����ϧyk3g�jX�Z�/4����A6��?,�)-ّ��	�T^s�R�f �ƥ���J  Y�e����~���'�f�JguE������`���Q�$2�|��?�+�. C`��H23:\�R�#�x�j��ѝ�H�n�C�^d>N�c�$ �s��l������I[+=��0�h�xJ��l�́]0��.N�Vn`���-�����)��]J_6�U̟�  �Yd@�q���m�����i!��7��i��-| �Au�4f�	�Q��o4��|i�e�yV`]r�����&U��U��Ƴᚷ��D�,xP��)&Xa�=�����"X��^"�3*R�"H>�������/	�^S�L4Kĝ�<� �6]@%U5��Q�����\%?qųX�V���������%�܃�;����e��ɏE9��R�X =5 �V���K��Wr|p$��� 8��ꄼ������������/ۛ[��_����׾,�/\���~F��b�j�Z��J��]�o}��_��!� G����2�I��g�������.��\����7�O3�<��e��6v�� �1��Y��0�YR�s=Y�.ꓗ�}��
�l�^���Td��R`A�C��hskS��̋ҋw)3���I���/�P=�ܑ۟ޖ#���@>��+�ڕ��boUF�D?zx���;ť�7<�/���A��4!��cu�u.�q�{�;e�9�v�!˞���b-`r��a��&��Cqs��>��W&�CӓY}'��bd.pEz���{�<@'���׸ҡ���6#�/����׭�	�U�<8���Am���ӱn,�T�E�8�v�NG졳2ܖC�*�3
ͩ�:R��t��?���rr4b���9�mJW�R0IS7���%c�k�<�Z�������N�m���r"0�I�Q"��4qS�2Ũ�;SQ#}v|f�$���m��ٝ�T��r8Z��1J�����u��Y�u�f�����l�\`/���CY����y->O���bƬ
�a/�n�4gd�1�� h(���G�"# e����h� s.Z��# 2�W��53:~��[�A�>Qg��D]_��i��f0���d�Jֳٱ����C`B����F�A`�ϋ�k�x�Z�qT��D�#>��	 �o���V��|En���P�TM|�
�z o_��Y��G�����{u�\�ʿ����	5Z�����Ϙ�D��]���z�����8U��\�%|S��:а���҅G��0JK=�]%=	Dz��1��Z0 �Xn4v����9
D�Rg����_���o{9��Fk��ә���!lpj�63�̤ym\V�j�@��A�5��>�W� [=t���B���2I����0h�Ȣ�,#���Ad��*/�^���V��R��d9��랏���Z��}���^|�c��A�0Ѥ]Dڠ&b�1��>/�w���2��l;.�Q�/�Qx���S�^�%��y��E�����[J��Q�n;$"�	�&J�I_N�[N������F �{K�,`���K&�T�Cl@� =��A-[�7\e+���U�
M�3Z�d<�#�S��	����8P�qow�-��*1�$��]QQ��댏��χ�Jh�ѩ��
��n�n�{�.�A���ʋz�/?�<�~��ƺw�ݚ��t�����}��`�ؚ�&�-.����1���u}�r*/�R�:���S���j;����K?�hh�&\ܡ��^�\f6(R)I�*��IP�����&�7�'5��d�?��.
�1FPA8�~&��pL�)c�����1,3�37P���,�ap��@Y���k;!1��H�gz$�2����v#ǀu�D;�2ZS��j'"��_���2"���lU��Β�[PV�g�3����,��d5�	��X/�Y���W �%���.{�@^T�������rpz*+���yy]��/�g�yF�xG��|���k_��\l�r<��G ų�8���ө���˟�����ʆ|�7��|��䣃����������w����B��LQ��*�~z&���΋�}�Z��F�r{4�YL����֚�NC��^�B�T�����l,�> %�3+卧�W��Uy]A��{����˟�kkr��m��;o�^5�C;(�=Rб���8_��e���^�UEHR�������F���51���͙�A�i,=��B�h�zc�cs�5@eQ�
�=�0��X��ĳ �9��s2���4e(t�d���ljǖ�����)+����/�P��wIes$�G��v�`�$�76Wes{�T5
��1*��* L�Vv��3>㦵���k����K��$�c(8b�� 
s���� ��]ʃ�ۧ�2�� f*Z�;� �9��Li������)4�[��٫0A�*����'�`ŀdf�(poz�.ĝ "���.u�?3[:Q����ŝ��hv$����n�օK��L��LNP(X0��{�� ��q��K�f��r�ު�i��e� *������m�H/ZD��o�
� �v>���{��)[�(t��^�I|P87�~��>PSq~��L]� `��瞓_���/8h9{�x�Jn����{4��\G��K���������q]8h�������|��3��/~��N��NH�`P`�e����((�P=ڵ�!�>[sྡྷ^cB��k��߯^�J�L$@�e"�s�@ܞ�����L��ޫ�b����^+��N�$�	�&t�8/&ȖM�q U_��-���J�%����J
����w�l��Қ���>�/�
p>��./�R�R�Ԃ;�3qRa˦j�.f"����i����笚s?����ī`H���7~�Z ���[���k��<*����]O�JF�8��6�H!��Z�*��5��կ��w����J�]�:����j�@ӟ��e��P�{��+[� ��Zmj�lx����<�>c|�ŏ� :�l>��0�=9<��A	���,wNM����p(L`(�܃�%.�I5�|��
�`P,sS�CI��օ�Y�7_ҷ`�f�ݞQ#�=f��>�'�A (ɸۄM�M�5�E��F�,��Ih��M�=c�#�b��gk��올���5(�Xʒ�H=�=�dL�P�eVP��o�Q xΤ�4e֌�cQ69��Yg����X��tn �P��n��`��eфQR���/� g�jw��5�^�I3�����s?�ʅ�%�xѯ9?	�cY3���<��҂Cɩ����,e�9u�?;e���s��Z�:���b`KcD���̐�Q��9��i����+���>Oj-��	S+�4��/�1+�uIΧ���HIFa4�uZA�l-�#�@�j5�F},y�x�c��&�o�B$vrpd=�}u�o��k9���bW棙\��g���ƞ�kL������?���!��ߔ����n=��;Ӆ���:Q�V�regK6�[.J�u���&u��m�8�}~��_�W��5�u2���젘5�%�>�@���!�$K�V4�y&1�-ZZ?�Xd�,BD��q��[��$)��gg����ьTAJg2���@�����M�����E�%P ��=�#̩:�PdBT
c>��t @�
R�|���?J���o�ߋ��O9h1lG ���F��� h�4V�����SD�^�l��J&��"��@y�R/����*��!@q�U��U�0����Y8����'p�g�����,�)N��h*g�þuN=s��>8���r��@7$�v.ɕ+���O>�u�V	+���඲y��.�[��
Yf����(ljJXؘz�b(���fU�هz�l�4�0\�� �I���f�b�q�tc?2w����m��6��l�MF�
G��=�� ���A������S]O�����	郗���r9�Ou��<#�`0*`��3�	B8�i�f@"#yޥ2o�.��^d�)YZE0��
4�HDo���5�����r��m��>������u���C����J�H�a���URa �����8�F�`.�@�@  �.,Ӈ���(^ly�Ꝭ� �mB2�\�JC�6R���SK穞A=�җ�l�Dh(���b�؜W�= �s+<s�<���c͒`����T�� �q:X�
2�]����"@A/�qi�g�Y�x�����X�"e�Kf?m�*�����A�C8A?Zp�:C�O#�=��Y���F�kY'
i�����5�<d @ąL�zf�q�9ի&���0�T-@��<y�H�`u
��8{��~��2��V�k`�-���2 �M�x��o	�"��Z��_��:^嵯��z��T��̏���'�Fk�0���n�1(�[�WNY����ײcݛ���^����Ж��e���GAKe���^��BO6JW�6��VO"���Ŗk�������	����(��=��#v6�f��
���!����9�,�L!�g�4,)��BM*�{��`��j��0�`�P�{��4z8�S�{%�������3�%�YK!��y��5�q�^�)4*�%T^���U� ��hy�~���C9U� >�V����� �҉l��x�Vv���-Sc_�*�{�R'3�upQ<�'��
_>,�-�n��l�!O%�	��^��{����唹jUc�*��2����g5��o�x[�y���������ZV��Q���SY0;�,0��a������e���P7����E���+��0\~3< Gы��k�F|ƌ&F�o�
]�&V���:��/������_�yd-��_�c����~�v�@!d��e���їA��Mn�9�ڐֵrN[eq?nDW�x�t�M���2���= "��1@�^{���@7^d'�T>���]$�W^�z~ӂ�cP���6�;���i7�St�[+�RO;�.-���զ<��/�,�6�کn1�S�l���	�ho==A����4��C�)� b5�5��K9�ݗ�ݖϼ�-�V�(*sz*#5*��7�K7^�+��2Q�y�[���M�A�F}���j�������-�6 �ͻ%(S�!����I�'.�UD��	���!����b�v.
��9�K�Hv,�W���=P��Ռ����B�U°ד�R�r��ˣ!=��
��e2
	�"Ot��<�Ŏ\�&-Ia��� n����t�9�����P��g؇=��!/���.H��ÿ��,3
t�w�z�ǧ�z��h�4��	�)�a��)2�M�|�D���/-VC���59M�� �1}������YS��������c��T]l���>�\/qk�)�G�z���l����\���:#dl���BOF�?E{��`C���%�+s(4�YoJ�g�;P���tj������R꺒u�-�]�&�Y#�}��ۤF"+��0��ܠ�.Z.ܺu�mPg����"����Vb+��3F����<�_��1����Z ����
�&w޳��YV�����yeR� R���d�"Zm=��8l݃�0j"��y;3�
���{84��=������((�#o[�����Z�ZI5jqN����}ҫ]?�P�l9�<iY$@��S��Q@c�h1�`2�Aj��e]3Ty��{�����p����T��{wɞ��iÄ�	Dd&f#�;8���U�� �����W3V��V�F��[�s��iꦥ4WWZH���3AQCǳ���z3ȥ��fU5�nT.F
�d�,��PQ�8n� yV5���TN���i�o��_�c�>O�[�`���@�޳Z�W<[!���ؼ��tЬ��K��ͯ���FiIYݟ{�猭mz �,o�k�+������p}�	��Ts���g��1X*C��e��`<C��*�	�E��g�Md�P{��2���PVW�V�Xc�ZP�m�=���E"-�ک�6��V�����}J�+������C�(�(|���"({��X}��]�MsR�+���[b���z�7�m�o��g���o����e�Z?�o^_�J6,��#c[2�B*8ܹe��H@h��Yϕ��^�	��Al�Q�߸�^��`a���/M�Y���Z�9���q�$��=��fPi���<��&6,G�5OMBB*�4�,YNY����)&f���5��W������89�#��{{߹�_A����������콁��y���v{��;\]o	���&���ծ����%��6f��M�_Y��v��-���g�U����(���̑����bj��(W1.��HNg��z�������,\��=��}��8Ƥ�QoCM�,9g��{_�����Q3�n�e�:7=(��*@)|n�[���;��F��,R����J��$��xM�|m[NP����\�_>�#���P��.��+��0P5�����
#�zS_P�S�Z��oB�S�<࠭(l���r��U)�,��Q��n+�/�0)dY�P��'L9�F���)F�Lл�Q���6�@ 
�C����),�F�z�t"{���bE�Gc)��ȡ�A2�ֺ@��K �vz��ܐ�K=n�]��Ph�eNI>�zcG._���SP�\�ocF.C�[1&ԫ������:�Y��O����|�����B���l���>�zPw���%����Q �(�P��S�g��ǆf��p�[an����Δ�7�!�@6Q�p.-? ��np�^eY�NtO�X3�ܵg�w|�k|uSz�6~����K/���w�N�b��WP]��k�5���u;&*��d6j�+��]�gCt7���T@�.A�Ƈ�̫�����׾)��WTn}��'?��/r�8��9�`\M�B9�L��'��� �sԪ�I��� �&���7�	,����;w(�Ue���ʃ�ئ�F�ׯg�߭�d�E-[�5�Tzƍt�= 	NI�5��f��m��Eg@k�H��?�y���ܼ����-�ㄚʨ�D�	�%F5jBy4TS����>���E\Z��Wd���9������LD$ka�@QvQ2뿡N��t҉��ή���"3vLԀ���X����2eE,R��|ё�߉^����f�>���p�ͩ< �k,P�;��En��o�qLվ��v*"Cg{VV�,%����/L؃�G��[Ř�؂��T�̲�)&��ϡh�N[f�6.�n��pb���,g�_E���3��ڸ��E͛����P_F�ͭ����ۑ�'��f�=�
�y��������g��+k|�Dj�\KV���~�=C�&�Fd�/��2���3G~����,�g=������'����L4+�$H��#��{h�~꿻R���6.y�";w�mݒ��	X]i��Y��٨�N,Hj�; ]�]���3���y������DP���)賔z�ˎ�gT"�ά�,��E�b�ʬ�3�Y�^ɛ@�%�-�C�7�[�j�d���X���V9&
fA�]`����?�أ􋴟�V"��I;�� JKp����C.�m���Es��E�>ByG��B;|��Yj|���K�
�US<����x� ev8oK�E��{#�\G$�}2���$�z�ϥ���	���,5M����u���4G/�}1v�����t���㚠�S2��Hq�<��1�������z�5��b�@�t:�l���T�ŧ��g_�ao���Le�L�l^��K5U�8��f��܁���RP�p��J��M*L�,D�0��5�6�P󨤹���g��Ȉ��j�<@�
�\9���_���l9�\߸ �d����ʪ:��|�U�8ؔ{G�dj�J_�O��`��l)XX�V���x&��#R�N���~X���ٸ�S��N�����K���#�X\8��c�Z�,��ǨPC�ˍ���׾"�{���{���hO��:g�r�ư��������NQ_���d���lٓ��I�D%�9x�0Yzoۃ5����J6�6�Z{�hON���k����\K��Odr8�%C�+ix���W�4Bd�zz�
�ǖQ�����5#�� t��d�&�p���N���m;U�P_�D��ں�Ee�q�+:^x�9�t����C���ߓ��]�qB;u�������+�d8?ѓ�Qu���,��Jc��E$�6�u��`�����c�1k��S �~�-&f�9靨�,�:9��37������w�]��W%������N�4�ׯ˿�o�[�����U���MJ�wW�g_��]FyǥQ@�B�$T&h�0��~�N3����>Dz��K�t]Чݫy���ͯ}C��=���}*�"v��%y���	�:�s�]Ÿa#�P����F�-B�`�A�;�O�*�
��9����BCx )�+��aɞX� -\"���銡�	�+�>�fO���,�qt���� n����fz��My��7	��y���!1����+2��>�Ȫ⚿��J��tϸ���59�kzl�{P΁� ������@���D��i�=��q1*�%T\a+����\j?���d�с�્%uw}E�?}�m9��/�rgW����M�%�O��w�^YZ��7�NB�&wz�;c!����:�؄i���^s�)�QZ�L��koQ��\�Ə�fwo��E韔�xlڹԪ#�0B�Ԣ��QJ4`أM��yI���#�:ܩ%c	�5j#:��?״X�z߯RS�6���je6MZʾ����T�B��^��Ev�	e��ʯ	�F���ۤZo��-�<���Z�A�eM�"� \�9���Uf�>���{3�Wf��C�Gf����������)E0���u�
�k|cnhg3k���k7��r�㫸~�\@#��H�>�r���YL� L���P�%�#݋N�E󖙗e�B�2��W�JF��~
���Yȴ?g�#2и�����s��{�ʩ���2��	X5-�|4��5���`�2���}�cP&/ѩ\�'���`F&h�lI��.�f��2t�%���G�ϖ&��.�ͼ#BV5~�p<$#�#���O�ڎA�܆U�3.�9%qT,NY��y���6 ���x��O�"���]�*��~~��f�u�x�4��8~�J��kR�����bX�v}P|`�Tp���Yu��4��M���.�8ؐ��������U�4^)�2lEGsu�/�lF�$R��w��mFT`��fc�vᒬm���7���>�
(<f�m&�*q~��/6���96��)0NӒ�.!k�Z�����Gn��ųN�h����}ģ��
^<)40^�d�vյ��
��կ�W��%.Nȣ/OF����Ó#y��w�Ó]�^{k��f>�ˇ���'G�r�is�"�\V�.]��v_���htW&ق���Z�-��]s��\m�q{�T�th]���ּ�l+#ꈜ�&r��|�d��*u�?�{O���׶ek�#�d��SC�+��ﰖN(j0�� R#,�r �T�JׄLzvD��J�tn���o{�!?��=OdKA��O�,_~�Uy����x"k]8�S��}B-�jO�0��9)�̶t,�QxP�P+��H�cߚ�T�eG6:� b�L�,�̆#ɦ�IVuz樭��7�Tv��e� eB�=��9�;=�rᲂ�ge��D>��	���r�������:��{�3r��"�c:�tjc��;j�ĝ,7|FQw{��fC"�ܦ[��\��۶q{��Ԓ� +f�VV��	�~;}��?��lץ�k������ ���}���R��)��Q%�|nl���ƎL�Frv<R��#͑}!K��u���UПmN)������r;��ޕ�ڵz<� ��"Z]�<�ǧ�?����˗��"��h&2M �P� ��5�S�����-y��?uF�5,�̦r��]���!놬i�z\�b3pB�?�g�EkB��jgd�|E���^?�}G!��/�K�� �
�T�m���w��u���p�P��m ��zя�@V�>l�촳�jg�&�P��7�2n�%w����0�m�ƒ��`?F{	dd���rx:V�/��>}�W._���r����>��Ne�}��y|z �D�um���!`�7B6ec���W�&Ѝ4����4�V9l��me#%[P%k�1��J�B�,qE�]��X��3�cUZv2�B$@�����/b���Bp���&H�!�S�t*����v��V����t���^���5��W.�% ŀF������+�]f6��ZQ��.s1���]e�2-�����u��J��QKؖa���??�<3ی�
�e{oF�٥��Nm�ٜM�=��� �s_y�[(%C 
��Ų�Nv�����X`�ߊ�q[ 5��A�����Y=�e����z"��3�s�����4���pU�XN�-�:
h�O�)����2c�.�|��Y`l�:�(k��E����jɁ��t{-��H���%uI�5�#��	��>�I�����.QM�%$�pS���w�T�o�lf��cs�<���1ON�8O��D`|�������)�`��MEy1�Zyi\�]�y�Kڎ�.�M��ҁ��<l�P��F�=�'|I��)����D�_
["�Oz����#U�>Pje�����}y�#��ư�f��˫�\ȶn����e�����penWMߒ���e��٬�!땜��^^W��7�XV��_�ӌL��鱜���G�oɽ��:f�H���u
:�}|��C�	w�R�pȨ�0Y�.e�f� dI�]�M)�_FU�FL�����c�%i�S���x>�Mil�?���T��
2]u�@/��ӱE���eE��T�ω���~�cy��{�qy� h�&�]� ���g�A�?U���yC���G��׾,�z�m4�>�όn��bM��1���*��4�,a�7�ަcjM�f� ��ib���u��7�ނ��>�+��O�qh$��ߒnesj�xRP#�^�?���F�E��RVz����J.gGTó.�'o)�L<Z{�v��ꦼ?�%5��[�^���Wo�JX��f��Է�֗���n��T��*ZDj�Xk��Yx�E�t!g�D%��j.�S@3��g����w��)��F��"�@��
�e�P���u�t��݉LGc7���Dk�#�c]Ck
x�䭮iH�Q�u;V�@ ���P��x�B�GKn�j�,�����`]�=I�V��q��^���;X�˗v�읜�HAS�l]�a�	�9Ext\7�e�����t�)`;�$�����(/��u�`/����L�1�d���v�k��^\�J��	@-�H�̍瞗��dE�)?
��џ��K1�����u�w�ޕ��=R'8=:����i��#��2����p�}�J� ��<6Dlna��
�� gu�'i�^Kބ�]����������������RX)R�L��rl����d{gG�HJ��o��Ϥ'�����":�{-
\R==��)c�ng�{$�T��'�����4���R��� !�ʤ �3ҭP绷w(���@f� OG�������x��eUmMWR7Io��������{:>�D�?�O(�v��e���^W\���'|�:_ 9�@���I�	mm��+�ߖ �)��U��<�P�YK�1ϖ�,�X��u�r�)s�Hw��A3d.`'V��L.ho}V�j}��:X��"�B�A��Z���n!��LS�������y��$�0L���<��'��y�Z 8�>�����@KR�(��hdX��2�:�N��������@�����dy�T���͈��K�$VY��Q���d��~��o�DX�U����~#�az�a<Z�7���5l��
�+s��CdgT�������@BT�/��LHK�ս�`2�S��&.�eD�/n�޲2V	������v`�q�P�J���;M��3:���˨����2i�-3g�5~m
���'���PU�E��+`_e�~�ew\�K/�MR'�Z�=@h�2b[[���}2c���H���������Z}�����Խt]�_�n�c١��y�fcf٧w0�ҧH�U^�Lނ'�,{�	��������|�' ����ì��M�$���}5��2v�W��Q�e��$i�����FC���M��p}��Vx����=-�2���0��l�ߑu��F�M}��0&i a�PY	�X����"z�-3{w���eJ��C�p�Ǉ�r<9����r81ꎞ}k����p�Ӈ�e?P�,�0����IJ���f��k��`u���JGְN�3A���cy���9�c�+�#�'l�5��K\Hџ�;8T��ṵt�#}p�=�YC/��_|Yv�>8>��} �g{����?L T3�F'2�F�:���ۧ�.�����d̼�YS]�1�[�Wɍ���s7,� �y�G��ۃk�0j4�#���輥| ���i� �2�0TC�:  e�4e� �t����%w�����ERpу����:}��foH�3�X!�C/Y� s��@�^h�s�@J��(2���3�:�0%�=47��`@c���1C��5�ܳ��3,d��^��DP��K��}uN�7i�Ţk5���X�HJ֣���$��:�ߣq;V���S�%� �x�f�Sd��6��%2�W��&�F��̓E�4�h`�j�g���,���*�$�����)8\��gA��\ �T�8D���]�S�B��?й�[�pc�M�?�wG��*زy_FMcDף{��\��g
䖬1��������nDP��3y��!��׮�O~�s���o��| h%3��2~�&5�V֛�Z?��	�"'� �M��1��S
� �G�����^{M�ݻGJ)60���� x�30�Q[m3�G��Q�М��t:&����3� � �X ����Pb.��a�oo]�o}�[r��<�[o�ů��3�j���׿��Z�ׁLg�;@_�ߢ�0�����F�s�_�ʫl�R�y���6�)F1�}|[��{�M�IG�s2؂��}w�E��@����S�Jډn���\���ԁ��!�^��s�§0��	��eE-�1���b�}/��t�ȼ�|��L����}�J~� ��
gF�XL��:�oA)�5/�ȽAvQ;�Q��	fK߬�3�W�6)}�b>�Ʉ!���/L�?k
��L|f�~:��f��v���eessiۇ�,P����40�1���z�ʁB�٘UK�r�9z�f��^�I[�Ų'�)^�*;/�$ןȫ�w�yo�*��9�����sS�`�����Ad� ,}������3&���7�x����$�܎������?e�x=�~Y{�R����LF���޿,�g��1��ڍ쒹b���I�!����^�@Sg�ǃ��U�f>kV&���5SءS<�������I)��h�Lg�ಲ��d�Ό��u������W�?�}f8\�1����!�co{���~����N!:��pWyf�$c�׽��#��6��k��f��ϼ,�/]��Ӊ���ln������wl��!�f��N1��:9BK��gE��Bz��E�C�؂IQ1��i����u�N�n��!�7S+�N���K"��=���M���B��612�-t���sf�8�pà�Z�	Q�,#��M�qw#;����Q��i�;YB(�-�s���8��,�><���|���_��"�U����J!{'G�ԧ�"ё:�Ýd��4���[�a�{Iq	�~
�赝�S
�F6����=�j�T�r���Ip�1f^��?�-�QW]Չ��c��6�lc�D�嘆�@R��}��뤇C��}���<���Xvա��/��l^�,�������d�,݋+�~���m�%���Ou�����Ϊ\-2?9�cWlmQ�c�V�7�&k$���l���x2Sf�r��Q�!��f?�1�� ��s^��l:�a��3)x�ޅ�w���d9�^2���T����?C��p2�O�r�����#~m���*Б�vC��#�2�x�WP���*~�X7����������3�wp:>Q�2�L��֙1�ҲA?�qXHl�!ߎ�����zӗ�@6C'��"K�{Ł��R�i=X��wt�����B�I`��z/f�|ϋ�پ(��1)p0�g�B�A��:�Z��r^@�g*�=C�L%:�Bd㈯��q~������92�1�t{�����3sNp��r��Q	�Q��;U'}\�-+ u`�Pǰ�>��j_�v6�y�2s	��Tz���!��+R.�DO ��T�ѣ�Ҩ�^�g9\� ��y�mj�n���Jg�^�g�:;�}�[Bx&k��)Yw4f�}���2dM!j��������@�`��4�O�7q�awBb�	�Ϡ���p��ߡ3����ɭ�n1z��F6���?�`"[	J,����C��1Q�����o���¡Ɵ��g2\Z�އzö`Lʴ�?M�>�d=)�'oLm���e2:_�w�18����ܒ�ί
�ފL��OF�-L�>]�~�
؝A��鲬�X�F��O�X��T�_�����ؿ�+2maYE��b; �z*>`�۷4�r�]��� <���`����X@˲=���ƾ��ef�W�l3���.	�������͚-9�+���g>w�j@U�
@(�Cs��")��j�^���������������#��!;d���M�")� �$ b,Ԁ���|�!3������sQ )����s�����{�M)<v��TH���<��K�X{ŝ��ss6��"Z�:b.$��������E�ey �F[���k�{��x��y���#��-�
����}�h�G���&���̣��hߏ;�z�`:w�a��!����)� {TB����F8�i[�+�bS��ȏGT��=�5�a��-�0���l��V��$ �_j�p����u�M��%ԧ�uoB�s�9�5�1�]/蓡O2Z �E�ft<eX6�k���M����X|(W%n��^e�4�����DO���C�o��+l��5�y}Ȉ��Bxb������:&��ra�LDʪ
��To���GGj��������wdw���H�z��]�N�C� �I��x�2u�a6_��>�5�x�@_y�������������3�#Li��m��ʲ��s�;�et½/�O*v�?_u�����f��	6��/�Ѧ*,Λ�W%� O��I៭�����sѿ2��ʔ"Qy����W�^�(�0�~ou��h��H'���:xa��Y?nb���&!�1�>�d>'z�����^��׮���a.�~t$ϜR���JS�叿����}yx�@6W�d����d*�i.K���]ݒ3G{2��d��<�M��'Wܓӛg��^�� u��� ;��!_}�3j�ewp$�LZV@=���C0BA4c��(��A�.V  #*V!�W��LX5œ����o�!
�㼈"��@��/~�#髑�'���=�õ������� �.�޾!{�HwmE��Ͽ"���\f:r��]���ϓrxg���M-�y��BUk��UƗ{��a�`�*��0��a���'�7_H������"��E䢶t�h�:�CG�����]W�l���j��!���6j��X�mJ�sH������#g��{�uQmk?5s��j�2�L�0m����VVNuL* ��5�(�u|�&C]<6�sfF�miV�<σ�J\x�$�{����I�]PC�F�3H�gu���t�m��fS�F^�'��d��<�4�i�6����tUֿ�3�9c��S�O�@�}�@�?;T��R�2V�h�b��~�$_�K`/�<[P&T���f����Ca��Y"�!t�*p(���v� ���	� �ڊ3RNg���0:�I�IK��|�?���=���BMLX�S��X}���F���`,�G=y�@`�����^��o����&�G�&i�#�?�Ծ�9#��x�YY�:�M˘�O�I�7�=oG�W>�����v�B�!֗ԣ}}/ɰ���τ�P�0�╠'/�4,�����G�^3�e�) �ҥK��[�@����	�:�q��~_��� �}ⓟ,�K�,�ao��Px~��A '�o(1Q��F��3T�'�sU Y��`���f�p_O<�A52f:�}�v�ܽ�[����dlY��EK��<6J�#A�4rP�XR#3�u�Y������M�V�T��yD��7�.7'��!gt�gjƽ�鈎Ĥ���7�O���3b��ܘvE�"W$���FFK�����+WWN]ݒN���!�"z;�:a�`�[^���f���D}�ü��d�s����B~3�g ͚��Aģ�Q������9ͨ�Cبj]�_�Ө�������:�A^}qC>M��H�9 �g�� D�$��O hEǧS����ב猲NYH��Ϩ2R�`�#��>����f1nt\��?�!zG^��"H�i�q���9/D��,]l?
��4t�ְv�p�Zڠ��i83��p`���?��b��]�9'U2v��Z�|/�26���k$�6,�J�T�q�ɱ����9+�Q��rqv�;nL�r �v\���V�&͋�d����x7���އ_v�s։;��^�DtD�Ħjw?ړ7~�K�sOg�d#�����!˝e}�ʪ��u(&����	YHh;<>�~�_��3�[ٻ{ ��������ʋ/>'��lI6�s��H�դ�#	N�ũkmo�|�(��@�O�,-_?��G����ݫ��tX��IEy2���7.Lޏ�U}r��*%p
��NR�1���>��ttBG^1�I��9=
hFP�K�#" h�|�vDx"�H�k̲ ~_�n0a\�55���Q��Z|���.L#EEj >�ɭ7�nO���ɥ�.����rk�����~_:j������&���J�W���O��0�Xح�D��~��O_��|��a�Q:��P5����{o�_��=��6�{�JC�}�z���j�%��x�'n`l�� �P��7m67����0-)/�mDh�F+a�&M���?����,��j����o�,����5���/ȋ�ߒ�v����]����/���e9�sJ��׿)�l*�IKF:Y~q��э�䵃[�����V]��bQ�Z�&x	k4S�{����TU�Y�ӯq$
Q',�!0d ���Q_Z��t'�L�CS2C�j�E��7�vh�h�
G
r����葬�x�~_:+m8Qj�@�x�Z�)��
<c5^Q�/��e� ��.i-o��ɦ�0KI�++گ-�m� KR�˲�G`���EZ_�jeN�	�,�'��G:'�5��Xj�r���/5l�S�.��R�E�i�"q��[KK�@���Y�q���6��b��	szu�m�d4�/7�1�#���^A`�͍f3�C�U;k�;Q`֐��@�V��:����QLD�襇�	 �N� ��̓֩j��n�(Os��]����Uk1:�� =en�s��@rP�)P������]�+��s�ɍ{wdГCl��'s*�1�X�3��t$��R�0���& j'�i8�R��Z��q�<ߚT�o5�� �'Ξձ�+���	����3�ȳ�>K/��C��{�l�ha5ǮJ�<�O8����y�?��z�.�իW��bSFN���*�oww��&����1��]���N�.��tXPEh�����-A`	 �J��{��uN��pިr����Ң�����2�$�/�z��}bN�g�_צ���0��bՓ��6k{��Rf*���)�_h�R.�������U<R�����#w��B{.`ΈB��cᄶyO�@l���)��\C1:��H�U�*�nBY��-1%࿡U���'�F�L2�HXQ¸p��)d6ݡ1JI�6��K���Fg�b�z�T�H���u�4B�� nl���[y�0� FH���d��ф��b��9B�`�0�%AO�x~��}��4^c/NN�Q2I@1gI��m쎂�aS
�PQ�b��O<���/o᧵u�S�Ǒ4�SM݇�g�8�,V2� ����RTl�{ޭ�������}��:�YE$)/�E����z�=ݏg����X�x�@ɥ�lƕ��-6�p�\�c\��*�jH�
�����qb�X�y�h��'�o�2��
lbmf|i+CY���l��ܓ_���ܼq�����.���T�?��#�[�iv��n�:�RU��g�?A�����eK�@���?��g ���Q������d��6S��Ԟjɪ^l�J	�c���O���B9�_A���C��8z��n�gт�3��U���5�A%\�D��-�>��-�s^��BJ2sA�ںiv���P�wj�� Q.���p�ZȝI��p�?��P�	�D;��{����r��=�@j�)�bdG�ᷯ��:,C5*���8'����Xc����3*��
���LP@u������%c݉έ��x@�>�(޿{S~��O卻�e��$�2�j��@Ԉ5H@���x͓
b�'�U-G�<
j�yÌI5"����U��yX��+�n������㿕T�ۛ�=�6b�)�Y]R�n"?Q`���`�����;��t�P�[��=�+���'>g\P���Q��;��̓��+ jץSG�B}��	�c�A!]���<�l�آ��"Ҡ��y^YZ�E��q��hGd�΂C���7�7��.��=9�)�eZ����'�7��!����z[V6��s����=ɛ���b~�u:�'�ܔ&!� /����j������vޑ�q.�U�ƈ�Me�	��Ȅ�d�y���݂ǝEYz�́tBZ6G�O�M�FޠW�S�JcI�����_}�4�0����+�0�R�e�V�mym]��5�ؿ-�=sQ�V�����ښ� �qS��Iӈ$$��E̓�����إxIr+��_g��ǆ�g����,�1oI���ը��` Gz�!"' ��Ta����S`����w� d�W�΁zS6�6d���|�a>T���b:�<TDs�:V"��Y��`2bm���mY_�(�9F���eƼ-�H�R�N�gT�����Q�2W��z��  ��o��'�F�N׷6�j`G|js ���x��E~�*�g`��9����
�xp���
���E�N�ۙ@̤�?�Ί#���P-���{��> ��y� v� R������ dB=z!'�X$����x��|Y�d��'�
+�&l�Y��U�+��3ֲ§�O�]�<�u_�]�E?iv�m�'�R��""��9��2jY�]�D�YeK,�:�f������d|�õT�|a��!B'FAk�:�!f�8���Kr�[�q�V��J<<ʝ���,H�"Ɖ9d@�L $�iQ��{���f㙛?�,��!�la�td'v^q1�̅_���s����Q"#�蒉�; ��O�8�U�m�)�ynsI��g�(4�;���H���� �Ǒ�ɽ��Ip�dE[�S;���9���(r���O���΍���zm�1ͶItD^$8A�`P�y��#�����1o_��P�޺*�Ŗz��`2;($��ssj�a�����:�����]�=8N-բ|�SD/��0�ϙ)h��Enƽ{�gf�5��Ɩ�M��c��l�)h���]$$�K'V�V.���>Ap~Y�m�����T�<�� w�o 4n�U��ɽ�c#*�1���:�N~��Qs[��C�Yf�� [z�t<���]�W_���=ܓ��e�c�ַe{}G�7����,�'-Ry��@�~jL����q;j�Mv�\/�}R66��¹������$�������Lۙ��@2W3wt�a��ϟ{���3V-�[��m Z��W��X�Cx�6Z�pg���Ӡ�5�\#x�$*��u���^����X\YT�z'�^E��E��W���#����(��"�L��Q(~B�"�YB�d8����|1�T���8��a�X�Goߖ7~��ɡ�zލ%^�>��^:��[���wߖ��
����;���]SR�:r�_�Fa{�qg=�
�ߗo}��ҥ
�/ɱ��k����'�j���X<��@l]�������Fl�s0P��a+����d�֫E,�&3 ����	��A�Ȋ��ͺ������W����
��ȷ���^��#��揩V�n�e2�Ȳ��G=��K���T$��&j �w܌eT�aR������IN�'������I�m
�4�q�j2�9?�9��Bu�TW�����������hRG_[�윒S�uɻ�2���v�	 !��z�ݸ!���fǀ�,��{k����h�I�,S1��b*�}3C;�"�0�e��2�:x[�/(0Ƚ[wl�MsB���֝�{�}C��@�͊�Ϳl��^�yD)w�Sұ@q��N��W����oȭ�cyow �iM�P�-� &D$��[��lq�����DWP���O��礱�%�ǒ�@Z�z�� `Y�؁�H����6W�&%�y_nL�u27#�ʜ�g"Y�ޥ�%��� 9��#)2�%ʃL��`Tޕ�a�����H��'?#�Á�w݈�'Zk�/�6������<�q3��L�݇�7�0�;7�2+0�y�&`�'r��h�,���XkX�s��囒���0��]�:l��E6,�h���	�

�憂u����	� Ƃ�(�h�P|������Ɉ��z�9~5W|��M���ySr�F�E�r��~�]YQෲ�"\���ʢ(����&]o��D�Z�E���W�K2R�>��ǐk��a�X�ÿ�s���ڇyj���G\P{�qt/��盋E��`�=?��0������Gzξ�"�:I�|�}9�M�ɧ^�uwYǄ��vM2�D6GC
9�`�L �Fd�8c�J�ͯ�����>��=X���(M��־`
�4z�n�o��/����{f�,��a�&-ÞG���r��4�@�2���.g�k��Fe��c*v���B��Ĉ��Ψ��-�S�B��ğ�\C#	y���q�,`!]Q,�1q�)�H?��j���.v!���0����-0r*b���P��?�#�}�����>��AQ5Ds"W�ίz*"����Pd��[��cB��O��ݱ���r�#���s� �Nw��5k�d�s�����]y�{PA���fJ�o��̱?�>r
$�1�P�<�MJð��d�{Z��f[���H��8��5c)���	�b��J��y(�0+l���۔A�>*�X��=}�% ,���̯����9 ��^��:(�N[D� <��k�˃{���i�\ݐ���ȕ�/����t�R{ �#}�·��)&�ˠ=6�e"����*�^~��]�����˯���_���짿���A/_��ڲ��Ej��:���\L<(�ְVa���K�=l�as�R�o X ��)R����Ѿ�at��	ʨ�ʂ(M��U8~�C>wχ���X� ^Ў]��{2E���Pt�*���vv���KMTi*8j`ӆME����p�76�2-j�ǲ��)�ژ�k8D�b���j�Ԣ����K�	���
�p��c����O��3	��%5�0��\?�Ic;F!�ڲ�&����e�&��0�� ˊШs��M�dj(1�	J��:1a��]O��aޛ����l��2:@���ڿ���H��a!�8���a\�
8������p �FC�z�2�E�����ޞ��lRV4U��(@zr㌴g"��.󗆨�yi�FW���0L07�H�[�f�qs]�Qѷn�C��f_�:�'����n�Q�� *'�ӯZBp���"�FDC������Oɨ�@0Ԙ��۴µ�!C��Yo(�jX�_q�5
wV�-���ʑ��=�O�5+`�r'��juF��}ee�{x�����'���sr�w(�=�f �
_�8.z�mQ���h0*Q�j����<J�)�,�Z��	�-!|�ä��&����Z~�?�O���r�J?��ޖs�,Bg�8-� ��s���T_�kvZK4��v�ʧ>+���D~���Z�]Z����!c%�G�S�/����]���2?yv�YTR�k�x��ȟ ��Fڦ-i�l���@�.5xm� ���<��p����O�NAT3�PEVtv,����7�����z�%�G}��"�uc0Vÿ�ͣ������`�ѣ����Q�K�����٫���}ԎlJΪ�ꡮ�xZ����͎�K��	��*��7��Jo��X^��DF
\�!"i������u��\���T֐[�����s��/�(���gl� Z�h]�0X��8��6�1ͨ�^��+(�X�R��П:uJ�7�����uy��:��=�r���\�x��>Gȗ�͡� ;�!�T�[\	�q.����W�Rݘ��ݙ�����.˃�
�WZ2�1g��W~�sֱ|����G��5+�Ԇ������#�k)D��Ο��%�8[��:hF0����0A\#Z�ߩ���[?̋�؂���{1�
y�&f�M��I�e�<��#+��bwp�U�[��Lq!�"�-X4�46\�"�\�ԾOEG�ȃ�;2�����EܼF��`�ӆ	�-~o ���g4��j�'qTDI��#��j�c��� ����
5��x��1ђ����N��B,ߑr�J�okJ����i<������'�B]BR�'/X��Q���#dyTڪt4&f��g.=k8*��8�/1�0�'j7���V;o�ۥ�iX�u���des���m�H1Dd�υ�:�0&t��^#��1B�Iy�A�t�VA��VUl�,f�7H��@a�|1"v'3�����H���.ˋ9#Qh��]��&r��ȁ�c�$u���� �ָ�E�Le{6��w��72���'�#�ԓ��Ӻ��wץ���]�n�d�(����-�su^��z�}����������l�S[��}I������7�bj̓�������>�i7�~su���t6Ғb�U!DV�׼��(��#�z�[x���WD�s�'OPv���Ž�0D
���X �Š�\�
�Oz�#��AA%���;�Q�ޚ+8��re�<{��\�pI����$�A�����������t8�����!$b����w�jt�+�?ړ���?�.�j� ���H�|��K��'�UX���M	�����=y���(~c@�V��	�^",A�vf��	h��Q �޺sS����Fre�	���>)�_|��(��$���at_��f�D��l�?����m����_����r��2��ˉ��-�Hu����|�rq}[f�>rASSD/S��fѝ:O"&dޛ噫���]���,�ч��/�oK��K���]��j.�YD~Ց�a�W`>��TG� �M����=!���7�Z2=N���h��pN՚����5H�Ԑo˅SgekkCn=x(�����wf�3�>0s]�� �QQ,2xf�"܃D�������,p齡6J�PK"51����Y?p���F.�@5N
� ��r1�&=g],^���j6j2W`�z��l<���[�r��2hu�Z=A�1+R��Z��,�l(�X�	R�ZL�o�MYn.�{�\����(Q��}QF�˗����> ��"e�)�D���e��Q0�2̱�k(`�;��g��{X-XfAU1'V���h���S��7Dm!m�I����X�"�-�X�hڧS�հڟ��@������پ�/����ҏ��'����wab���GK]X ��l,W�$,��ސ�����x��%^j��ֺ�-}���v1G�gOAk;�r��K��X�f�M<o#����]�98v�1�F��m����������������e �N��3������{���C�H��k�� �X�ݻi����<r�Z:��G�LaT����D	�9 ��/��8?� ��]D":��a�|ꩧH!E��� � AY���\�&�d=ΠX�p����-C4ǾP����hF�Q��?׶E���=�P1�~�\�׹Oq��h��>�H4�iQާ���h^�P�g�p�5#��ᵥU�jΤә�F$���뫝xޏ�p�#
>k�XJ���Nf�S�W��؋��i�xQ`�A�����j�L
BśK�����Y�R���������y�q�Jȹ̳�&y�
��x��'~��ֹ�5#�q��a+$b9����Ԕ���������q<��QT8y�p���$�*�9e����`�~�/��3h��-�����цL��)R&%�6�hs^7� {XU��A��b��$
;�i8��*}8�r�?��`��R̯(��EVRc��t"����^bώ:֑;��r��w*!���6r�ԥN�d�^�9�X�2SDE�QI#/�I�)B�� ��⎏P�ݯi1Sw�=�fv�g�Ӣ_�c�N
��1Hd`6P��C~��#�}���&0(�ؓg�#�*�?���9}��\8s�^�K�n�Q>!�-���] 'lE�#�������h�څ9��_�;?c�b�{�Ȉ����2�}�?��\{�:uKN�;M@���ڼѩ�Q�g.h�Z�)ז �!���d2a���P�JI���w|(�C��|�my���;�����X���5�;2_����M�Yp�^��۠�	�(�%�v��Q�ɽ5���{�[������/�[YRu)��Z���3E�9�|q��\�ɗ��hąf�[���
��j`�3���nm�������;jH6e�dͨ�t��Ύ|��eC���ܞ6s����HH���"�4|.���-�PN��5����+�sO|�� ���'35F�{�|�+rnsGƈF%s�P�`Ɩ��X�2?J
.. �P�	F�,8��Ȥ���T`ъ�#@?:8�%��^_ڈ i��ڒji��uq��z}���A��֍v�M^+�PҀ�m%>�)=t�����F@� (�Om_���~!!�Ӫ�V��w�OV,�V���m�I��5�2o��}��X�-�ߝ�L}9u��2�7d�84ը�#���<#O$&�U�rJ���t8��W����'��U�O���&]��g3��$&f+b�c�s�>���5��=����΋�?/��}9���JOzy�c��r�Ď���d&Ar�rM�9�(�IC� ��xF��:)����}$��O����XV0< �������o�� [c�����tPtL�\���h��qw��S�uI�����Q6ַ������X�I�p���o��^�3#��&m<��/+�n�rt��W��<E,�/����]D�Q� 6�G5̱��@��	��{FF��� ��"�pT|p����}�9e��%(ŸC��P !�G��wﾎmK�7��[�7���\�Hz0`��,Y!��k���۲�?�N����XA,�c��Ԕ��5ё<��NPkB;��6o�)�Gu�޻wO.]�(����;�󠪋<���s���E�\�� �p�pT���%�q��R쇊��h$"�����ac����|�k;@��#F� �1p��� b�HL��b�3��c�>TE�`�
?=Qv���E�w������߱ge�Մ3Sd�;�5���_e��-�B�Z�1fS��GدrS]
��F_�����hH�t��a����k�Α�7�*�`a���?�A��i��o���;QK	�J��=w63UI���9Eq@���H�?�.���x4�1����:f�"�{���Z��KꥩP���b$ ����P}5��̣>�KcI,�C0�<+����`��QO�H��ɑ��q�k�����QV�׬��iF-)y�~Y�6R�a^b�q(�=��5��l�2�*[&��4	v������s'�R#Z�ĺ��(�ON<Y5á��w(/SUw6ϋh����X�Rl�4�;�	J'������+Jɐ
�`_ �+�����ʝf��mi�R�l|���ʿ� �/�otX����En!�8kch��P
�L��jV*�����a\��B���a�)�N` �z=�����j�A��������k���&�N��'�?s��p�̵	�Iѡ�[��iq^��%�%�æP�w��pܓ�ϙ�C��P�GGLw��=��x��g�H�����3���mYQ�0J�8������.R��ڿa��"׀-�>�w��>�Q�����"��8���ƅ�dy�bC(f�����gիcM�R#ь�Q�q�eE�P+�<g�NC;b�ޒ%�o(��15��$k����c�$�e��'�r�2��a4A�p ���op��\?�<)4:���T7��eGESK���%��ߺ����X�Ԗd��$e
|f
D�����􅜸�lZlؤ���7�LF��%̻��9�%DϬmr��|0R@<�N� ����;�{�}�lv��L'6Gf�1 �=�y$��{�E�I#�°DԮ?V�lP�_�љ�{�������[à�NΖȵ�}��W�%�I.k @z�.�f)��hC�\0n�P�|J1w�0\��%
&a��u�<Wv�+XYU]?7�2j��$%".�«%rb���V��B �r�:F1yTCT�'k�˲�@cF�7�� e�!�vG��D��Xuqx��m9����e %�Z��m�"Y�gI�u��:��躑�je4�r�~_�ړ55����'���|p����%���X���c��tjϓ�>?����-8X��,��4m�.&j�A @���:ā���Uio��EO=��,q�2� ȫ�� Ď�=�T�^ѱ��مx������ᡂ˶�ú<���,���g��7r�<��]�$P`��(7��X�͌�m��+h �meiE�鄑�:(��X��_���^���&^�`�r_󗲦����ϲ���=D� �<�(� M���(�Rp�·[:u��\A�?�j;Bp&_�9{��n��m�����:^�l-�
�ޠ��R��3�iA9=$MP�Y�1e�q���緶��G�ZY^!��ڵk���)�>!�������)�T�	��p��&hd�k ~P+f�G�X	) ����f]B�Xю�S9Y��H1�F������Q�mw�A��>�=�����=V ��EqL0 rD~��iIA��E����� �P��fSǼ��sP�u����W��wߕ��G��ܻce@��:�w��p� ���D�j�L��cL-on�s���m�/m�e��ZC���+[�����TIi����6���?� �I�V> ޹�֙)�j��D�E����W,O,x�M�%��hN�w�yq���v�:o���E��DC���k;�9�6RJ��gBM�*x�QX-�N�rlQȘ��~�(��uU��ֆ�a 98Laq0;p��C~��o�:�[[:*�}��[�k�,����.\�ӤJ�>'`�4���FB�j�G��y�^��J�$V�)~����E�` l.�YK��eR��'K�f{�=�-K© A�G�sQ[{;��i�6v�
�1`�!���pebT�t	x1�����Nt�	���3����'�fD��S[��� Us}��v�G1�
�s1���� �����<=HQq�ʍ�u��M��+����>%�=)�wN�]ӵ�@l@���<Zl�f���bvG�U��Ҏ��G�};E9
�Q���n����s`@��6�����/���=E��Y���:�M�m�	S�a8!*�3A?�!�����T���+��X	��=z"O��m��Ӱq��$��*�[-;�1e���Bb���4� =9���lYA�g5�3 ���g�������i=��L�P��5
|���/~�7��L�.So�N���"�y<;+��h(G�B��ϋZ] 0  �� :�s�%$�G#5�u�}p�oޗ�H���l��ʑ��}>�8�hLBD�Q<D`Dv���P}cn9� rmH�4�K���_��Wd��Y�R��b4soˆ�ٻ/��/�\�=TC2g�o��G;�D��Yk�虝+�E�xJ�;�
phd (�ޥ�%�vd�̽f�Ct$����֣�r��}����=�{0�����՝��LHN��jXQC ]�P�Q�2:�S+O(�~�zc��-
��6�g�Ngj.q�BH�H��q����'d`e�ߣ�χ�6!�0x�F=y08�;
�z�MyX�ʱ���2�w]<����کK���s���M�+��i
cP�f��P�����p�<q����&���cK�1�~u1�IYs֧�j4v��T��*�mv�4��3�x������!W�P4���x4`�&���3��|��ݓ;���xM{�5�-caF��D�n߹#�[��^]��z!v&����Y�ͬ�mͮ��X6�9���?�ө�kq]�|C��냍������q�j7H�D.�t�����&3@'�;k#��5u��⓳fԜ�,X�( އ���󽽇R�V@e�`α\o�b=�C5���d:P�֣�=ٝu�MY��t�oj�������T�18��A��tۉ4 �Z�tJ��U٣�4jh,��Qh�]�5M%���� �w�@ń�5�<�_�.��k:�v�_�"KA`��&�P�/�s�����'���!�KQ/�U
'&2�(X��{ ��sO�*
`�k�S��8��8��@ޫ��P��dt�$�5�Ɇ1�M�W ���
})�-+���h�}:3�w���|���{�~I�����.�بe	�T�o�^4�1.�őѽuq9�:�&�'��6����[��gW�}����bd䮄���|!������?~�u��.� ��|��i�Q\��`?�X�ef#o>1ᛂ�F�!D
^:(�o���ċ���F=m�X�G~��q��B�qn�E.S�9�,
'�.�U�� �G��p���{a�KP.Y1�x�(#�Z�/�Y�� `^F�~����|~pN�r* /���muZٍ����mne�\o*%�x6:�"��Rlu6#�G�w <���p?E��#����r�R
��}~lqN�t=���E�,��ZXr$6�z:�xl����Cs�;��4�<�e��T��L�����-v�ʸNՑ��Lw�!B������X[�c��� ADi����򨄠�ׯ����Sj�M�<DK��l
1ɉ\�z�e&._zN.��(��_���uPב5��UW��9Kak���f��Ǒ�C�mK�NЃ�}>�*(����{�z?�,���,\�)K�-9��Y�4����}<�]{9�,�8/�N��P��X�4��(�<3np��.IB��5A��J�HpX�W����wW ��(��ma@�^h\����8�]^>cm����N�N^5�3�ԇ2�+ �W7Vx��O��E>s
l	����`wL�����rsz��s:��G�>=��
��_Ѿ<w�l�Q�(�C�V"�G�`.��~��s�'�9Jt��涢�&s;j�յ��9#O�;�z����߽W�p�����	 (�ATd� n��P#<׿(�=/�ⷤ��KR�քB6=B��,;����'��[
J��P��A[ȓ��@p���َYF�ѱAH�2�	�tp��I�̭j5��<�{:��5u&i���\:q�u��]Z^�T�?<��E�
u0���u�θ���H��.�Y#3G�N�v>e������l �kf8�  1J	檫^��Q?~QIb>�+;i�&�.�ӾL�TΩq��l3��9s#.���5���׶�h�-L���&,%cy�3x} � �� ���BW[���B��������}�����*0�8	�'�-��k�Ќ�a	�gϗ�HK}��X�9֥�#
�ң���h�gt� W����#���\���oʡ������I4uY�*�M�]$Vt8x|�M���Y�H
J2*p����=�յU�Uc�
1�#���F��<��
�mF�r����h��L"}]|�����E�O����<��d��.�y���Nu����cm(��۩���*�#���[��C�g���ˋ������>���@$���j	#~#����P�X�GS��{$���2W`G:Ol>0 ��Ա�I�R�N?2%�&FTD@W*h-�S�h�f��:�,�ש)m��+����<��`�TݼyC��7���c����>+���/x���yi�bU��jb�N~���\#�LZ�;��@?�u� ux�Y�
�_����P[1 �j�0�q�_G����J�g�l��$�T*}|��	�޸����@ׁ��c�נXD��ڊ��9�͜�dŔ��*�᠊��L��"����Cy��7u�7%ܕ�>��J�ӷټ��V�����9�^����4���r���@�����a����,�`�K(\T	QJ��nn�6��M/��`D���U 	� ���������S�DM</���I���x���>u�kF�FI��s�l��(�F^F�o�.�eh��-O=��EѮqi�������ljѣ9�hL&������1�f�O�cnT��Jq��������<]Ⱥ+��ɖ+�?��%X_)��Fŉo| �H���C�-��.����&#ѱ	.��I���F��N��<�b�*;l�^a�ňX0��hxb�cq���➫��W���c��9��' Yn��h@��5RW@�����F�#vR�-�@���UfG�	~b�l�L�{X���ʣ{���i9����>-˝�V��u�`W�ಭ|��Y[96��yνcgm?�a=��d%؇�v (=88�����)k}���r��]Y�\e}D�_��b��^��V�eAT�ڿ����GU�8�~���������%�S��|al��&a݊����w�/b��{�iuc��@���vb�4�����x�9}9#n�ĕ�@�Q���k�^˛a}� u혶��ѸYD����\6��lD�
��(]1�[�2�T;��"4��^|�i���%��&��ɒ|��O�f��|�H;5�� �tsm]>��>-�km�����g}���7!H�o�ޑ;�C���?r��QA��G���Н���g^I�?z�c����@���x�����벽�E��\��H��b�,ѫ�A�6�X_'� �_�w01"�$�w�p_��K�."x��h��h�a���@4�,zC� b D������H��:=/X$g(Ƞ�
pi<<8�a�Ծ]���	�?��U����J��{Z�>x�@�A�fO�ɱwپ�-7�ǻҝ�X�[Y�u9s�SƱ7����Y��#����G$^��(�:H���.�B�f�P�hnY}Q���Z�v�q& �2�ꂲ,[��-l"Z?;u�h9�#!����O����I3jR�fs]�{��������Ç��;o����eY������"���'͑�Y'P'��Ո�B�#�f��#'7�6x�VWV9N�ww�H �l��Rb@����<�<��ĘL�r^8�RI���t�Q/�s�1*����.#����H{�+/��3���h�]H½͇��J^�v���?gC��������s�ݺ)����eymYǻEL�lm�SO]"��6��F�ž��d00�
ZMck�����k�_AɎYL�y<�D�s��z���o�cj���}�'8>�u�<�d*^��E�Ҳu��"+���ߦ���1��o((Dn�֩m��W�J��͛7	���'��|��K�6>�R[&U�0�#�inL�	�����6#�P;���{�gxnn������xJ�o�� �s�K@؃
/7�)Aռ<G�������Iq�We���)o��颬��%����=#�z�������>��
w	׃�fG�G=�[j:|;����<�w��Rx���0���m�C�bQY61�U�E��'�J}��%���V�������^d��
��쒋rĞ�o�F'#���E��kzQ
�����XX�}��Ŧ�Q�H�|���U�j����$6�f�q�&AA����)O��@G���GqA��x�����Q��M��3���z��,_��ܣ]�����PټH�L�d5\�pS��k �:�H��yي�2io�,���h��,���p�L�!*�zw`-��<� CN�G��;��A��c�����Os�_E4�)X��^�9F��{繫�V��a4��C�q��<��fr鎉}�X�%t����\�����q����)��:��\p����	 ��������P�<{ENmnQ�!��sBv�֑�J=�R����J�6>|j�-��`V���hO7�K;([q�C��H.?��d����p�����q�j�v�;L��m�x�*�y`c��. ¨�y�-�W>����x�H1�r٬b���E�><���D�3�W<�坅1�f$�����N�؃��in5[,��&j{�FLP�P^"n8<�{?��-��j�vdgm�Ԩ�B�`n"�������P�}P�G2>��K���GG�f��<S0��`(?xԗyoHሮv�׿�y�+r��-�����]5V���ߓ����C5��ݾ��I�Ӗ�{2z�uy*,"�z�"��|3��9�%}�}���!� �Mm��>*d�W��#7/��s����\��,��ŵaX<s�����ͫ���o�����E�������?��)�d�l���g������D�K��\o-�����a�A����]��0�u����P#�#}5���R %���Fc֑;V�t<,���P�����!bΞq%��2�S���(ٖ�hsO��n.�G�2� ��1���`�<V,\j|��Qi�@�D�EH+���3!�9�'���ӫT��C�c�P#8:��Ohc|��ʤ/ݕ���������lj?l)8ot�XԾ�ͅ�G�l��N�y|x��Q�ʛx�t�6�����ᑜ�pVN�;+�NC޺�,/���ܑ;:^Q�u4ۈ��VI� �R��"M���q5L�`��Hn��bP��P�]�mO�ӧO���,���J���E"-tQ! [g���)���ͼ��_��m3W�������#�灓��OQˮV�R�����2�>�
�9#o_�*��k,�����X���@v���v�k�!�Q> Bԁ�pèqSO��^��d7��@��D.�:���#�U���1��
��C�^L�l��Ї�8�+dex�L��'>�R���)Ho)0E�#�u�޿��4;-�I��P �R8x�Pf�#��a��niR
��r�/OX�d��;gy��9��|�c#ӵ�� ��:��� �Ss�"�� �:�ϥ
��Ɠ�^���b������Bu��0�S��W�����^�\�Vx���]��O^�wJԖg���3S��Vx>1�41��Cw�N�Y�����>�y��@�+��~���1W��<��D���Q)���e[��⾄��e�f�y���Y�[��Jd���m:��ݩP���^�?q��c���]�f~�Bh������ /�Q��X0UTq���n��3.�!����&�ڿG Q�P��������|q��K�6�
Z{�dI@��YphT@�[�MW����bu��{�r����OZ|?�A[��jc[[~`���Pv��H��>�����'N3�9�@)6pFC8E��΄�֡Z �K!zZ���W\"yɆ������Fx��/�nl]a��I�v�{+h����F�;1�~�x>�rx\t0�N�^���~~K!>��Β�8{ܸ��	v.���%�L��j�=<� �v�^oֱ�[m���y��m��y�0�t�{l�X�ͮ<q�<�L�4���/�Ѿ���,��u}/fD��"�<�B�$
�ꘓ���Ƿr9�\:�����H
ޅh�m�F"�
���=��ɒ	��I��^�A�\�
���˙�XBTŢV�)R�����a b��9�H�g�?)W.]f�ŹSOH;���| ���oJg�
�n]}_��C�,P2�����xN��:xc�KJ�[���`ϻ����s�?"Vm�����~�K�Tk������y��59��&� 
 �?5&@̈́�
 �?Q���r�����xC֘諛�xƨ��]�P�~uyK�W��TsEz������,���\VWےז�g{������H��� a�3�>PQ�M�QK�����X���ߐ��Sl����$ek{��Ͼ��h8��Z��҆��r��sJM�.��4�yx�Ϩ-��H��i����uXI7/O���&t���t,�RM�6�}�Ӛ�浌Ea�l�نx��}����T���D���< �%�&�ǤC��dmaNC6�%Bat��u���Ql�� ����K��sr��+��<s�{�o�Xo��
�Hփ�߃��Y_V�n��ⶬ}����pГ��g��)����ʪ4G}�9�-�Ѝ�%���tԺ ��A�����%W�<o�;�#�c�su_��z���&����؁�̋��P���<�r�9��iQ���`|�=��M�&'G
�#�P�3%-o�\��6���M� �����>����'RSp�z��l$y��3z �$>�� *C����ht��b�U�"0�m�hf���}m�d�4a|�q51�VVn:�Ԕ�}��8��� #��rI�-�g&
C�Ff�탇emc]��ש�<̆T����d~��!0����8��	��{��Cc{!�V��ERD��\���u�L����۷e��C�DA%�� �/u�kP�D��{�:*"�X��=�Mz����(GG�
�j�e�C�`�fF-�� �G@��x$?z�y��oL�	ʉ�#�{A��)E����A� PS�
$M˹��t��c��{1Y�F��3������s���w�,DHC�"s#6�XaO@ȶt�PG.�E.�"f���f֜<p�Y��~����ϓ�/H�ͤ�B�7 U�9	����Y�	�**{f[ �P��2bt98h���:p�}#	r���"Rf��RA�"�ܗ���l�a�ʘ�Aa�>L �y���BIK���`��yh�
 �C���A��[�����SK�t)xdx:���2c�U�9��Ϗ1`to	�׿���U�`���kf꺮s|��$O�9-On�(�j���������=�3��&Sh�5�rO'a�?%l�~��s�6��9�\��A����{<jGChmyu�����([1wO������u<v@�Ԟ��J��ݗ�[�	PQ[��	�`��/�N8�jd,�犼�"�HL�^ʨ��*�� �� ((\wKCm�U�A!�)ϝ:���1�����wJ��j��P�`N!�	��w���H(;���y���(4�ўO�T6��Ɠ��U�S��'fw�H���5+�8L&��U�3a��~Oq�x&,����xm���0�rMS�y�w2�Hd�h/��dq&�T.�QY׍��t�L�#u�n/���Ɩ�Kr�h_�C���j�dueY=x$/����X��70lq/�vf�����*�����^ِ��?G}/� �"�E�@��PSL��'w�ȅ�Sz
��ܟg}_���Z��� 2����
�l��~2@Ã��X0x� "�r���
�p�Ο='��6���������X�mIe?u�]������DXk����4�@��~yV��\�j��ˁ�C��00�P�bD��T�=�Kj"T_��' ���N�����;zگ�9�}���`h�S��5�zёW��O����U'���Q�W3+y��K_Cv�^�$��EO615���C{u�����r/G�0���̅���t� ���dIa������zq��6��v���L�c�L��q���(z2#U�j�	`��bM;�|�<Ơ���z��C{E�=�>��a��#�����H���ґ�����|^F��6����
ۄ�F�P��*/�ކ|@Q���=y�;���)`� =-r0��c�r�]��� m#�(��PHJ)����[��<�L��['E��{�{)KMg>������=6�1,~.TAͩ���r��<�Yk�QSg�{5'�9޸Nd9��$c�MA	��k!�7s�昉���hA��z��6�˟�Y,�� QTD� \����
O4�g�~���|v��e��W�Jp�����΄P�7HPg&Єv4�W��VJџ�D�q����L^|�E��w��W����JR�zE�X_��*�h�������!"��'�3�y&'<��w)i��J��{�?x���A�5r��[�rڞ�{Uޅ@�`*5�dI���"�j:N	m�s�������P�V��܈ kN�J6Ii��x��
�ͨl��8�Pr&DO�7�*M+��r����Z�9��?O�W��G�"cf�%���ȸ5�Z!�ww�%%p*�b8�}V�'��Ru�Wd���¹�D�y`�.�3SW6����{g�u��TF����Ο�gxGy^�����������}6DJC�>ԁ�FA�ςZ;/=�����%��/����xTت���?Zao�(7?�-w��5���J���y 9SFH���ʑ��GƋ�|�d��ӟZ_�+g����<�V�14��~:�^���"tjR%�ȁ]��Izf��x�C#�����ǚ;��9M��r�`��>e��n߿G�F�SN��"	�7;hG����w�u����֎�.��
�.O3�����.�-�����@r���!��n�e��p�M��?��V� ��Pw�~ 5�3g�`�](v�y�bY]���J[���`����斵�|&]�̧cT��b�a�V}�&��]\�ʢ�p�%����{Yi7d����S���ǁ?�b!�0�U8� �q5�ї�tf�4q~5���y��'����Hh9�T����m!��Ga`�h�S(���4@P<S5���O��s/�;o_�
�qMHӓ	#p��	x �f�I,ތ�
��-(Y��ǜ<]\�(ȵPA����K�(��}��5�D޿q�|���rk`���@daN�� ����=��6(� ,`
�h:�3D���K����eELD$���:��r�
��R�>������܋VV�(X3�[���d�	�	IP� � ��1�V�%���b�	VBDwfz���1�bU���YRK�Z� ~�"�4G={�GmGm�N�j��ܢE��Tf�)�U���p濇��3�=D���G�֠��A���%^ڽ�T��X��d�I�&��Ca�>B�*A� J[��$���<70�=�@���k_��Ȝ &6FM����`9�*""�I��_�H���L?3aQ���kV�Kl�"��w<ؗ;�=N���u�+D��`��c�:�ƺA�}������T�@8b+2OU�Ȣ�T��>�n�Q�0�0���>Yݾ��\L-R*^L܀���"����\NފC��N06��s�[���쀴�p6X3�����qD��h_�������J������Y�tq�iH���$�It�Y����7�h�X�����$N�Y�L���H�]����Z[^zr��|a���P�DG"�uz�'�a���@7N8+P�  �8�&�� �p��%����}FѶ���
�m�]w:m�<- �4"�	� s��,#�b�i-����lmIO�\�5��uq�Al	/\�� ��"P��6@i�7�'k~��Nɣ��K�Q J�ޠ�'L�L-ꩳt4:���y[^~��G�Y�k.�9��r}�́FzoS�5����h ���8{��t�4v����`Q@���^i�EY(�'1�=l��������P�����L��8T� fC>���RQ3u�`F�8�5����¬ǯ03�" ���$
0���J�L�B�hTp�4���q�HB~\\^+�_w�Z�7� ����܃�A�	Z�k�?Q�ۘ��hh��r5 o����T��> iIaĞ��EW{��,e6�G�5��y����d���K��4�c�n�6	5�Ά���X/���vW6�^�z��N�H��_��V�б�B:�GP	R��-�D�@��<5�q�Ȭ�Q�X^c� 3*�c�荶u
٤n� tÜ�_Y������i����GZYWȃFũ�E���2�=��#ڜ6?urփNt�~ㆬ�M��`H�ބ{�m�6#}:7'ә�1�Rpj�����߅�\�H8:��	s	i�1-��=i8`�Ԥ.���d�Ԏ\�x��4q; �Q�O�����țC��6
��)��D���U�ϣ껏9N6���qoG8G��N E�>vYʃ�X�eM��n~�ۙ�\+2i���H�l����h�9 �����Ċ֛�pX{�#	�'��n0ܠ���6(���"WD��HFqC.�%�6�?ɧ>�IY�ܠ8ǹ���o˗��Ez �y�i��w�F����\�8uZ���꿖����X�d<�SX���S=�$eg0����' r�&��a�'�Ԩ���+���פ��>H�V?�D�&E�D:53L�����H,GQ�.���'6��i5���mi'-��0ѓeP=si�-�޽�46����8�[��ܗ�(.>�U�ח;��*�^�~�{�}�y��I�֦1��K/QHap|$�j�u�m��B5�*B�ť�(+[��$fuI��)j������T�4����ov���J��PTkJ�, �#F�/� ' jc��3Vz�c)��żd '7�(�R��ܮ���"I�,!�5�DpSp�9D�F��B1(w!�fI�N%��n�zzs���u�@e���͌Ҕ����e榔�P��N��@K��D1U��"؄��P�-j�,�W�()/V�QoQ&��%_3�׀�N��hXb���A�3/z��g.ܓ���@�b0��p�L+*WDD�8A`�V֑YF'��Z7³�IŦgb6��[M���a�#I錁r��R*�O"�5��oI^�3'�s�B�{n��o�_ӱP���0ll,�ɀ>Φ�����`P��m+U�Q
 ̈V�[�t���i���1�)*s� � ��#q�U���x��͛��#�۟��ʟ�ٟɻﾻ �`�����V�ޜy��8�פ�8�q� �:m`*g�=�c�c}u�τ� ��5���GQ��/�g�|� �9~�ͪ�^ܺJ����̜��PFjj��L��4��Fr��������{���Sm�&����Z&$N��kfb#���h��f2�99)�xGQd�x��m]�(�<G{��Ib9�y0xy�!��s��*��SR�����YN#�E�FP�] ����L��pv�{���|H��(��q.��$0��DE
�� ��q�] �����3r�
���p��.Cޟ�,ҫ��� &���C e����j�F%����^���Ւ�M/@"_�)���2��i�e ���)�`��!�ЕF�!�4�'�����zi(����ǚ��E�]Vm.��6��>�"�",6ez�b�9EBK��k���S:8��`υ����~�]ښ����#�=�F��Vk�:��Y4�Z�W�l����ظ�_��,�����-?m�q���~�ٱ�"
�e���M�Y��(ϖ{[��Ǡ�_�X`�To��')A��P�][۰RuKI���ܮ�>��W����;��mkk+�?�/�ý����ܜ㰟�9�`=s� 7�`�P1C�����Oȱ��&]ȉ/�E���r�p<��yhHe���t��R�-���U��܄�!�{bk[���SG,O'M(
h��05C�`L�Fs���LV۽>q\I#�$Z��Y|���$M�Gߌm�k��RWM�#���0:23�m9��BC��� ׎�Zd�BzǼTt�NG�V��rb�V2D?�V� x�������c��?�����e!���ʿ�w�� �uG�G����J3�#�!��h�������K����\]���/���"O�;/�h���֐��z4��X��3���>�����"߈$@Uq<
��ݤ���%�٥9#�ʜk�>ei���{�[B��?ҘGd�����l7����1�q��+r��=y��S��˯�[����x����˛o�.�F�"��hlo2���c�u�C�����U�H�Y:a�	�5DB�W.*�cW�e5��QΣ[MƮ�V���_8Ǔ�ca�t�b�A�5��"6�5�J��"+��eb�"�WZR�(����{�.I��Z�DDΙ5u�<���H��H)����(�=�˲-˟�I?������zK�=���GQER� c�ntwUu�Y�s�����Y�N�E%V���2##n�{����OO�|8e��E�ٛ�ɎZ��D�(��֟-Dݐ�BAĶ���t}�
4��42R��� �ބRfΰv@OŽ�`��!� ���,KNAD@A���D���K�
�[�7ݤ%kj̨���Z�d�KTh�Wa�m��'J����4ʴM�I�	<T��{$�6&�j�)ԙ�чaE��̩e��"hPs)�g�����k��B�5���pA���HĜԿ�u[x5�97R��b@�jJF�1k1qPӝ�c2�����؎N�^��>���e4I��l���� �v�F e�]�g��e:�p]G��2��E�.��C5�< �k5n:�Ӵ�[+��D1�uagA�w��.]��<���ZB�`� �=�����_f&`�$~gt5���C����!r��{-����/�&Tݸ�D��x�8�e�-�BD�	�f�װ	G�g����G8�s����"(�B-Θ!�]�@�eoWn���|�[ߔ��|SF�`*�z�u�V䈨��իk���)�"8�Lja*��(Q���:�:�w1+!Fk�cSc���d��)��?=�pE���?��$�P�H#%ۇӸYE�C�Mߝ�P��r�l�㩡��J���"0�:�@�9{ V�?:G��D�@�)?�9>"?"����٭lj�]�y����>wvl�O��1�O�.��{򕉴���a��_�/<(�TT�Y�x0���bSL�L��=5�"+$����g����(M]M�k��Uq|�D��/��y��9.�bv���g��P�ƻI�D�%:gޫ:ސV��$~cL�$��>����e���ZDb�ŏ�J"?�T�����
h���4P�*Y����
=������o�%� w����L��vY)}�q>>��0����3g�2����ĕ��~�^�J &d��.��� ����x(
�a:���`�̥�W.�\�ʮZ��!�#�1��l#��W�x]~��������M���1""T�pGc$k._L'�e��xj�W�OU�=�������Ĥ�qCq!�7��8��I��PU�r�	At��x2��8�h�%Q,�M�͢	i�\\~��|B�	��
\��EJ ț�z�LǤA��1x2(�dO�f������f�g�yV������|�&����/�����?�/�@���`'-� �j�F�Ǔ�s�����N2���t��dU�� �|����y�p֠xW͑'M�� ,��
���)��F��<�F��U�S�v�(%�x��oZ$~���J��К��y��Ύ|�ߒ�:�O<vM^��w�KWY�6�y�+�]e?�v���?2I��#b�j��}C�L�C����
��.�C'�~H�7���IuՄ�������A��rƺ��8g����D��jk�L�� �m�=}�

��z&��AݑAx5:��g���Y�ě�&&�a�Q�:ʇ�oQ�8�e�;�����!S�йl001�b�������>)׮=.yǮF��q��A�t8�tr�%�&Q�{1OmM�6�(mM@��7�#M�v���d��sP��:F!u�7�^�"u�2RwqmhO*,�-ւLY3&b��'�?%�����2SM�e4���äs������)'zd������7d/�ڤ9�������/�)tg^g���6�Y:��.�=���l�"]���YO�:�=��_����Ͼ(IÚ��u�BЧ���z8A���^c�k�P�ԂE�����S�Q��&述��{8�;��A&��@-Y��r�GY�Q��S0MQ��s�^%�����iae�W�����ڮ������1�o���/ 6x���^z���( %�*~�b.����+� fc,�������*��1j���~����^�+��@`!�����L��c�u徵 V2�\q��p&�Q�ՙ'�c�;���!���7��|_��Nk2B������![cX�����e�Q�T�U�'�;�;�1�3�*�"ѵ��s����J	0(�L�j~�\;��E2�W���E�_	/���}�ʛY%ŀ����N�I�R��gE��Z\�p:��g�\x&6yE�κ`:PW9a���c�{y�ޙ!���uUcav���E�E�91>6�כ�������:y�B1�	�Y1\sa�e(���x���zꕍ%B��V��;y'����sL��W�Ģ:�G�ࣨ��:3�����
����Nb���G��������'	8��D;�o�7��% �%�Z��ۃ|�X$'�TYoT�W>y8�$�0g��#���L�)��#���p0X�9q���s���`R�t+�0{ײ���)�O����C�*�
�%\Y^���>i�UpM[�po��Q#[���#zwc��22S�-�(�R����Ӽ��=̮R|*X@s$�xe�]^�Ώ����j�P���(sif���A��9E����Lc�K��Z�G��^5Q����<?�1E��ibI�/�f�̯�b��2bTn2�l�H��-̃msQ4K�2e��'+�MD�|��b͚�F��՜԰�Q�Iju���Z�I���V��,��dD�kpЗ��g���\�����s^�YS����US��Υ��nșsg��ݻ�� @��AQeQ����59��e�7e52
ǣcfSRd������b�k�n�O���{`c5x���鸢�4@�3x�3�dc8�1ޯ�����k�c��o~N>����o��o�)/��:L{��^�ٰ|iu��5 �z�F�]�( >V��j(wЗ�z� �޻sWv��=a �	�ҁB�T�M� ]d(" \� +)������&�C"Z�:��R�6 b}��,?{EjKM3�2J�~©���.b��v�E�'�aj^{F�M!p�Y�Y3�%��㷣�}Y��dP/ȻG��	�
�g$ԧtޠv/���.�S��t�*X@f�fd4�$R8�.XX3�Z���(����$�*8�ȼe��O+
��lb���YE���>ss����[1f�H�Л���˙K87����!�u���	̡���#֋Q��\�W\���ny�����ڢ��� �cM���U� �R4u<Q8A�|Ȍ�H�7�ĊURY=�./��:M/�ӑ���1�9���Vw���[���Ɂ"��/Q��<�Ya���`,��)��#��ە>Z7�5���9�B��XoB��I1W��M9pN��G�5�b �in�(z���������v���3����ݺu�^gd
��������W�ʟ�k�� jGfZ b\	΢3KlC��.�3x�&LG�	�m`���Ei ]��$82���0ԓ���I�'F-�swl��������oD��ĸ��o�j�3d5��6I�{�߼+�忖��C} �'�R]�{,�
�1�]�W�~��E���#i�W\<J��6��D���H��*�@�f}2�U���)7ҽf(����~��+���
�r��q;y�l�1��y�D.�`4iI*Y�d�:����O�Rw�M@"�-����B��@�^	
lZn�\;v�յ�>��ߌ�I�:-�F|,�Ø�SIV<L�t����bdp�`��8B!��� �")��=�I��ZR�)���Ϳ��Q_'VOYX�e�R̹��hL�`��F���D���v�}R��Q8(ȃBCgg{!jɰ��U�H��?
�y0Z�%�5EET��q
�>z(�y�kǵ�=����Y���� -+gU<v��c�����Jq1�������g����7����6�,O�����yT�1����K'����D_$�P��%2u� #	��� ��2� 2;8�x����ju86�}����ҩ3����? 5�buf_��+�հ�T<��R(m�>$���@h���(?*���VH��0��%�-�{�t��Ǩ���SG,�mHr�V6H[��Үv�ȩ%چC��:���$ڄF��T��?��$���t3	�ĔYC���$�Աp��M��9[���Z��p"Sqњy�R�J'6p8��{{�8���7?+�N������?d��*��D�4�_��Hg!�����j���uL�9VT�C�PX4S� ����֎���ٳ���+�S�S	p�R�P/R��P�3Top�GA�Yڨy/;a�%��F���g�FA� \��Ĭq1�(ڀ�l��7�0����Oʋ/�����{����:�����eO/\������C�- :�.�ԐI����L��E��o��	C�̘�+W̬�%8�"0�C��d~uz(� P���E�B .�����o�@I`u�
6�?󌜽zI�.�FS4���hn(�^j�)v�#A�$F������ f�YDB����3l�p��e����p6�
'��ӡ�PJ�v�45��4J*.���z���"S��a������(-�;��.N��R�b�O܋)78�D�a�/��:�О�Ю6�֖s
�g��B��|ÕG�l��\5�Ie��  ��IDATu�=Xnv,�#�ƭ����\M�j��<B*R�o+�I��e;�̕�<�2����̼a.�C��@��Z�F%_x�)������9��IEY�y����c�cm#��0�^�,!(��ޏ̫8=;����-�9�-�֩w����P���Q_�K��L��ч&�X�7H��a)(򔲀,6��tYQ�=V���ˌ��p���`�r	39�[�CZ�"S��@K���~���˗/����^|�k_��ţ��7������=ɳ��I����������?��t�d����0P#j�e�Ǚ��i13&D*&���D�Nd�<oW�DQ<(�uk�)-A���a��v�q���������P8Ǿ&�:��,F�!v�X�-N-s@��	2���&���"�����2���JI��^[�M;�舚�U�S����ᆗ���^E�mNS�3v~�Q�Q����"e�p��������F�����t���p��g��3&�]LY��.��䁡���&t��5%*h�	�>K��BaMc8G O��b�`�����_���lYqc�� �<��w�}�|�X���p��7u�,�Yr�{�T_�������3;f����*؉������T2�M�lW%Y]~;��r��5"e� �u�%��� �����_�QU�d�ǦZ�u���F���vl1�_Z�'�����`/IK��X�� E4�����U�[YK#C�A��|���!Xj>�QP���@�V>���k���'��y�������e	A�5%��D@x�����P�pG���f`�6��7[�ǉ]9��HJ�Ϣ�W���B'���zVQ�7���p�
�2� Lf��J2�D��"7;�s�
3�WT�ۃ��f�l����-���NY�psh@��NY_g�k��ji�O�HF��8�9'�j""�P�3��O}Z~���ݷ��^Eq8&�6#�p��\�r&��:9�� �p�q�3��Yr�X�9�p\����[�IC�
ll���B�S�,T.Hy̠~�TЀZ�ZS����>�=�0�JgY'\�a���	�^pGG�[^�4�<��˨��c����x��uS5Do�F���Y����;��jwIG��

�Pu�!��*��Ȝ`�676��~m������-���伖`^/U�@�\
�&u
��Ҧ>�C��S7�E� ����kq3�[(�ۓ�|��7����5u8¡7��f@��3{A%Cfi��pNBI,{S�,�g]��=�w"�z���}�9ܕ��$[ױ?�1#5��`:f��;{۲st���Z���@�u�6s1��1B�wЙ'W�e��Y�:
VK�B��gIRϦU�T Q/�E���@K�1�"S��5og�W���ߒDz";�]j�<2Z\GA�r�����ݽC
�$�`�3��@���Cu�k
�߻�����㠶�����kZB�lU�cf6���E(��#��ʦ���F�e�s�s��.5�rQ�޳�=K�5z����������k��[�,��L]}�����<G�(�	�BU����tV{R�6�80�K;UXTY�fb�a���5��4�����tm���u��K�G6CRu��O���g�"x9MJ�(��f�~@0<]�HDf� dF�B�����=:I�qׯ_�?��?a��/}�K�L��CJ��hjkaӫF?ͩ��#2o���a傠�g��� J��K��Ź�NC!�MHS�ZU ��~�	�B�cpl����?������w���P�F���3aa���}h7���(.�,$�`M0�>�}g�&��l�.��dft&���bIi�ʖ�3��f֦�}������+��3f�|-�����ȋ��Ojue��yu��p8�z�l�^X+#�% ����d�=J��s��V���>$�T���{��9�Y+ AKj}!Yþ�|
�O�V=V�b�=���&���������Cv�
Ho6�`g1�LeYaq�n�/���:I�G14h�����k�(96N���o绽LL�G�p�̅�
�&ΖI<�m�G懟wDl�gσ .G�x-��*���x�w�oSڲ��?��Cc?�#���m8��0-K�8ҡ��T.���V�~����>��/��䑺�YZ�1��:�@�ÎR�X�����>�������wž�~:��)�&, .�(��l�A��uNfLvdbu���@'���i�
�qF�)K-NV`V-�,�6̣�>�RW#͂���|ƞH�m�����A�Q�ض!����u9ͭ1nQ7't�1�r�12�q�m��L�NF��*�+��5������~�EH[�� ƛHd�/T�bs�L�F��C�7u^�����0��2E����" �Ù;p�;d��ww(��~X��{5�w����sOD��]�d�3���O�K/�##��A�"�$P�Ϡ��-u& Lq��E:��nߖ:�f0B
�p?MD�g�����Ȓ�}M��7B��$P��(��3Pg��ֆLĵ�:�+�d��?dEfV�f���ԡ�y}uM���/���B6�mʅ��("tM����.��h�"������SrjeMƨiT@ӇDZ������N�ǯ`̶f�kMՉS�;Ng$���J��I<
� R���7��@l��OD_�\�Ȑ�ݓ�|���wfSF&�":�+
k
�����x��9��z�zR��֡�}S�-�9�cCl| оB�p�+�T__QQA�Z����bh5�2���tW���Ⱦ���bLX<�%c�"�i`��@��'�E�P����	��(T3t�]��w0��]<
���U�{�מ5���p6pWϬJSg}��@ m'�����߿��d ��WP�B}�E�W��15��#O��
.��}��Ty �7�j�&�xHI!tp��}DFv�s�����ϼ��\�)Spρ&�?�8zf�Z��	P2S�;��̱� s=���"Hc]�-�&�F���0�cK�@��_� ���L�gӚ�$��X�����`G�;�c�?|#�s�ʣ�Va4���Y���}]���b� 2�x��06�;`��_��ڲs�����{|��A��j(��IjLX����hz���:�G����N�x����U>����3�� ���^l�Ɍ`0CoT��}?<���{��|�o�V��o�`�DJl�bͨ#��5�g���:�F��ZX_P���� ��$�텠4�&��|̲R�&c H\���d�?x��U���\�cdD�;��xК������d1����ġ�� �2����#�!1��<��pU��@�P��=?�:~�����W�Q��%i܈���I,țG�����޻z)I����z��x-PԎ{6hz��B){�RTi�n��!� �/ep�ma��HN����ړY�������K#����1�V�*�o}�MH�@?S�)�f��>$"iD��LB	�����b(�t��u�y�IRy�e�Px|��F�:.)��>%��GȒX�Ibj����G����:&?����<[k�ֶw���=��>c��et44�Q���ld&S}�u�qVV�x����>�����+��¯ H�����y�i�9�4B�#�'V�|�K�G�#\}�i2a:��5�A+�!�$��l��	�* ��Փ70�����k���@��"�'��8B��tf��`�f���:�)J�H'mI�%�|@�pr!�P3���d(Q'H�(����#����r�WaQ�+с����P�r��� �m6+��|h
"�*��	'�N넁Z��֐�)�v�z�p����o�w�����An��P~�_�����׿�M:���v��u�r�*b?���>�q�;T�Ё���Q`y�N �W��ݖ�^ǭ�M����f0U'�Y#cȐ��$[kH�ӥ4=���N���H����UP0�x�poܽK���K�)([�,��f����b):��H�)bb��� ����r��y���]Sg�O�ܿ��/rY��6V��<_�tQ~������/����tp���{r��y�Qp����ꨍ�e{����Gt&�e��Z�q���T!P8��Hr��ýRR�b&9�J
��r�����A��i��
bԲ�j����nO��4��6�|�
Gz�Ad���d$#4����� ¤]B�S?�z�<(�C]xnKXj����kdj`�i��� �	�x�|M�ز����X�0�隳&�Q	�9A��@A	)�������3g��;`�t���]n��t��LX˗�v@��CY�t����6���<�9cwmM�B]VA�ԹV�QcWg��]�s Sh�������a_�$h�����d��@).����/�$ց� ()�sQ�8s
F�8�R[�qN�6�7�x�ph�u��h�� �5\����c����zvP}�`PkJvh�$&�1H,�T�\��
�#O,�����h5�u}k[:Y[fǨ��.M�Hv�Ά��6��t�>ǂ���mTu�D���.��rWm��儐"���F��?6E�G�~�iY__gd��/���b�V��,μ_�ՃǨ�|3��\Qr����|�~�Gά����!q�t�D�L��� �v)5��E�3��d��ߺ�:�6"6�@>����՗�,��Gd2�X�ǹ1l�h�g���O(ލ��g��Q�	vt2�1�٪�dX7��?�~	UR��ADcz:z�����������rL�8�!�����0�1�TȂs֩�a�V��8}d�T�����H�3I,��Qk`��.��@�Qnr���Gr����뿇���s�[�X�8�c�/��ƌV��Ic ���Z�\A�G���~�a)��Q�M�+x�Qj�&~,qh���Ss� ;��rb\�"	s���"�/Q�%OloKbH�s�˪�s%�N��(�!˨܃�l�i��17�������������� nSp��H�J��É�[y�8y�w�u��u�B�#����d3�p�Z�t�\iꟉAKSA�g�kK:<2��P+KY�_\jTZ/ĬX+������	��I��y�'�MeI�������+�V��5�l�׸��K�b0h/E6����d�� r��v�43��X�|�I��*�L`���i��G=6�H�o`?�/3��Roi����E�(�'|�Hq~X�u��ݍ3i�Q��*�j-�gV��z'�qæ��-��voҗ[�o�4���s����99�^���_�����y������ȵ3����S��懤���:�i��܄Ͳ>�8��L-B!i���.^?h���`�&$��1et�{�:��#.���x�m��y�x_Rd6�Y�t�����V{fuN&�Ǔ����H�O���-������Y7�?��_0���`E��N[�����^�6�HxQ޸�!+k+
u�V#8��4��Tc ���ѹ���WW��+wTw2���X��F4�G�����n4��0X/=DeRuf��Zb(Ǉ��Ľ|��l��U31�q�ã�:sGƙ�����.���������Щevk2���P���B#2�#_��W���ޓ��
4�X���Oxo�Y��g��|X��g/I�ٵ��.��:��,f�Ec۞e�8�!d���̍�Ɉ��o��iv�k���&R2�H����񝹘
���N����ɋמ��̊�Md&��-���ߗ�2��*�|�ڳ���Yf	���b9�����=��)�����?��#9��@�p��=��zYzEo
@��� �7���(� ��p�,�Q��5ēRs�`�,z@��!C !�^~�*���g�,{���T��u��S�5��ڇӬ����iy��Tĥ�)j��͌d�fi�N4 ������?��Sr����	 Alj �yfY^�T�p>�x���>h�Ȫ�!�me���<ÎJ��P��S�T?4�w��R�M�0�����3RB�
�ZoY�Y��F��u�]�c���#���ؒ��O�A���\j�>*���AMl�P�_c���'l�QĜV�����$9����|cHl�4�{�����T�D�sZ�3f10T�z�S�Y'k*�8�6Q��=��Ŷ���V��op������u�����矗W_}U^y���u�;N������0s�+�kR�!T���I�?oN��rϓ8��
��ƖeT֩�͆�렪���P~���֎����o|K���W˭�j�m�����v^�^�r=������+�v3��=B�g�[���)u"�7�=������Z:F��E�H¼�s�#<@{�����7,�=za*�����
#��lz�bp؅ 3�/���'4�$
I��
�����C�?��Be�����ǅǦ�������@/7pR
E�A�;�I�A�V�䬬`*��?c�Dt�O����<��5*�%�e=s�ZY�F�|���<��� ��$u�lǴu�R���u�+�y��?����wP�פ�
�1��m:�v����z	`�=��)���	��X�����y�3�⒒Ia��wJz���X��y����^(���nz�I�D�,�k�b�>�l���=�����3=PY�
-wN�^�����rA}��7o[�3 �@�4��@�Y�����Y�Ӓvh��,��hB��̙s�Vf�l>Z �l~�O�B�f�egW�����$�W�K}��a)�;�Ѽ��k��a1�S��$�2;^0��
���h���)[��u�9]���<�i�����&���)jPH6f��CuDϥ�r���H{���~��,���[�0uALx]Lg�V���'�;[�++�SO?/ߚ(��RgC�F�z1)b_-\d濓�@�l�E��Ic� �R�HL؃�}9X9���#�VoA��.��}�y�CY҉����zs jA#cFDc�ې���> `d�&�!iIA��%����P���c�����ۥH͚NJ4`�i%�`������w��ܓC��~�X�#$��7�e�!}���em:��cu�_��])�un�����#Ɂ���*e*��R�55<ֺ�ǽ�yW��mȠ�=�Z$��^o��+
��tq�>�~c�쩣<�{��u)%~��9w�������˖����, kVs�ɂ�dL��}O��\�7%��>?�(ni�3�̜��ǆ��-��6��h�sǠf_϶��I���S��e�)7l���e�_��|�p_�;2:},ݳm9���x�����R���7󙧞����Z�P��ξ�u�����d1$5,�"]]�(�=qM�N� ��3�j[�NZ������D��w�$^��c��qz���
3��LGQZ� =)�f[Fz�P|��<,�9Q�f*��|D�eXk��Ҳ,�>y�:�����Z�ƼE�� R���C�M��9�PlS
λ7ь��ͽg�`�Tc�$���1���&',��TA�b?�yS������++�;{���~_�����ޓ�o�M;�ӹ��)P���͒9�H|�܇���)3�����D��>Z���F�Q��q�$j��}���6����RI
�,�O�֘}��r�H#��}�YA�������� �7nps��z<���?�	���>&?�я���[r��y�XF_�Bf�� 1�(
�lJ�P�K�_{t�.k]�չT ����2[Z�Y��t$#8z]}ݸ��}y��w��PA�[zF5i�:���lX�@LX�����&P�k��,weme�5�ә/b�ϗ�����dI.r' {���)�h�f�d����gĬ6+�Ɵ(y�r(�y�|^��4����Џ}�1L����!d&��j�5)7�P�ĥ"�O~;VRN�DbM���K#.h*q/=�	%ψXH�����7UG��-]^ң`ՙ��e!�k�nM�-x����W��u��/��mL�>f7#N��c(����I�f@!��yp�늌3b�@�)l=��D�&}ᔿ���y� �Y�Q�p�w�<KQ���L���C�'�D�D]_����D���ٕ6:�J��'��_�W�v��}��SbS�2���ј�I,�C�\2a�z� k�u^C䰜����=�-���G��R��̸�����6ec�_9#�[��ZZ+E^�3����������c �{$g�3�+#���]�*}@�j<�E"{�Yk�Ĝ��z/Y�'�����}diy��=0��5��)����՚���	�X��kXJ����.�CM_A�n�-	�/���z�W�'�wn�+��n*��n}*�fV��ҍ����]u�jr�ޕO]V:����𶼷qGf
Vv�3��ߓq1e׶�͞\��3��I!���ւ��Ĥ���7!RS�@�h[��>V&@��3mR�ZXG!6vu&����ò4�Q�q� �p2��ё�L�+��D�Q?�D7�YTgSd'�o���a��Wܐ�������s���\lͥcӖI�w�i^iw��@�uOݕʹ�:�Y=(��]u:eo�����d�lk��S��3��Q6j�(�Y�2o����TP�PuP��Ã]9��� �I�ׅm����( ���!5m��YZ��8$H�)#ڈD#�2�cM� ��q��i��J��������C!��ŋ:�C��A�C4������lZ��@s��/6
�(�E0c��`�*�<�<95a��4��� �Lc������q�k�F�z��Z��⿑�fW^��?ʻ��g�ly�'���ȅK���}B��7��Pn�o���ɻwnK[�����ۻ�)�:��/|V��O�P�RwmUƃ-#p�k�.[NL����m�k�Q�o��OA 7�`m���A#�����9��k�:��b����9�b�NH �q�Δ;>IV��@&l0��ޒd��9&PzM�����qCf
��t����;P���G�^�j#�X�6�X�H��
����0�:�|�؁]�,�Z	�3�sv�賅���'FM���+����`J";���@7�gR��a AO�����ŵkO��W���uy镗e���m&&3�6��b�%��� T�j�h�����,�� �@訽���t���zC2���&�� ����1;��Ny/���A�!	a��S�v˜�c��	A!2�x�Yʤ�.-��P#F�
H�b�_�zU^��g���SH������a���X�0WA��}t.����:��ᴹ��>e��	���(nH1+h�E��{��d@Ё ���i﨟~����ǯ����]iwz��)��]��ru-�qb��0y���R�!]��]�̚l��%���c` ��dl9 r ��h�ɣS�Yu�o��������+4c��|��h��|��j��5^Xh�4�A��e:C�W�xd$t��%5�N�S��!θ&p.��7�9:n��$���.�ż��5��S-�kL���O�i�-���/|��̈���5NcﵘDJix�U��e
b&<�����z��Ze��Ra�_�c�=�JFs�{�P��۠ ."���ݖ��,��r	��,��'�Nq�x�Σ��*����D	TL:P�;&��@܃�_��s}��Z����˿����9�� S�?)�=��a�.��<��!f'M���@���}\��a��jsz��=�=g��阼x�������G<�@fa\Z�JG�]�&�����ߐg�?�ZF����*�>@=e���0��?Լ'��]j�I�z���t�n�Ϫe�nk�1F8�i�P���.6�M������~��
;ּ�,�"�/Ǭv��b��m'�O�:�1ڕ�����0����� 8ȺY�Q}��%w|_N���-��\9Q޼[^ٹ#���*Xj����6�7d��/����Ʋ|�ɧd�Ӓ������dخɾ�=�Vڤ�!��(R$��S�&�Y��K�����Z���H��tr��Ķ0YR���#��Ý7:J�>P5h�:���zr�Ie#��e����L��	��z��'�q[�ձ����V��V�q�� ŭ�0#BКY-Xp����T�<��N�{�3۸i=fc�%�����>�s�~~�B�b{��b$��`����aQ�	�:�х���t��N�#���^���3�:�Ym&�d$�fΦ���|����?<��p$7���>�'�١��ڲ����3�f�p~P���*@��� *.���Ƨc�N�T�����ߒ�+�@���-�}�/���#���wd��{�Ucc������L���ܣ2��hA s���,�#W�'�͡�G����8�i2e܄"�(��7�5\j,���5 ���o��`}(ӎ��Ҹ����<'��e��-zE��UP�w������C�u��i�է���~��IIy��7����J��X_V��˦���~W�_�"���ZWЉL�P���9�F�U�*(��HBA�d�=�"����@��M{-ӎL%�Yt�11SR3�Գ��>g��5AMb��'�vCV�=�ۻ'7�|�nHz3bwtn}�����ʚ<w��,-��l��P�U?s���7�	C =�@�Tf@�T8=ҹ�����$$l�aF�j�赆�
�=���?��Y/�Bzi�@E��0����@6w�>_[[Z���}:�(J��Z&
���k�.��Q_����q��Q������P6�)k���@)���j��2�;X=4�cP!r��Y�7)Uu���E_��(�YR
��Y����d��=��P��ں����3D�Bl� ���!������۸'�;�
/əӧI7�W��_�����<�	+�>{D������8�լg?���X/����YB�]��Y�;�Gl���~���懷卷o�ݍ-ٺ��?���jw�,Z�v1*��	V��!����<X�4�>ѿcODp���}L.辋���;7ߓ���b�&��&$qMqˆ��&������0�Ml�D��4�X�����)"�|�^!k�,�Ϩ"�I��S�i!F:��l�˓@�W��F�g=Z^���*`Z��� ��ד�Y���b�9�|��PL� ���ItҒ|�/�z	�����Oa~9t[�{���Y����-/߷��k+�/���r��ދ�����C�
�4��q F3������� Ob��$fe����:^1�.��U�6s�3)�7b��葕��C�K����GNL}N?�6�r�"�#�������P��r�	��|'�/�q*��y��#�
�G���b�2�Js�L�N^���=eC����9)(�p~��?�%��l-!(?�F����]�o���ë��ܐ��ϓ��yK�c��?�3���J:����K�#̦.X�e;I`�TY��m�ȽN_dG�)�)�^�rY��;�$��}{s1�KlU��0������}n��F�#Of�Y0O>�@t�v��g�(�tisE��&��i��c<�Yl�h����@[�7�'<^ݥ����cu�!Ģȳ�-F�cY6�E٠��v�u��AF?���n�(��O��-�kP�L��#�zhJ�zVz�tz=:��28� m���{?�o����d׺Kr���cN$��8��PF
�.�y�`Д��׍mG�!�qZ0�'e�U�_h����X��v��<:��Ft�ysة@XO�H?ԣjVO�Z���k���"�!�q��rd%�Y�g��[��po�����F_fzl��:H��ؠ|+%�C��;����O���P}V�Ǻ�d8����:Ǡ*9><RC^�W�>�{�z}#��������-Y�ݐ��}R$��C�kn������DS���h��RS����8��[k��1�beέ]ە��-P2�`�^lޝؼ^Rp������e�S��F- �`�n_F�Lh�Ѫ3*Jt�SC�Q�Ŋ������ʴ����zU���o��G
<Nueo2�����,o�o����/�s��O<#�Ͷ�c���?F_ɑ���3��Z���'���:�Č3�"@�@���ll��h�0Q1u�=5>�m@=�~BL�:�S)أ᱇�xM���/ЀQc�PP���eX/�nA��<x��M)^����r�ѱl�xʚUp�A���$���#8T`��26y�'6����ѩP�cM`I�kQ]f�kVW�s&^�Kө��E$�L�lS� �r[�nm]~��ϰgӹw�.Ub{KK��Ԧ:NO=q]޾�>E�؇�170��7@4�`?@x�LGA�]K�����΁FV���%���m�U��j��{��H��x����s�E���3�����xxX���4J���-fkqon߾��2���hxK���Ȑonm�f�!�_���@�u��u�����(��.%Óy�_��Q����T�,�bQq�����2�Y;de�bJ
����[r��rosSA�ܼuW��Ԛ�Q��������X_�JE�/�nm��m����t}<v�<���r��i�:�PΰwtH|��	�Kq�P���kօX(I��~Y��>R���^����F���k! ���BbwZ���)�����sp�{?J�iZ�d����q�s�J*n����Ct܃��_�R*|�࢈g���yV����g�Ԯ5�����?d#��Q�)�i����VQzL��"�lTя|�]�B�'f�9�W�N �}v)�� a0��/�B���1��I6+�e�g�b/&]8K�#(؅$s�ST���s�y�b�*�x�vU�4���*���dRB��v2C���pb���k���j�L��G��ߘ�r���5�6n c�V6?U�q�:��!������LR�:a�o��}�ǒ��\���=�j#�ЁӬ[f��c�Z�����9����o++���ʡ�b�Ú͚��Y�����k*~@���н�=9��y��jSz�d�!�l7m^�@�0A�1��h6L��i4j������Ss�}��lO����z�P�'��M9�K�'N������ڙ�S[b�I����&�5��cƢ0SPYٯD� �q����XM)�N`!�s���ƈ�u���4���8���C7��Y�J�X�-(!�jlp�����w�0zp̂X�@o>����#�~1�>��2 $QPh��/d���x�_S��z�ŭ����T-֒䱅F¬�0��$��GvO!Q*,�O=k�T�"2C������qD�uP��C9F���X&]��b,ۈ�gS�Z��W��ֱ����;�Sa�ڑ�A�������c��ʭ�c��et�Dǵ������X#J����w��ү�8��\��{r����h��d��:��bs(�)�1�biw멧��Y��Th���O椎y�@R���UJ�����H~�^v�TRe�r/�K]5Z��0��,I��(/&���g]����Җ�=���ֳ����v�m��7~(o�ޓ�^&�}?�xRQ�6���#�n��wn�e���NJ��F�֐�U���:٧�I�2�� �dd�P��C�������U�n/�g?��\�Jhf��\8ɷ��my��dz�sf�e�'F�B�#Z��q�u�.+x>�D'�1RDtl߹G��l�"T;�۲}��7 �a��)ԩ�9BeqM�-[m����y����Ff��G}����A�S��V��,��`�l9�+@O����y��4q�B���}O�\~P�A���p��oo�����O��e���5���"F��	w�h��:^%.!�c�yJP��������s�KH�d��CɃ~@�{�0Zt�_�/F��>�1J-F����`!�R���3�P�ԸB�c�y~S�\�̶��D�2d���pR���q�����b|���mҥ�C�|�X��ͣ��ut@�#�|y{����@���w���ܓ���ͽ���4�o�C�{�=�1�b�$�49 Lĳ�Bej<qoѫ3Q@�zt|8���k�^_���ԛ�e� �R�
�3ݩE�gl�5d��E��赑�	E,N֌F��<j�����G�kF
'ki2ˈ&�5��T�0���gN+3Ϯ%T2v��:Cq����p�����
�e�˽t�����8.�}-�e��4��,� �� �M�`B(1Se`г3Y�U�hr�Ј>�=�PP����{��R\�1�U�����ѿ���~ϒX�N�$?9u 8�S^3�X����[��Y���@Qa��8&�(M�~���9:�`�TU�_Rڕ�D�bѼ��ډs���t��c�NJ�]�Zp<9��,�Q���>41Zy�Q�х:�Yx�s��`c��1-��#}�C!&֭+\ZV��5ʨ��u����x��Z�� ��K��L6n��~������k\�v��[�n��	��$���:Mo&�k�먝��&�=��t�R�un,yKZE��c��x�9ؑ-�'`��^�"K��J�9W� ��4̤��^����$)�R�s|�Ic��3�0+� !C���J���6Y��x�6^�c�M���$�"�ݮC�J:�(�����(=�e"�U䤉�ɃtG�����,]Je��:)$�Y�O7�8�Z�ٌ���
�mPR��TU���n�E���f�)�Cu@�ѫ����L:���:��42�J��d2T�<�&ިw(���,��J ��I<0h^s�����Լ�E�`�gh�=5�V`]�5��A�m��ӆ�/�b���B�+��>��C� F�Aeey��-�Ł�%�`��	ivȦ���5��Ă��cu��N��?��҅�{��`6�<��A[`���R�o,�9�0�zm�A^`c6TC�*�P��͠Aj�c~�8�{#k�#��S�Da� J�CAϷ�8��4
��#h��?�&�n���P0e>�SRVY�9�ɶ�~����: �X��~��h�RH��q@�h��7��䙜g
?.��ԯ�ë/���zEޛH��@�f=�8����m�t����Mߝ��F�=\�T3����B	(�g�xZ��������.���T zp|�NsKV�te�}[6�ߧ�N�J�'�����\:}��y�(�"z�j��&?|��U�3`�@���,z�lu^�Z��{gAPP��4������:�(B?Թ�6Ө�;��Y�z^6�ݓ�ш�%��̇�~��O��)`8��T�U���έͽ���^��~�oIcmtSy��c��3����"�ݟ�0�`���l�}���{���D�VD7� {�wڬ�EQ/l �D�@Ίޫ�g������]M�}�,��!$nޅ��ǖ�Ĝ��bo!P6Q��{�S��ڼ���N82Ѷ{L��V|�D��Cߩ�̢TT��`6$s��؏6f���;����b�-` ُؼ���-�v����5n�K�7W�m�ڮX�t֌����<�ކgEb���ҙJ�>I]x��Sat4 vP-':G��C�@�@�֭�����}RꏎGƠA��X�7���[�A1��d�5#ά�jTN��\�pQή�f����P>��߿yWu��u��^�=�"#F��j�I^�:-i���L(��=J})$>�)~h-������R�7*��$f��d���ы"�MU�2�B�I;�e2���N�gIͭ�5� G}��C�D��U{*Sw�(����Pfh��1�u�	��~Q��Eˋ;1��h�1�g��3��~~�͵RM��U��SG?'z�|����p>Z�_��S��c5�qP�wq�����;,��|�#�O���F�_^I	�<x}���恳ʷX������T3�������ROi'n�Of��j^H�9H���iei%����ʼ��)��5*!�,)`�^��>������&�DR&�u�!� �hb�X��fe�5��]�ҦU3���J�_'cH��3��P����X�}�'�7^�������?�M�w�4�]*����ti�{����@c�Y��t �n�m'��SW�=�C��^�J�C��c �xt [���?l�^W�<vY���~��/���x��քi��}��MRT3�cnqi2g3ȼ�=�96��uyȾA���,K�ʠx����i��"$�{�ߠQ�pl"/�ԣ����ڪ�4��L�PC��d�Do8j�Z����򨣅f����D7v6N����!��Q���Ľ�o
�b����aŜ,�ESo��P=��If�'��y��@D��NJ3�sK�|8sA���A]�M$�HiM|H[:. 5pffN{CЂ��@�:�ΰwH5�Vl�`��q����{9�rZ�iSHCAL��R	������e���Wmfￗ��YR�z�A����Td�4Jf�Qx+�9��hY���2���@ 5B �z�Xd�F� <�0M	�3M"ESǨ�[)b�n�{O�:�j�~���X�f�`f�ZK7�q���(*���c$�1ހ{o
d�5��E�������F"��%k%���$=��QS��ʻ=�wg��|����kO�Ԯ����oˍفl��X��ͱF4uml��D-j0�,�i��kt�G:A.��y���˽�҇���`2�B $(��B"p�/��<����ߐo}��r�w�w"�p*�����}NV��d��Ώ_��*&�d}Lmg��&����$Wj޸��h�fmfڤ��:ԉ�i�|��LyA���u�{R#Z5���?��ߗ�^vv���g0jJ�SLE�E���!��ڗ~��_}���ӿ�)�ڷ�!��P�wt��,��ƙٙ��	���0'�B0)Һ�8~f}!���m#�{��ի\#h��ݰ�CpBf%�U;�DbM�hʜ1�U��xT#8#��I=3��&X�)�x�5>ĳ����G�2^���(ڄs)��� �x�,au�a?@�@��E���NJi�kG�&BU�7僛7�����(���1���"S�Z�f������Gė�K{�=�*��$P�N��Ͳ�GP�,�@�
*�w	 wv�u�?`m�+��S�3�q!��1�lB��<���q�P���}�HI��$3R[��ۭ�4u����>W��HSBOλۛr��]��ߓA1�hY),�3�]�>_$�C{=0��}QetA�/��s��L�p,��-,�x�4/� 0� .���ʓ�kt�1�D[T�l��}2?�;�R�gt0I)�R�n~6*p&��S>E��P�^�Qc�.f���h_����r����?����u��)����:�J��r7s*�H��B>�*�n7���s4��
(�-���}D�=,���V��k���W�٭*���2�!�_8���|XӅو}�m4�^� 8"9�P��e�K$f��W�{���h�#ت�9Vz��`�+u&��Es΍	�"�Q)�τY��,C֪0%̸+�L�D?�"k�1�@Y�w8{�Ը�u�t\��E�� K��&����1IYӟ�>`φ�a��eIE�y/ʴ���B,B���I ���S�7k��l��ĕ+�d��*�k�������~���Ů��a!��  ���>j���P1�'���ی����̫��/!����{�rw���:�?'�+��;���Fuz}p}���[m����Z�%�&o�.�#�<�E��!&��U�{2�A7�k�g`t �=�fJ�s^��Y'��{m:�i`��n���6�x��d�j������J`����Sr�L-� �GN�I�Z�rF����;�`� �I�Z7��ð�=���NP-[�x�CqS��Z���6�3��)BӢ�6��$�o �(@��Xf�, ;VPp&&���	���  ��{�Y*��g;��>:T���)J0#0H9^x���z֖&2��𨑊�>h53Z{D�WtRfG\��]+�H	('7+ �
f��i�iI�!N���ap����|���1Z����e���x��^pp����g
㋺�cu��S�/`�9ܷV�E��oCfP��rQ�^j�Q3��^G�β�U�;�w�2�c����{�x`~�u>"P �j!!����b��)�}��݉�=���a(��\��|��u��O�:�u�����ҍ���پ��R9d�:*S��	��#l�R㒰q��.��@j���}z����7��;�wX���;5L�2.Ǉ}Y�����u�GѤ?��W�o��sh�k_�2�/y��59s����yc��ʈ��"}�8��F�X]�;\���l���زꎲЊ��7 �1�K]�j,�yG��G��z�{�ē�9׾��_��}�
�i�Sw�0��
 �M�����o���U���7l2��bn 3���jf��`��_%q�d���D���ږ���n�u;m���:>;�F+i6e���v��0ߞq�\̅��~���L���7*��d-]�j�nj�)��DƘ�� F�'oI]u:�I=[DQ"�gp�p0WeGfI\;1И�� c� 	��)�S���*6Y�D/��Υ���`��@ �
Ѫ�$��1[����n������6���������
|"�
�ͱ>ֿL�F��=W)P�� A�X�ı�f!É���������Ւ��^)cczk��NF0 ��3��u`w����VSz�t ���v�V���=V�`soO>غ'[
H��cDp �%q���z��1�TC���߰w�u�/�cQ���Nf��y�c��<�\��LypoN"�?lD�p2�wތ==Ǥtƃ���k��j���Bz/|��im������>�;�س̕�.d�l�s	��caE�~ܢ(�I-ȍ�k6��$����\�6�)�&�u��g��P80Mh�sLGh�P����_��&�����0;e�}B�}� `�k�D��+r��&|R2��q�-��Z�}�9�2��oxM�f��T�6��NN|=�(0�gX2f���L)m#���ʼ�%���\8ɃI�L�T?�"w>�e�^EU:/~��?����pq3H=�F\�ߓ)�U޺0�5��h3J��k�-a�:�-$,�M4�7l4e2����$��x8�R��ke��?gT��%�����Ԁ~�і��Ψ�VW<�v���phK����59L�7�*;z�f�Y(o��v���0/I��<���p�u����u��Ξ�	|�Lܲ$"��t�Ě�J�0O������FГ��[#rO\aG<��#�Z�s�	bp}�r�~�޼���0������fM�3 �i��<�b��"V�aƟ��nZ-u�;z��n���D'f��1�{ jԙCۃ��v�PC�f��y,����5F,� #��ij�2 �g!c��-�y^?}Q�����i�j��c���z�ԩ�&�Q�N�`|,��PB}i)���t$=��o���t����i���O��ކU��40��R�gT��({�Q��d+ �χ��<d�����dFBl"�F�piYN��u<Msfq��.�V�� ���YI���Gӂ��=c���fa5���"�D����^R�<:`2�I�
�G���?��� �S�����_�˹CK:jT���ȃ��!�^gS�Z�v�"���D�:_0���!�sK��L{��P���X��EL��Pw3+4x��X��̣��"S�4�൳�ҊE�*��U)m�}�K7�ȩZK�Q*=Ы� �Hu�kY�����+��Ͽ �������w,7�w�`Y���9��
փj��H]Y5��y�)���A!f��Qd�AF�/�H�6L�i����z^ӡ�֖dg{�E�_��K��;oɫo�.�&��e|<akP/��c�C$,$��f�ӭaS��V�p���
y4��itt[�$	M�����,��6��uH�,�y��}�`G� �gz�ts�JZ�Bd�%{�w���)Yj�X[�&�,�#D���e5��q�e�k�@�@��n|�nv�X� (�Bi�z�+����a�k���ѐ��S?Ϩ��k�	�rZ7.�x�Q^L
۰Hne{EL���D�REU��PF�~���5���(����ʜ�VM"���&�ף�x)��a�V ��m���l���B�#
�q�Џ�-�<#��tue�2�FB;�Lt��y��|<����2-(�UJM 5,�@�w⻑!-��}��N@k�~��<�^װ~���X���n����c�"�G�IR�Dk���w(��νM*�6�\�|��ڐ�����6��m�~a�hTY&S�)"�t��2˞�~Nu��3�������H�2kbˌs&q��#^���ZLsz硈��l�V�L&�\qN�M����ZX�*�S��C�e
�(�p�8fI�X3��^�$z�9�j�^���>�:7}ֈz���r�l��R���vM�	1s��
�%Ԍr���5���6��3wPC�\��25�?l.�������5cٳ��'pl��\Ž���eI�̨�lk�"L
�sF'���qM��"D
o�}6��[��ȓ���n�(J ��X�!���P��6R��'�JuQ�<3{%\����m����u���"��Þ�7��b6����"X�T���󱎒,�?��G��[��4FG{뉏o��ۮ�S�N���S<xȵ�S/���p?�'��֩qAL�Z0��שd���% Ҕ�� �(;�Ȟ���S�}��5EY���ʍ�7d��@�}�Yy��������ղr/�r�=x�t����Vj�ePˡ���	�gfOM�Q�)��9#��oZ��:�7���;���Ca2eɜo��&/�<
aT�N�Gd�+M}��̺�F��ZC�uBp|{xOڄ�;�d:�&�ꜧޓ
c�r��&d�X'���'�M�|�@{��z��,%���+����^�M�ԭw
DB({�?2��1�
�����}=�qm��"k�6c�w�7D���?ʇ���F�$a��Ա~��%y|�,���<��:���0�Y7Ss��5q֬94'�aˉ*��8�� uw��,�v����,��#F-�q�N�3Ǟv5L�AbFL�K��\	��q� �0$�H/3j:�&���D�Sg����kwޗ��Hu��yV��=�krm���]�,QУ@K�"���,�H\F���fPzjY�7�e|A�>rF�E+��t&����e���y4�W��%�fh$3��N�б8Ww~dit�q����0�f(Ì�`;�ɲ��l�ɪ�'��g�>&lݖ{�7�|�#���3r��&(�x����ѮΕ@ �,\��  `��GÝf^�i5&�@jo)�ه�ACUJ�?�=�jtBJ�S�����s|H����4�-�� ��S�|jb,K:w��tI����w������7ߔ{ L�I$�R��8��%�o�3F!g\S:Ms��Ȓ��1a�#s%YI�Z� [�ɇ#Yiu��y��H�߄6����jF
�:ܗ����q=�����R��@��T���W�lŌk3V�%���T� ���X�s�t�x���޶�����Ng�e��!����@�Yx�gA>�oz��X���.�S��i/3� ��j�cP���c����l���r����$����Y�Y$2u��<Mb����8E�Шhf1cX�1�O�<d�#����$0�����c��@�#2s rx>3�+8l�����U�i^��bMD
�9�FEe�;}�q��������c?2�,e���~�PA�H眵5���y���U�<-�g �c�Ԍ��kA$z�(5@Y@�e�����(Ȇ��|��|I���%Sԍc��9;�,C��q,8�l!���� p�u^?����kM��z[O!'��8��{L�6o�Ѫw=�O�<J��ܽi�%�q%�7��/������ H��HQjI����mƦ?���km6c6f�=�ʹ�Z#�&R-��� $v�ګrϷG�?��FDfU� )J��LdV�{�"n��׏����1������<Q���a
19���t8#<��e6�����p��j+�a���/Քٲ#Rg���W�ғ�
�`1��k>	Zp��Ϋ�[_T6b� �����kNk�%&�b�	]8$T�v�E(��u<������o�h��`?ա��۳� ��Sv �쵃�Ef�H���@�e`�@O�"%⃆R��KZb>k�v�@�7J롞�5N�_����#�d��Hk�YC�ǹ���^�\��ٓ���$F�.�g�fi�KYI��/��{S:j����1CZ��m��e���:3�X� �EQS�S?�,4��v;�/�<� 1��7mO���\��� >������SZR�ݸ���As�G���kꏀ-8�MZO��Y;6��Ss�g@���G�ɝOe�x��ʳ/� ��[�?�}+Ղ�]FW w���o�����������R$�#P�%����N���^*�����<C�������a£���ץ�IggQ�N^XI�:0z�-8CuX�t��݀~ƚ~����.�� ����6��f�`WF�3ڃI���Ɇ�)�w-f�ya����ꈣ�7 ���yIZ�AHY���%)qk���?���  �ț5b �* Y(��yz����@\P����87��Y�h��]N������e�ঋ-�⺳J��F�'���z�+r6I��P��U��8Ae�2�0�C�[T�WYvQF�c�y��P�A�-Jft���#r49�^\�b���h�jFgH �5����Y��`Po��x�F�����lgq,��\�ݹ!�z���1.��/�KϽ(�,�:@P���U�_ `!_B?� �e~�� #4CVS���k����j]��i)wu��A&�K��AW�'E�37[�u��g��'0(��i8�0 ���*�
�-g�dC ��_}]�ߒ=������.>&�_yZ�<wE��ޑ���<}�y�ғr��M���oɇ���-dJ���ˊ��K��@���7ƙ7#[с��1�9��3v�ќ>U����ϼ W�>M��Q\ɟ��{rc�ε�mA��>~Y���s���\���;�+����ܼuS��?�G����q޻�z�����(nkO���Ʈ�,0so��5��~�:AD���q^�t��!3��R�Ρ� ����󷣶hw6�����l�#�ЎG�o.���=�s�*h��B�����J ɭf=>KZ� �^� ���uy텗��&SY��(~�~�Ӊ�����O*�	>&�iXCcLn����^f�)�gu�A���dcs���3HѯOvf(�T�6�'\,)�`��i��&9~�L�8���=  ���hk싚[[Je��8�˨��(�q
��aj�ܙ�ro�a|n��V*j�ÕL�d�~.��ޖ�~��O+�9s欜9g=� QS�����k)�TC[�>W�+ݹ(��I���i5��s��|B�r�ϐ4��ՋCV+H&�T/7�����F���X�k��zq3K	�KeP�����dܗ�&�����-��mR6Sܕi	C�f+�=���xk[^z�e�^���S[^�"���(P�EO�v�O�H��6������G_Kj!�~��H�+�>k���*�c8=����X�?q��*��V��E�d]U@��X�Y�m���U+-�7u��v`[�����������x"ߚԀ[ ���}�#سˌz$&�*'U|�S����t������ n�'p_xz��szVY�o�K�D&���7�KI�^g^ƺ�I�a5�u� ��)��i���P5�Eb�whRo����A:�d5e ��Ú���ŀ"�����������ɐb�.>Fg��I �G`���_ɽ]ư�y�Yu��d^��QE߿��B����Y���	�f���,�d�G�`�;���x^��f�c�+.�Fn֥7��1'� ̵�32���!#�}lz�z�w?z�L��+/���\}�)���dt_��^a�fh.�`9Z�9�oi�vK%+u�*dG��9�'�;D���@𳠹�8�)PQ�C���Q}S���FE��^9��"][*h8VФ�([�W�桂�m=
�ru��]��^æ�{�7��P��\W�2������:�P�\��.'6��ƚ�us{��w�uB�I�	��PFP�T'�<ܕڜN���J� �u��r�#{1����ݹO��.��$ף����ɩ�7�����qX�n�m���!�S8�e��N���<@��Ֆ�5LXj�GGr퓏�\g$��u$��\��H��䤋сP@6B0ˣ������&r��uK����ǡ��졂��O��[�L�d8���u2R�QF����;&,c�V=��G��	M�"4�/{�:�w�),(�n`�� 
V棻
*��Y��!*%��4I�����衇1+u|'j����wWS9�Y3���AP�!�2�������psMw��H��D�Mpͨ#�K�@zf�A2֨��p� ,�	����;�΍������o��u�t�@�X�S/�p}]�ׅ��pm,cD|C�s| ��ܐ[�D��T^�3�)U�P#ӣ��1 W��1�����-��e^ʢ;c3�M]C�<��dkC��W�@w}�G*&2j#��0�ѿr��A�cye�����O��۲��������w��J�S0Z
w��b�f��<`�MͳIp�3񾃈�.���t� ��rn��z2B�xHKE��<)�o��s9P#�����MAل��k��A.��຦�c�E������"�
�){nj�e���ct��kd�UnM����?�C5��x�5y��S�^C�4����{�5dag�XV4�%ε��c�̺�9DRE.���c�-�]���)@���˾�l�=+/=����o��^ 7�:f,(��Z!����*lݚ2���̒: d���}��	�gɭ���P��(��J��h��͗��;	er�}����t
�G�Q�e��_x�[o�E1dYG�?C��)�,Nu�w.�FQ��3�E��nVF���ήOPc��A�l�P��ϫ���]69�)�hY���o��SD(�����0��h8�6.�	��:�G#b��+�9������Ѐ�:��J�����y�IJUuǜ���n���#�㺜t?ߑ�:�C��:b�{U���z@�Q�jy����Z�f��g
��B��un�� ���Xf%s�`���3c�^jb �K[z !zƦ�WMLR��Z 3V�7s��)�M7����&�ߟ��r*@���{r4�f<��	�Y��yD0�h�Z���ڔܓGL�G���OJе��`Ђ.�&ESm�Z�k1���i��l�)S�\�3s�,�n�S]_����Z�P<(dA�t�T&S%Th��)�ӓ��;��#��X�ېP)��G����xÕC�*a"�	�5�,UV'��]�7 ����k�(Ac��7Մ�q���91�� ���47^�:��K|��^�KK���2W<}�����i./]��r�?{�k�g�\,N_M�p�м�sO����;��ސN�#���$W��"k�+B��`0G�?���R����!4cb֤�!TgK�eE�W���M����U�D���JR�"{'��dD�4�<��M���l��s^��z�ww���K[�� *i���I)/�MmS�>�K ��\Z�f��27��M�������֨��C}��p�@G��o?�%��姸�z�������:�f*N@�E��#
�s��R�� ���� 1H��B�� 4�V��҇��Q�����ȇ7?���{rc�.3Ȅ�ȟm-0qpoz���L�K%��r��걦��H��ޔ�
8���;�W";�����b"U}���(wƖ�z����bb�� ��D�9��@��1��df��wn[͞��	P�����v��97t0~�꒢�&�?VM�R�bv`��~�{0.:�e�Ϯ�s�hW������H9�=�Z:TY4�?D!*�����F�����D�s_����Ȭo��8m�U� bH�̎���)�X����\���fp��Xۨx�� L4χ��
.��y���0&G:�]WG�]�����N��Ǟ���a���_r���|��e'׹�1��'�e��;rg�c��3!x2g�r�����V,RM?"7��|���`�Q��f@&��8�]�P�3�YM�͏?�k{�M	2����޷�1�`��q(���ߒ���We�@��?�C����rP-e�Q��a)j7#��o:S�::��&������<ȁ�JA ��YuH��E�!�g��5A6�s�&�;s^�{�y��:��o����M��x��w���̾~h���Y�����_g�g��T���S;�Kf�KR�
o\�@����mZ���}5\zndk�����0���Ϝq�.*9/Cy��U������{�����Cl�ZL@@�xW�ڋ/�\�O>���l�KBJ�庍��&�*�!��#C'���y����.�ɺ�~rX���WW\�0��jբC�r۸2wT2���q�͉M�?�~��D����[�:zB�o����X��Q0s̴���_)]�@�����ύ�UZ�HQWw+����7$QLѮ���⋒��㌟�n�z,:���?kk#�VP�����s��蜽:�S-kP�����)�w��玌���6m�k��ގ��J_�+����T~�מ�1I���4r���=��R$�iV-�1<q�����RƯ��`��l���r~�����U��2��Ee��L��m&��]
�%�}��N�u 6��_�V���,r~�f�ksP�g���-��g̤���f\R�d�~�a�Y�꒔kWP����BP�׀�蕁��{Wi쬿$z>�E�VgP�����q�^�����+�<�]��aa��pUy�6)؜�L�{R�L�������ח@l�Xc	$vP �?�m�L���BSm!?�u���l��4g�yZ���M������.J�
&Ne�mP�ϣ���R��@�,h_��k����4��,��J�=��
�d՞���� �Ɲr|�dj��
�6�@%t�c�<����(k1
�g���/�޸.�޾���L��o�s/<'O>���o�\�A<��(��0؞��9jk��V��f���+uf����rC�(�:F�ܣ$�UYq�=�~5���?�����b#k��5����p�sCԠMh������5��������ʳ�=Ǻ�>h6���0%�٥�:���Q]/�Zg���h�i�:{}�� )��a�(MX˲U�$�\Z�~xp�W��<�bQSF*b�j�9%pW3+dK��F�=}��l����2�ޗC}�(x����TP���,[�~k:At,��H5<��;�#*L��s��;�0P�C�\F��rir� �R �$�� +@d,\���TT�P(�]*�S���_�ey^�;2�}8���q���W �N�k������W}�S�.��W����X����a �����>�@��̺���STV�Vp�[]�*��(|�J�R��x��}� p�})�ꙋޒ�r�����8�gH��@�T6(X׌����( ���a)����c�ʕ��_���W���;Rlu��:�\,����;�����ّ��G���tcmM~�����
� �����:�=?����_��t_������?�+�?d��%���nO����+�M9���εS��~4��o3PU��*��0�I[��w�����T�g. @w�d����o�H�ۿ#��L�M�HǆJ������X�عk�tm�ܽ'O����o��������{�������f�D*a�u>�$��L�,��>�`.����fU&��M(�F�Χ&`�L&6A4��kx��'���Ov�H�u��0a�:�,;��(F�����@F�'%57*���E�?���hk�*����@A����V����{�H��Y�P�A%j����Y�%X��rYt�9���1ȅ���;x��A�{w0���Ǎ��:��؈UO��wBK>������9�@�}��9-(At8�l�6�Dߢ��-�e{m^��ӚO4�Xo��|Q�M��@��ҁ��"m�������M&
�e�k66Mk��I���~���^��0K'6�s�_�W9S#��?�л�g�5IC0Km��O>Ƒ̈����� ��B\}`�k��՟u/����e�6�\���/{BѶ��h�Ak�d�"x?���9a�"35�L����}8��6IZ�@'��Z�Cǩ���|�V��ipc	�D��CPʂ�5IE��xnK�/s���,�MZ�jOL���N�@�2�zΟ 6����L�%JY��dޢ�`�ޢ&�	a�rs�\q��ꙩL�_�-cUo�R���W�8�_j�Ӟ7� U�	�ch�Z0�g�HE�ׁ����aA9�M�+�}q��,���:��+�B�h���w��]c�!���p��fƎ�JY%�i �,n8QH���̑f�V��d����r�[O���9U�Gֆ����&0X����vY���G�0���`�e��+/|��,ӎ%�*]7A�^�g���ރ)�����-��k+*�P��X�l56��82�@�����=�mb,ۙ����D��w*CA�(�X���ShA�$�fϮ�?�2ԿߺK��ޥ_6Xȳ�?-W�FΞ?���iIp�i�u-��3�-�О�~4�2�C�'��3�f�q(���Ca2w��s�Z
�UȀ0+����`e�S)�ƚ$	�ڌ��7�����.�1�U�=D��vwv%�AB:Y�r2S_c�]jh���wF��"3�6�� �
��b��EȻ)r7�Ϣb�lD�&7Y���	B� ��� a"�.������qu�E�H�,�b;�d6����+���x��$_(���5��gU��#ig+��ØN'����@F�Wٱ	���@ Y�j�͘��T�D��FS\(hfo��z�%���gdXAar�,
2�h`>�1~��GR���r��)�rS������O�(#uDacT�� ��គ�,n|$���ZT0*��"9�N
�]̫�Q�IO����3*�3��.y.�4
!�BA�}������%�ϤsV��c��pKlʅ�X6����#'X���R>�o\~V>Zv�S����խ���ūri�%��bUo3���Ν�3
\���ߕ��XA�BnܾF�T�0��7�kp��#
(�9^�z���
 3�+�}��Ũ�]Fk��}�.���C$5���O3cs�^�/�t9����M�9 ��8�����'Gr��%��+6�����x�P��������kLs�?:d�Xz&՞ G������{�C|Ҋ�Q����2P����u�̜`��
D��u����{��;����;rK����*`B/Q�5��D���D��ާ�&%WP��������a+u�礮tL�x��^��\Z��S��@YQ�2��@�kE�p�P`�g��5�<l�)M�C>nye��7�6�ӟ�+ǇǼW�C�x#�@�_��o�v�K�/��[ U�<\i�����f�psw����L�^�RAf��Yk�,�����Tz�3���C�^��@�m���<zL��=o2��
�IsZ�J��f��Q{��Ԇ�f?�~���w��
��:!lSo��/��%����s��Z�^�ɑ�]YC�
���)�F�'���Ճ���L���������ؐ�ј�(��ʨKa$|f�O�Ɨ5ä���:�@���D+D�)~�:�9>�l��?�~���>-���)>|]�M��v�`HpN�	�VA�)χ۽�<xT�_O��+g�r���h8����ҟ*gF=z3�y��k�;���@��#f����@�k"\�F�/<ӥ��!�}U��ȫ4�38wMq�N��<v������`���5�1�c�F���8��M�)�k�56-|Om��X��|�4x6N�YWR/����LE|�7�T�B��lf�=KSRG�y�{<�{Ζ�w��t�A�4��.��Ԛˢ��P3�L��Y��[���W � +"+�~1����ZY��;Vf�g�F+�=�!' *V.fb� �}l�,s�^b��f���K[I�2��lM������C�@X��g�JeI�))�F�i�$p�й~���(��yG���f����$�����KO\�*�[?���ϛ�n�7�*(�}�e���f�GdQ@*iw�\�̋O3+x��cH����5�ѯ��~����	� mc��H�- 5�����Q��Ѐ�V������_��tr��e�e��ai�Vp�>�1�L<�O�e���}[l�e�t;mW����8z��k��߹�<
=~_-��u�"�c�&d�>Oj����c�����ڠq���8X�j����L�[��с�kz�Vta8V�Z[�@�ZQ1S@�qҰL�.�P���el";� �sտG��Dr2�<|��u�*�[k�	����ȇ�?�lsLy����
�O{Rv'rK'��b./?��<{�q9P��'�o+ ܥ��3/\}V�<����_��:7o���\?k)������bD�;%�%mh�d�k�5�*���{
��
.�}c�$�]��+������F(�h�0�a.s������}u�PǷ��-���������;rk����N�/������s��G�����\mH��	Tr��x�
���5f� $����3?Pp�%��ƅ�p��K��������ӧE����I��!�Lt_�J�nn�ݝYu�|�j�F�c+�Z�$NV�/U����}988�7������t��a������2w�Ń 	>��=��/����B��t��>�sgm��1آA�<�`'zR�����S����f�^]�Bz�,�>U:����G��`��1�|�,��(�
qU��F�u�����*�y�����XP�����ЂE�y�j���r�E��1��7Fk�{f�`�\Ǻ�.�3B�,2�%��!3�� �P�DW:aH����8���	�ܖ�D��8���7����32F;��}p�������X�V���p)�h�=KSd��6�g1���\���(�h���v`��I�����1ȉ��Y�7IRܩ��(Lu��)%<�U����M��Ԏ��T�e�V:�����k)��0!]�B��x8��[��"x�?9T��'�8 H�B}8��Ղ�Ε��I-db���#�>�꽯b�Ӑ�IC������Ԏ�󕿫���_��x��dH˥o���]��C� �帑B(ް<���먚,"�s��1��EE��K��u:�h�%e��)w�'�YI�F`S�f��ϟ�6�n�I�I��<KA��'�8T����N���= l�`�biu�|.��:FL]���ЈA���ư2����9@K5Pi���3Iপk?��fJ�H{�L-�5y�Fp���=,���;! IY���я��Y�~t;�l�O}����1U��F
������g[�/Zɡ7&qfa)��sx�=2t9�QV��#����$Jzد�ͥV�v�Q��{u,(Q�X��^Ř~�hh�w��5xVN�R�3�'�^�&?�4����T��G���T�/^'O��%Ǡ�e`��m�IwM}��-�w������x"�
����e[�$^�d�/�挦�ϜF�\ؔ���~m�X� ��*Xr}Iy�T)��zȫ��$'��Ԫar+0Kq!��YJe���I󔊍��)�����L~5X�&T����E`QeP��9�ź�`��ˢ�ʙ!��:�����{*�:^��ǘ:s�n��@KJk����:�U����إrr��9׾� =��UF:�|5�7>x[��.�֘ʰ�����:����-Ol]��|�L%z�}z��ܼyC޽{C>=�����`MnrC��?�}y��9�����v���/���zJT�2�Sy��{�8[��j$k�o_�	&�Y�4T1E��?K#� ������;�OR;���e�\
�#+]�����`�{?��ܝ��	q�ά�-u�^:�����*�e�L}����>��|����l��Y)2�{
�޿w]޾��ܘȍ�X&�	� 2�7�Fyb�6ـ�r9�	TDwF=�`�rb͋������������!m���L���՟�����߷��[����'2����������ٛ�����v���o������� U�,NڑV^�=�E�r��X���_�0�Y~D�a[~t��=�xQ.�Ǒ��O���u_&��z��7�k�?�����\�|I޹���.��LƘ �pG�ʎ#��6��C9�6:u�i롊V8�X�k����l��T`�A�������	��?�����E�+Z����ڍ��������;3�;�$�\R s+s��������@����^�'F�'n  ��c�8"�dQ�M�*��p�v1^��'@�G-���p��P���a}�ŉ��ɭ�K�X+�:5��!��a�9�y���K��W�U���)4'�����Д��p��P�,nwCt�K`���h�Ax�G�{�$-�/����rr$S �=��\�X�S|ʆ��H�=8f^@��F���`�g1�����G��0�A|��c�o�|�ճ��V��C���r�B�6�o��Ӆ�Xp��� p��N�x��R+�e�6՚��̌&�qva������ͅ�7��ʃ�X/EF��sk��e*��BXs�Wq<ۙg۱x7��kśR[3�C��E}�Icr�Ѹ&�d-� ��]'��I,�hV
R�pf&�SEKG�>$)�����HG\�����1�٘�g��a9�ޚ�
3�e���`��3/�)�x���ة�8]S-Ç�ʡ�ڿ�f+ؓ�l�s�xN� �F7�sUR����hM�ق��2[ɭ[�e��g��~������ܯ����d`���O��z*�s�is��O۳�{�(�~5��J����p��!$��h���i��0������y����$��C��c��w����`�'�;+�ٜ�P�>::b��T���#�k벵����� }Ǯ�z�O��2��^�`IVe]�����熓c�/�꤁�O��x�%K@,}o�"s��Τ���_���GW4�_Y���h;��g�9fV̨��,�gdV�Rd��H�������nH-)]�6�ʝ�<������Wdy)��h�0��&����t�Y9�PZ�#=�	~{v(�\sR�Gs�?;2Z�1'`@o�\{���ʎy�G
b���e�v)����)Q�u��ʣn<+���{Y-/�<��9fUZ���]��T��'	���U�G�,��=��B�1��:
��:��dWn��#�M�rw�'��-{G�齃3��a�A��R6WA�����W_�����Uu����un<��
�[ۖݸ&�;�䰚����c� ���Y/yS���vh4=��jLvIkcy\�Zg:Jf�V
�@����}�v�C���8�ʹ�mY�� ���w�F�<T?A_Q v�X�����Da;�U=`m>����j�f5���c�T�y��5���[�AMx�_������_#����ek06!,}�{��|�;������mnȿ��?����e}��a�������]���o�L"���5SP�e���oB�?Oq�w�l@��t��&���y�=��ƈH��5�\$մ:��Y�	����TP�@� @�f6��gf}]ўsV�	��{z6�f����E��Sr6S�9�(w{Tb!��P?���W���O�r����d��)z�����'S�3�ǒ�:r:k�g�db���JRV%�� ����^xք�=�w-�.�=�@��"�����z1�PԔ���-*�m���^:b6"�x��e�K]F��OC\+�ysP�LH7-K��W�ץЍ5ef}�ӯ������{�rS�ꎂ��X}2��2�����(�~J�7�,!�X�s�6B�{�C�ނ4�(���9U,'R�dx@�CZ��[ɻ1h�0Ȇ�y�#������C����u������	�yc���䛟�n��X��J�@��H�z���&����.x:�xL�a����%�5��AM̥)��R�S�_�ֵT?k;����r�\���[�.^$1;����:���hhi5#�
[Nu��'��m���0H��H�a!]�vv4��(�D�<����]��ڀ�`0��[xMσQ[��.�����>�X	�ua-��U�K�*�@��X�s	����Vfh�����`�a�G#�'��$��3["��ɻ�o�L4q��K��WKֆo��,�@�i��o.,���	:`-��yf�N��[q�z��c�+uu=8bYߚ���@3�Ӏ�Q�>�6��~T��]��LpLU��wn���x���XB}A��Ad�׷Ʋ�orB�:Qb��U�W:F!����^(HC�n ��`\t�&bf��~��!e��\/�P?�T:ԩ�9&�fd�ӿ�j}z�0��{��N'�����g�B7yF��L���,P���.p�2k�Q}�:4=�9�[�w�{CA7���7��ğ|�&kn�B!9�e��X�S��2T[�2g?��EV1���P����S��a�[d2Sgk�bs�K�5����է���sL�#��qIY; ��#�	�y�';�s<k��l�bLd��l�lS�G��[��H�����z?�B�ߑdE9�jQ�9[��(�p��sٻo���QO6�o��t�7�Ǻc9��ɺ��7���Z�i!W��~Y��qY
}?�!���Z[�LΩ�8ھ��e%�w��=�ӎ�(<c}�l3I7��5���ʴ9�IR��G�w��O�^���Ŗ#Ya�g0�С~k�����째v�ܚȿ�(Cd�s��B&
�O�="�8�+��ब��� ?�~��g����a�Pdm��B��{��4��{| 냑>������<3R)��X�k���ܻwG޿��ƾ���r��U�7���+����ɞ���{���)��uCsD�X}�юCl�=#���g&�)��ֿF&�O��nמWYօ�����< �iC$�G�m( zp}�|Z���
 ���s�Jn��.��w݌�l6���:#{a��+�r��;������bVrm����r��:'���@��.3����ʴ��2~IAFw�$��^w�^�ea4Y�=:�M,(T"[f4�j�*�^{�,TvA�&�'%%�:�,�H�O'Z�df�1� uxM�����[(P�� �@XV	�ǆ[��,�0�s�u���`�ˢGfʪ�ԘBK����f{ơR��"�g���%{}���9�O&��c�@}&Ty;��*�`�	���(q��&�z�v������l?�z�H�
2=������
|���K��c�E>�#���iA�Tӕ������2���d:��	�1;�
֤K��c���UC��Z����.[�{y�RYh�Ԥ<9�	?7�#4��A �V`X�rUݴ��f3�V!�\�9x���b���)��U[�t$7�W�hm�VS�0�$��ѩq�d�����h��q"�B=�E��O�9��^y{�P���d��{����J�͊�`�BWE�b��#}D�dH�L��bj�P���Z|�zkbA��\6u�=;���~c�Z�B�vˍ۷�G�?sV��5���5����ܢ�D��t,M1,�*�a���^m�00���)��8ؕ��}����s"2X�V��ZX�=�e -����jӼ�	��A�:�?���a'�ڣZl}%?;��C��eK����3�(�"^'X��6ʮ�mb��,X�QH��;잀���#p��Z@,s_�����;���' \���nL�P��4�_�����s�v��?�y!-�%xd�ʾ����J�ԭ"�,�6
�R�~Η�0j,�ڊ~h���t��>6�N�QRB�ͳ_!C Չ^]0#`�$Cd��\�F�E�lP�'�~���VtZ�sd�(�D���g����׾!_;{�},Q։,j����.r	9�Nj��]��o������7{�U�����fC�
v_	�D�����ÀIҮL�&�o��N�+�z]h�z�DHVK끣�:\-dҳ�Dֶ�[�Ͼ.Ϝ{\�ꧬ#�� 	})��@��u������9��V���1�+�D���{�l������xK�ٻ�V*TM9A�MI�~藶�kl�l�&b1���=�v�6!6�y�qZ��Cu���V���^���7�w�e/R:g�ޤ���̦�/f���z[�r�N7�[Z��w���m=G��BV�#������y��(b��7�c��ؔ��v($#�jxՉ�7��o#���E��d}Yl�8�E��T#b{����1E�>O�=�[T�G�MWUNy�j�(n�= "�)�'YĐ���DU��G
LY�D��ӥNa�{}A���Q�<v)j�T�X��TP#P�w�Tr�_ (��E�jy��R��ّ|��'���Fg(���	��;�:��G�N欁���2��*8=��o'� s�������T�P
2�������hm��k� �iHs،�Y�G�1��t�|#w:((8��^�}��W��FY�F��(����m#i`�SJ&��R&(c���tFyoZ�s����)Bf5��jE&�P�����xЫԯН1һ�V�Q��}����"g�&���>�����ӉLJ]�@�����i��2� �t�}���/c�>�Zx�o�Z�Oe��b�t���!��W���s*�~u�yF^l}�)�t�>.d
��˸�q9e�j��7��ep����b>���w`ە\���iJg����&@��c�6�c��C��'���M�D�kʁFeu���:,����j��s�k�c4Ƃ�Hf�%�W�>�*��)�T ����hΦ�>Oi�beuұ���Q�0��"��n\R{��lJ��V����<�uV^:��\�</�7����3�uf�������ȍ�u�|�<��U��u��v���q;8ܗ7�|C��^�����D��G��'PY�1�os?�m�bYQ�8wp�n4�&�Wz��X��>�h�%�Μ�2LQ4�׼��u�nTE��z����3Q9s���h��~���O����Ȭ\�3.�`f�����8�}{�rie��b�;
���=��e��$'F��d�͛�7|��Z�Ѐ�C?n��|�NXDk���z�<,QX�I`�?k�aa{h �`r����s��k�r��M˪5�C�`b=�,�h{9�*hD�tԠ���
�k6�F+��1�e��Y�S�Md͆�fD��Ž e(�=s�_��9���=�9ؕ�������ѳ�m@��to�$��9w�"��0Q��h٢��[��V���;dB��.4d��
@�
�V	�>�J��E�+�訳���*�tfK�s��e[�u��c�C�P�Sg��7�zQ��a�e�5/���H}����w�r��y��PzQ|Χ�2=�k�$�,��Y�aJ�y��ل��R����"	%̭��?�m�!|��N��\�65���
�(2�ǀͮp��uj^i����R���0Y뉟�$���ڷvP�
��S��}�sqWp�+��� 9�^�Voڑ�NG6{ku�m��V�rw琠��/�>2�#W}��$����@�^Vz�v�I3 ����� �+��V�e�:�䣥�hӉ��l�g���}-ІmXb��:N�!�d�0���e������dZ�@�a�3س�,�m�Du�G�\ `�����7�j����}�u
yor_>��Ա�MKYSK3;<d��>Z���
jX�Y/����ׁ�>�w$�d��,�F�S̺}~���`�Ե������4�lmoɅ�x��?����\Yf9�z��Ob�(�r;Y�����0gP� �(�3Uㄔ�{~�)��Fz^�/d�ʐ(�f}��ce�X�?�M��8����'���A_�~�I9��|��x*�^?N��չ�1�����[� +j�# 4�.M�4k9eu~��Э4����11SV�Č	�d<ʎ�L��E� ���QL���*�}�w�ЀR�ϐ��l.ѝ�P�Y����ɐ0`Sof"���JX�Uy��ʲ( � �lB�lP$�K���=߰`e��HE�<K7�2��S#���~7�����"�ծ%�07o��l���N޼�:�3�u�Ƶ-���aU��4;�k�����|c
�
.P���-݇1�eՀ�t�hv��GD�Q:����e�QO�ц<}銬�o�O�y[�ݐM��a�?�%ݣ��Ɨ�,O����G�y��tW�}����Y`K?�����=̸�ڊ�ګ~N��!BP�w�����45��گ[x���=�p"a@���I>`=u��������I��(F��zn��`� 4u�R�)!�j�Gl�����~)x����8<�U���.j�CKԂ՗U��?���L�(�Fh��B\d��N7Y[+��ָ�m]A�����xY>�<x�Q?��+oyN���?���G˦AYP={֭�&�o��fѤ1�^4k�e�5
�&f��0�jp���\Y�z*'@�_A]J��@}O�ud�B��PQgP����A�.���W'=�p�ޠG�򲗳�*S�
֣F��qi�k���~�t9�?����{�oIO�o��Uy����|��7d{��lq(�G��_�5S$2�!�H��j:�����I�D1��ˈ�X�����j�*�����YY=%O�[]���t�j�>A��:�(��K:U ������YC�Cfogv,���r������|����8��)��z����p]�㹎��U������ɲ�B�O�K4��ĳy�`AYY��.6���T��a�/
�k��cʢ+eVu �rËV����������ıA���t���I��=�`=����(�D�^ٟMI[\2ε��`	Z_ }s�WG��b�u�,5�Vċ2d�yP�"���g�̝}�4��.3�f$���}c0��N�g�,�z�a6u�"1�R�<�C��:�ݓ���rf�6����*�H��!��f?Qw�!�@y�~h�惮��޺�;k�� �!���2�k*��ʝa��H�� �U�r�G�1z扉S囲5�"��@>޿#��c�mmJv������ �`�!���P7�ɭt�tb�+0��
@Ǵ�$~�}�6�>�Uא@ĚC�,<+ N����M�ݚ�w�%3�F����3�P�07���GF_�h(���S?!�Jun�u��̓0��!���M�ӕٶ����zq��I*96��
��BH俌��{,bf�cL�į Q��Tt��C�uu����%K�<��i'����=�����DaX٨�f�?+��z��y�vj�׼���Des�-G=-<:޾6\��v���6�g��R�	��q�8@?ҹP�eC:�U�R'����h��	"(̑<��`��2G�ALJsLhճ����*f8V���o!��\� [U�K#�g��k� �Y����_��c ,�.VxH�0�����ml]�k��y�̞�1�g%_�g.����`�]U�Wt0)"C�$�(��r�sO� (8;���mY�ؔ��yO}ȅ\9{N�})�ʑ�0wn�|�<Ygd�uz�{�(迡>� 1B��9i��B
=��ǅ8�@,�r�A�y��²#�]7kEv�����j�{`^���&��9�1+	�r��y����LX$э�wMI��pbԀ�2��VV�Vz�d �E�M]ac]���%a����Y�gMCZ�-v�C�{�$��Xõ�Z���J��'�N�o�X ��{�M������a�/rXF"�A� ���u ��׋.6(�Q�Z_fP�Y#���R^!�����>jk�	d8�3�S���dHה�jQ��,���nK*���ԉ��Z~d�z� �5��A�B=�MS�C�q�4��T#��1VgwCЇ�K�9+�Ju}�>�b=8��`�ʓO�����S���E�3Ra��<)��\��8Z/j���7'�N�#�듰ZH��!�2R�m�ʑ�+�֠��"K�z� ����h9�y����{2��p��������`���z�3���e��f� ��ę3���Y}���#B���YAEsi���u��EsD�sh����Ɇ��vxS[*z:�+[s�(�5�|̗|�Q��b�I`�!BǗ�G7��g�2=�$�asB�u�˝R��nn��
+��u�}9VP��J�&H#"Q��9{zUVw��[�#�Kw�yg�©P��9��+HR �G�]��)`�яM�Vok3kef��`�;�CY��jw��������PZ- 6숬��#�^%��\磮�`�Hv�R�;R�x9_��}�7內���ںLS�?&�H���z���#���尘�L2�-� �+(����u^��կ�7��u	
��/����?�C]�.�� ]Ŕm��y�t{�"f5���0*�g���h(k}�� nP�D&�M��2Q81`���fG� #�ZoC�۲,6����b�TQ�~8\�{O�l�̓�(��F���lI����JRέ�R�,��Tn��>s劂�.Ӯ�	��g�V%9�́�2*.�N���X3(��5��D��u�|����?�؃�b`�E# p#hZ��l���IN�z?��>N��!����rS��f^G�r�T�y-�S{�	(�I�I׾��)%���F9&�{�K���l
�$ڭ�)���<)���N_2jEe�Rd�Q���C� �m+z������<�k�ߦ�Jso}�?U�>�=���� z�k�Y��I��`4��ӄ��as��\�s�OY�,|Sg�j�]I�Hb�7��f���3�K�g�&��%k�;R-t���[˭~z*����9��=���E��U��'W�D�d��-{b1��(yP;��G2���=M����U�{c�ӽa �z�̿��ߕqw��u�Џ6�e�`_��Ʀ2�#��b�:�u=o�}_���j	 ��Z���#Zs!M��5�n��>4�ʾ�]��ב}��9�@[H �m+�q�A���t�%m	��KB�	t�l�e�'e���P��Ba�l�O�0$�D�M�ꇮ�G�ʴ���hc���J	��uוOD)��P��F�7	Dp���7{�tlcJ�%K��U�{�]�K1mN��39�������!�г{��OpBٴ�:J[>��*�\�f�@��!z�C��>?\���}�j��\{_nܿ+u�@�?�O>��W2��2@?ţ��>Ek��5��8������^�{�fuZ -�c]{�����c�%���yOx��$eܠ�.�{k������l�t6���xf6���}���Si��)w��--�0G��9 #ߧ�E�u�����P���iN���r9{ G�/v�+� ��H�1��oNƨ�>O�E�(�5�x]�$yh�xݨU��SRf�@d��0�lr��c}���lx ؾƇ���"j�NU�}��oS�����T�f):���^�u[���PP�Jǽ7����eSvw�C�V����)�T_Ӎm�f�p�3m�ٷt�7!Mb-�(�Hg�T���ei�[-"��qNGE�˾:*�ۈU���Y�*�J��Sև- ����u����*yj�|���uCP }��t�G̶monKW��ų������P��1dY'3	�R���(�~��֫�˕ˏ��O>~Wn߾��ݮ5䍠��m����ʝ�huz+_�u.򄂦�ߒ�g��:O$s`,jZ:f�Q�L����ߪ��XZSzD�Y�-[����C +�ɽ�����}���x@rb��עx���������P��*�}B:#LΌ���OȠ�e�"���K,5��t������F'X�E�����֩YE�����'�é�e����E��LJ�Q�Ԕd7£V�/w����@V�.Dx�y��i�d꟥�5� v2�a����K���P;�5[�Wb�=(�I�e�_�<�P��=(��PY��Smv.�>Z���0[ȹ���,T��L���ȫ�Yq]�E����(�D*pf+Ϫ&0������V1p�N=��S�g��G�{D���%G=H�M?�|��S�GEI{zs�)T��RO������b4<�}�w�����m�Wh-���ͦ����G\]���o+���PY�
��9�T䠨GkB<+����LaIEQ���p��=	
�P��y!�_���Ygl�f�j=?�����lno����׏^((�%�tD�3 ��Dj�x�t����X3)�=�vB��!Ù���޲cJdx���q��Ȟ��j�y'��͏��R��y�iy'1���������9U�_s2;�����:�'%<PC�a�+�s�������r:�Q~�\~�c�!�<L��m�D �X�{��6���7Tn�q�6 �e.Ƒ�F�=�J� 4O0���R�t@r����_B����l9g�2(��#k���>�vN�|Dg��xM�����/;�	��я��3��KW��'���rgr@�e_�W^~R�y�9�<���m)Տ�s��ؐb2���9�*��s��[1�ͩl����HC�E ��]�/l]���xZ��țw?�c5�[���֖|�g�����R Ñ���?.����뻷>���}��B�n_�s[�k8�Mx��F3�u(�2g�>��&wt�Cju����Mc@گ�Wd�O�U^�Wۊ(� B۠H=W$m��Y�MHѬ4EPW�U��"|L*�Jy�Y_�1��y�����s��v5O��=���{It�P��v���5���h��|u�G�A6��B���Bj�#��9�\eF;.+Ϥf~.�mT��t�of}�s�:���d���&\�:��!NYf���Ϡ�@Z|�lF�ʖFB�CaLH�w� R)���:��U�iY�� �2*��s�@��Oޔ���A
�N���o�KO<#���ߒo�ַ����u}��k1��v�E�����-��+��@/��O>���c���ޔ�v�X �(��)�σ�A�װ�r�H�'+A�ڮ�
�^yB�+sDFTg��ʚY� ���Be���Fˍ��E��h��D�2[p���O�c�YA!\��r���M�n�Ր��#f�#��P�k����:�:�۠7��U�X[��#��Nu�3@MP�}Bf��Xb��5su�h���׋�\O��]�s-3��u
�J�KS�۪̮���-�����X�2�g-ܴ�����AK�O���yϊJ���Q���}����l��-�Q�`�`(�����K�M	DյYn�eI�4_��8]	6Ym�k�M�)c��˃8�6���j^���6ߺ- Uz��2S�24X����ֶ|�'��G_�J�R{�Ӭ�Ʀ��0LE��i4ҽd��{�=`�I�$��Ξ�S�[����A��S�t�O��tT~E�MQI�~�x@͗�^�tE�Q��"�]���w@PBk%2o��ۗ����*�͐�-������x]ƫJ@y�Od>=�ը/��X���6o�얜����Խ��O伂�E��g_zF�}��t���5�{8=��J������ZJt�V��f����c�f�+�5[^�) ���?��
x�i[s�][�>4��i i�����L��n���S�Q�bt��T�d����ڋ�WIx��>��y�n�Կ�B�<���QG�ҿ������(��Xd�F*�"K%Xyq�.!�A��`5Rl� ]�
vS��7OmFB]X-��5bQ�#�g.*S�D�T ��7z���7D$�d��:M�u��+_�'��̴B]�@;A�ܓ7��'��aբ!��
�~����`Kn�S����'��y��?��_ȵ[7�A4s%�ɱ����PZ8��h�aƠ��r<`d��CM��hn��o�P��8'�	:N����Oߐs
^�����kߔ����S����H6t|Њ��O��_~���p89�7�=�����7�U�t�	*Wb�ϯ�������[ׯɮ:��a��������f=\� 4Q*�K��c��_�%Vq�F&�2����Ʊv��`��+ϛ�S�*�Zfd�I�q-�ӪU)OFKy��K�g��`���G���N��ԘnZ�Y[���1ݟ���չ�_��K]ַ��V���%7Yh�;�z���{H��'�5zU���=�4̼�@�� m{$#u�g�g\|���$�r��ڸV�Y|���dQf�CЎ�f�zIj�@���q����v:��F'X���s��$�o��{7�K�1����wn�o(���s�>�ȠQ������է����ߒ'�?&7?�D�{�]y������M�WI9�ZI)s� ����/�3O��TT�������)�BD�C��Bn߹'���1�t��e���\�y�f1pݰ��ڰ�L�
}Zh��+@^�+���.�V�������X��U���Ѿ��xG��3S0����$��yr�LlŞ�〚F�{dX��NX7�˽�Su좜��d���ﵐ��8:�s�j{�uF�٤�*mt�q�Ua{J�#�שeUY��k�i@E�ru4鸰���.�DɆ� b���,�M}����+�\���T����''+$��ʀ^j�u����S�"���.O�����A���1���9-�ϸ��v��=~杻}ݰ%@d��%���,�ݰ���8"A�1����y��>3�!�I/f<�8M��x��N<��Jv� ����p^O䵾�C<���?g���}�o?O��ßi�N��b�4~����:#�<V���r\�r��=y��k��:��Ռ����U؋&NB�__~<鷈u�Q�"u���IE��d�U_���
Ob��IO������JgЕݽ��H]m�7���c}����y���t�o��uM$��<�(�V;�}}�]~�����F/T����ܚ?cڵ�?��IÐ�i�܃��t����im�.�
����qxP��M ������`{�/zͱ����*�ɟ�{���[9��ns����=����$�B�*%9�)�P��Eb�:14���%�VR����׈��Z8���e'�O��B'tV!��Z2�:쩓��&�c�Z2T�q�Ȗn/^�����os֜L�y�{�'o|���wtO�6��8�s��l��G�/M^}�EyI?wɦ�Ȇ����;�W�+˵�,;h��UGe]&����gR��ԟ������i�66ѳX5!:�΄���)2N���|�	x���U7���^��ο��<T��/����/��T�W�r����߳���|�k�}��g-s�7t������^9�&#>]��eG\���s�lQeY��e}f�`�qobq^3x�B�yH�ҽ�V5���,f�$�Љ,���mt���[q<NW>4���H��K�������i�zn�k/2˔�9Y����X�WJ��&���9��#u�J����
�?d�PcX���Z��{��	�T��}ݢi�qCɳc��=�K�0��BO�
���򭁌t��
�Ț�F{��eM:bJ��z��@%X�o*�Ki�\�q0�=s"
s��+�PE�x<�n�~��� ��Z�ڸ�k���^��\���M��/��wߑ��{A
������3�7_�5y�ٗ�����Wo�X_���.�e� *�Y��1P��LL (Z�	���8�ƮQqS�":L�笵�TIF�Od>�v�����n��K��'�OΛ�^�����5��'�jgևc*�,t���B��8�3k�Mk�v?��{������;ȕ�ٚ���LϱE!�T_J9{��Úp<����Xy����յE�R��?��H���>���$`�O�������=}#:����i�֫�*26ڦ�y�KP����.g�n�7��k�#������u�����.�{L�g���I�5�L�h�� �e��G�\Ә3ѯ��٩�����[�&�aʢY+fm\IR�ڦ7-����o��%>�@>����ʆ5ʹ��K��:\6�6��@���t��J��
2��r��)��
����ܮw��lc��b��Ő��>jZ{P�{�lՏ���%�x���h_�ϏG)�(΍�o�2�v[?�\����w��4lKg�̀�KW��w�:���v;�C���ୈR�63�.�ZO�~q�h�tU�q0�Me����y��1ϛ��`d��C��P�7���AGn����D������E��'ֶ�#Q|0���l	��&>ݚ�m��֥�p>��3��:ܟ3�J��5�W����5k �Ck�Ld������X�/f�������~Di�H��t�����4�)���N��A�X�ӓ 5��&C�Ј��t����;{uvP���ĺ@�Λ(�6�+i"1���Z��@*_b�s*E�K3��`[6���ں:���r)��?���K`�&��� �����l"ޗ�y!G�!��@&˅��C�<v��g�Ӷ���Û����[R�����ځ�s�f����ym����ڑ<<�5����`'8�o�	y�JY ��� �������Ո��}��1&���Y�[�D��a�X���w���;̠ ��Z��{��\ӱ8�U�]W��j�"�
�9F�!�ꨶ�F㖬�\x/�T���
��}�1z+[�y+����Ǧ�%��֒��_��d�9���Xq��I�`���kczKj�KR�j�Q�f���	DW�Û��aoi1J �i+��#��gV���Ei��������ȠpÁ�ƝM��}��,���k�{O����3)|����ee�c�zʻ��A�](S`C]���<�rh<��2J˥���y���J����GZ�tɽw)�!� ���&�\O�:�! � P0��TÎe�!L���:V��\��ҥK2WGb}}�"JW���o��Uy��SRN$(�z��eY�dwv ���H>=�'c
֩@4����b]k��w�QO�g��Z��ˡ6���������}��~}����墐��]�|ᒔz}w[����F�����(�iŌ �,_��vI;�qvK?����"%UL� �,�pN��KI"0m��&0����>�X���-Br�΢��-�ʔT��;#��y�{C֨޹wW~�ӷt�5���i�+������3>�2(A���k��I ��Z�P�� ��:�WE]�$*m�j��3�_���v��iy��¬�v5sP+��)�n�u�1 i 9��	�I�9�P��a��N�)᱿僲�k�-Qj�Y#��y��pj�
�7�O䘰gm�~m�}s~����>�-���s���Zs��Rzڹu��������'>��y��O̙�/{��}
�~��ӿ�f�#=�Ө��B�}go_��ɛ���y��'���Kr~�%7nޔ��'����J�����>#�v;�ZFa6w���X��W��CB�R����B���� �����BHQ��@���ֺ�ԦC��p-|�Ws��R�0cT���5Sg� ����C�4�j�L��bN��v���5K?�cQ'eۀ��Xb| 6�ȏ��ܣ=}��j�Fc1��c㿝�uwzX^wJ?�<�)}p���s�鳸�L�R~��g	�<�x�3��r�
N�4�e=��H�ଢ�\��)+���@I��;ۿ����o�i-�g�h1�Q4`/���=w��ԽY�%ّ&f�~�-���=�2+k�"�E�\�PH3�@����~ғ���?�W	h#hF�e4��4�M6��&�M�^�����}s�#��������"�l�-DEdĽ�?ǎ}f�}FPrws��6�LH�PSv>���z�Ɏ;��]�������?w�t�h[�¨wZt��g�`G�A$�X�ͷ;/��>�%�G9>Գp-��#ZZ[�p���Z<�fp�-5jM�Le��4e#kc((R��.�(]�~�	(�wFk$�rQkU�@O9��$(�͌6+�FA�0I��Ǉ����mD�����)�p<�v�A�<&#v�G��A�R�"�Gt��$o����
L�8�&�_v�z�9����ܙ����;#�S���>1�ل��ɘ����h ��V)��F+Vj���j$���Z�;aJe��6�<�v�"�(�PD>�2j42�����g���FS���m�,B��vb�ʉTjt�
��ک|��O���q�#�h�7���:;��x.u�ȴ��X�g� M$� d`QE�9	0᳨��@]R�X������&ew��R@ͦ�g(��Qg�`����\=�>UU�Du�B�LTi2�P���KTe59���Rn�5����":sV[��I}�R|Kfr��@(�x�δ��f�ТA��gԼ�xlQg���2���2�B%`��{���[�_�7.]��������ƕ�r��Ɉ~�џ��Ǵ3>�9�
�p���l[��Z�͌Yj@W�i������� �p�l6����Μn޼)B`Aw53YS��tHm��u7�
;Au~�>O-b��K�̀��wz�s��j��X���D�BV r�s�\+�P9�I7q�G��#�}���9u�PL�^�)P��Zl=J������۴�x��~��o?���.��
ɒI�N�`�r����P� �������� 4�P��b�&fi���Z��\���3�2�V�-���} �;��)�9�^B���?����R���1���YG�����7wrߠ�y�/SXE`K�"��W�oKU5�?+�$Y��vȞDU�!��D��A��������i�����gN��0��t����OU�T�.{�)�M�9/|���/zNϟ�K��Nǂ�Z���j�PM������G��""�5Ƒ������gx�S�\EZV4�%ßZk
�a�flf���c���ǟ��S��|�f�Z��--1 �AE�X��Z�9Cy (���e��1�E�շT�3�O��	p�V�Z�L��Y�"'�z&�bv�9O� 
_D|���'�w:���l^'��O��ȷ 
��^�J��և��v(�=�����N���=�>݉�z�8�IQ�����?�����5Y^�*3��!��dVjeYHeP@�,�$� �'O�����l�x�ڙ��='߼S��N(g͘E�Aѡ8`#���Ƌ��ړT��A�d�ԡ���` Ҡ�זh��V:�4dG��_��i�����?�w|@��H�;�$�X���|�gVEɱQmH�!'�i�����ۣ�<����t�T�z8ƥXE5b�l���h�S�>��EHIj\@imNb�%��H����,V)䍿ʟ�����S+~� iHkb��UNձx��7Ҕ��ڄG4'�v���B��kmf	��`g2a��z�Dh�F��c��}��A-b h6
͡Q�=u3�B�A�'(�KF'�Iv*`��������2���h?�2��dNR��ZFP�'� Z�R��F��Ӂ�<	D�/���7b 
�t�ׂ�D�xF;�x�cP[,�MF�$�͛N5#C�17=Q .�,�HS�3*&\<w�+U5G�<�54Ud��?z&W���:�>dip]�9�>�ti��%4�Ny�Z��7u01�ӉV������C%s�	\��}�?rމh��5'�V�@��	���P�����F�1x�-�Po���xjM`]��#�����P�:�e˧�����p�Q%fÄ��::��J�\�A�'7^y����ߣK/ӓ�1�>ٕcm��S����}qN\�"�r<{c�t���>{�F㮬��ȭ�B�;�Yg_֬Y�>�K(��Di8әF�%PQV����z�������3�%��s�ɀ+��I�ɿ���Z�k����	�v��6L����8��CB����ċ񕚈�e�-Yk/����uN�M����D�)�
�g�t�t饫t{�	ϥ5ؖ�__�o�����������
�]�e�Bk�ML t <W�a3��K�f�Q������&+"�;�)�0�&)t-붟�zg��Y��]K5�`��k=n�'���Y�3�H)nZ�,�^C#�/��~�ٮ���XC�r�A���A�"$�5��.��D�4�γQE3[�J��H�S��|\���c]�M�㛄�w�9��1o�ҳ��9�h1@��.��8��+ B�{��iFt�o'r<R1����x�+p95���]7Z���YM3���v�'��K,�;*bX(WA]p`�(��D`
es���TE��d���	�G�&$XVo	{��ו��r�#������:�޽�⟀��:f��gf�{#�
��l=(�������]��E��Q���2�s쭱�������L�\v�H���� n�c�A���OO���f�Ϊ>�]�Y<���f�� @���	AhK7��*�F��D�?
 ��l�Y���Rt�SU�mq����^���U�ȫ�J��M农�S�<
Q��S��ǂ�i=���\�?pg�9�BnH)3��F������V�m��jB�3�pn]�s�wG�4�zP��@��,�$�� 2G������X��I���>�I]$�qYD�Sȼ��G�s �2��=KvF+N̇l,6+"���Y��JK�"�u�=�9d�&l$Dƾ�Q2��B��(�@���DL��+�4��l������_�h2�y��ד�f
B��� ����I$]E&B���{�kͧ#q
����z*P���Bp"��>'8��0�j���݀#$ q�P�1d ���W�\k�d��@
�e�%�q���3Ǟ��$���(}����W�(Mz��:
! U6�Qh}�P`C���b<�v�?@&6���٪���2h"�����D6�PG]_Y�z8�<�"e�C��	a ��)��ݦ�}�!u!�o�̹��
% 5	 ���O�7ݵ*��Ȝ/݁���%5Z>g4��e��:�4�ֱ�y�����������WikmC�I"��f�a0� �5�GM@�W82��Ov>?�df1��A��|�wg��_��~�_���� P/�JY�H�Ox��aL�TnTd�
�g?	�r[�sT[u�FZf���	�>j�{��69���d4\�֪���O���b#�<�k@�+9dA��2�?���k�.�$P�����C��v�-x\�o?�_~�1��F����4C��k����x���]ھ�� �)�CE�0٦f��Щ��FU=x%�Q�z[�B��I�=;W�Ν��~�����C�h�!�*��`�}N��L��Z4!����9QWj��� �ۈě(�nOF�%esH��4�@�Z����5����#�C�FW��T������6�D!wg�1� nln�ۯ�`�����?�~�.�J��H����#�0�;:�`���:;�e�J��DM(��Ҍ�tH�
�e̳�6�v&��e,��z�A��k�r�l+6LQ��1G~h�3�<���� ����%3p�|����^��z=/�a \h�A�^�Bu�	��{��N�	�3�2�T�k��4������i0褰��[�K+}6��<��޾,:�Ee����W��qEv�����:*��NY�/!�#-���_�
t}eG�4�G z�=?v:�x�n����{L��\XK2���Ly��C�G����t��A'/���4a����\pr ��!�K���sJ�DY�s΋�����i���{�MG�[@�e?Wd;�;��m��a.&石+� �3g1�R��i.i�O�2U^'#�;���"�"^'�=_$x��k~|᣶sx`[<�\��E�=����Q�� Qf|]���%;��rK`rY�Q5���q�\�7�dG}���Y��/1. 4zd����`���B:�Y/�9� ��T1u��
S'�t�Q����aO"[����5�XP���u��=Y�vq
v@]:�ߖ�`�tʎ�+P�K<hha�+��i�&.hb�ˑ9{
���40�Qu��D�C57�h>Ki�^iAY "����KMZ
k4:8��贤�h<�r��X6�MF31f��NZd���=�a�t��ی�LK4h��P�@3d'��V����=-rA.�F>��7n�q����{�2��"���3��tc�y���@T���� l����UI5�palc~@f�BJQh&�P�qH�卯ӛ��������t<�JY�f�KP)��J��������wPDƇ]Z�6�L����ƽH�@�p�'��D���J��8{���Uj00�38�c���t�<�����dX�  P�G6Pϖ�� �(�9�R��B����T�tx��>��Xrc�c�;��X_�zMA?@�4O��s!��8HL�Z.��ո:�8/R���"i��F-���}�=�����}�{=�XAy�^�!(��r�o,둪�F���H�l��T�5��r�E�v�~�S�+
�A�9J���=T!�Nd��m�F`
��R"��$*S�}�ݠ�7��T�Bd��=�P�Z)	��X�֪4t��-C�K�M��y�@E2��h�N�m�<'��:����ޘv?�_��o�wܥ:�-�j�~���O�ݦq5�,!��ʾ~�
]�x�6�W���`J�R�����׌z������R�ڲ�M�w�fc��p�
��G�;G%:{�;4zp�._w�<9�k��^�q
��*?�Dk�$�0�y�HPNʫ@�c'=-� ��K��$yџH�;�[��<��b�0����;ƦVo*�����LՕ�	������K/�D���0h�X�E-�f�� ���v8j���|�`���э�W�ݪ��D`�T�a��4��]b3f�<e]�@N.���z9Ӓ�L\V�Q�7M������}q]?B��zBQ���c���X����n���io����˜�D�3�x>p%`�)���S>#s�3yᖔ�e�π�	,^KaR���],{�b��b6�^��30�3��ׄ�[����G1wf�E(�x�S@	��,p�%��1l�P:s����|��!��M��ͤ�;RO�)�
H������Px�;�}���F�÷1b?,��`DӔ���,�W��DZ�y"��j��������;f�� I�ޠ�ހ/!��hL�RE��~��-#�m5�05��5Nϋ��-�}��o�'��~�̽{���3ia���6��t0�U��I�}��cy��6ON�1�N6���Bg�M[�%Y�)g�ގ'~B"��JU���@�Z	e����d���S~�B)�	��-�SG��\8�	���s��#ޓ9���JL�a���O��o)�����:�"����� :���*�>�K��C�����s��y!��R2m��މ�xAh�è���J�A�:�����g��L�4�78�5$U�R'Y�iF�B����=:�_��t�x�*�hT����Ii%�	"Ϡ|1�1�P�p��@@��*Ȕ���:���=�����o|��mnQ�ԑ�-�D�mK爁Y8L%��P+��ux���sC��?�#�f��:;c�Ԯ�����[����l��]f#�Ŀo�ʒ�(�QǸ���36�gS^���:� ��|�x�H7��Z�D���W?���)_��UkR��JX(�,sq^�4�� ���,���p}e���L�V;t��V���<��h�w��{<W!#��`�΍�<g!7�ڦ�Ϊ@g"4�z�N/�:�������  4���~|x@��χH�
8��bFF}�D�{�i�7[�*�H�@���H��_�q����+,K&��s���+v3j3(AQ����pܓ��v,N�#3�,\��!��z|��>�[����<'**�.���=
�]�V��N���}�^���r�X�0КU�5,duLy�ITZ�  ω�`"���Hڳ୒=㱯![S�
��%JP�������G럼pLj&JE}��ꌅ � ˸���՝��O�v,��hΏ���6��o&�,7�]�o��;M�����}���h .�������^��a�<����u��B����2�A}�������4�욷a2�Y�9��.z �*�"��l�C�h��'N�߸�3������s����W۴�@#^�/\�����1���ڬ1(*%l���8T��,.
�9�QV;����@mc��t�A	gYk�L�2"(�J0CA�4�P5�Q��x<�����n@��� ��k�l�W�x.���������5�RW���?\������[t��Ez��A�u��hL��L#�V�ֹ�����v��p\	�E�:j���K�Ϡk'_>��_h��<�2gЃ��D�<�y����sc>�HyzB@e^��F7{=-��BW�:�(���;�F�,����^�WD�$儠'����1L\J�*(Bϸ��D'��	��f>�����
N����b��K�(�f����0����X��dv"C�g
��y;$���BYA�������t�Jզ�ܺs�=��4�@V'-�ʜ֒�`�A�>��rW4d v)F x:�x8f����
���U��COM�Q�V�y�B`�1�&Be�u�T�C��*G����mm����%U����4����T�s�������gg=�<�W�����=�$�4��LX����r�x�g�Ӝ����kȵ7l�������c2���ӯ}��$�B������/U�N�u�J*��(��l䋽�~oa}[�W�N��¿��@г@Y�i����GA���7)p��/�F�3������N�����U��np<���!m=�4����BSp�mB��YC/��TT=��Id�/�TU(��2�\��B�����
Y�D��Fk	U�@�	@ì��6��i�\g@�z�*��:�W:4d���O��N	�d\�
����*�}2>�+��@z�!��i<	i%jѹJ�ދ�F-�����5�S��IC�(�M�BsT��'�ڏ�n��u~Ӓ��6�R�+5�?��dS�O83�-6p�1z���Uو����ٺH��[ߣu}˥
�HjܤnHV=��rS�:��:`K��\@G�Ϳ+k��|8���K%��4w�r�at�Y���S�??)��p�!�a� �J|Cw�2�gו�!orp̍�O�V��� c��iZ��:A����U-3�M��S���|J�Ã�2ok�~������m)�>�}����>��9�v�y|�>�`���L���h֌�i��L&}6���p.�U3���hT%�5c@5	�|�D �w�v����� ɑ4֍�j�YD�pO"����jUǍ��Ck7TG��(0/�t��an���;�~��aC���sS=)���j?�9h��Z���Vc�Dn�hG��w2�J��2]�4V�q��ڞ���f#L%U(�8�2�V7(�_m<MS'A�z-�#����>:>�G�C��{?ّ��������u1x4<b�w@�޿C�7��K7^���}r�&����XY��V�V:K���=a �Pv��	1�6��ϕ2V�<�\�*wQ��x�@�1A������2TYvO��#^��i���mF@�~���b����K��\�����R�Yg�;e����x&*=%Q���a<1-4��1P�yI�f���4�`%�-6���&ߦ�Z���\��Q�e��6V���:��6mzB;;۴��F��5�A�u��ju+�}X5��Q 0�N�m������=F/��N@�_[���W��#yz[�-�dԨP緯5�`�v��p���Y�T�3�a���t�"(,ޝ_���~#s4���6`�B!���ߧs>��,P`��Y͡�%��NŽ��f�r XsT<�����v�������D�Ʈ�^�V5��,0ZTQ�}��O�����g������K�Y]��iwgG�Psi����ث�*5= �3U�8J���;|��pDU�������=i����\f��̶��6�.�&?�#��vv���.�w�G��������1 ����v'-�ߠ�b����������P�l��3�'K�D�-�T)�B�,N��y�]�a]�v�(|ѹ��i_�/O�N	(4���@/�.���9s�ɀ}��d�%��x��'s��`/�gE���X�, _;�4��L���;��2�/ze�P��'�_0dI�F���d���(9!���
�I;�j:5�F���}|�`�f��W��7���ɬR)5��xJO���xx��QpHM�� H�XU�@aQ��΁7��R?U'1����4�\�=*d$Lg{b�ET%�d)8Լ��FEz����k��լ5�����ѓ.@�>�7;����=�s���"
ѝ���I�	�2O�)Of8Oc��B�A1���Bv��A%RǶ)�M�'{'˪;���2;� "B�
��;lm���|o�:��Ҧs���.��2/�J�.j����&M���AL�i,��%>���5z��Fu�}���d	�u��~��\���4�3���hC 5g#�W�Mm�#��	'�>�\�TԘ%�v'�d��U���1P�D1�5��>|N2��, � �'��)ʚ����� Y8d�l��M�pF�Ap�̠5�Ҧ���m��B��z�JǭU��A�x8�)�}:�|�p�Hz��)0�}�5?Q�0�T�u�5Ӭ�]��mH��C��Ɉ?�(�2 @�d%�ٶ	����v�d��P-���Z��0_q�PU��ntR{C� �b����o��I�sx*kS�Ҍ&��x�z��68V�,I�pP�J�	B�u?��OQ�G|&�� �:d��5@FZ{����jM�>�%�x�7-���boh���TϦS9w�X~s�A.�T��������M��� �A�Tw���ӟ���<'��?����J�����vl~�ᯨ�ֻtfe���fS�u��{��f$��5�@�����kAd��T_\�7D�@�h�C���X�S͠,mB�v�;��m�Cs���L��ko�Mwoޢo^���Z�e'k_Y�X"���E>	:)�Z��9Y #Qv����b���B�v$� n�#lk����d,J�(3Pl�5#3];�B/�f�s���"�l?�F��1-�n�����p\���y�
C� ��� �WT�������,�vl-��d�k-���3�P��|�4�g�,��r��Z7�lC�e�:œ� '߫�_�EU�Ϡ,����8������-�A�S��,��g��BE��Y�U�z_�A�AQ�B�����9nϿ�0*�u���_���y^�̞}]º���#��s�� ��l ��l��g�C�����wxOE�{w���Ci�$,��ZC1�s�7G䗬k<��J`_!(
ۃu��88>�Qw �s��KWn�ٳ�t#P>+�^Z�:Wu��U��.^�Bw<�j�I���g�S��'�{�4����^�%���kx�,��ȋ�0y����3����%b�A��14�䤝yt�]�$�!\ �vN�T W��K����1#:::�D�P�0%(�k%��v�b_f?�I�V���[�5rPx�/��j�:?���M��r;]�'���S:����z,y�<§�ܜZK摐���/��_�Dp'~m+S�r����mٹ3����F��q���5��"04̨����#��=��ԇ!r,�)p���T��1���qF��<J������@)�6�C�A1:�<����C�p����FDJ�����]����!�G������t��N!�#���~O���^�y��y��s�>�{H��C��� @�!F�Gz���L2i����3� " �l�����2!�
�W���j�I[R�فy����qV���Mǈ��l�+���F��_�	�h͕�Qw�f\�τ����a�Xc YJb� ��S?D�ל�"D3��EYS� m�Iay����a�h��k�hI�+'j��t(��L&hk�D�=�W)ڔ�Ҷ��6\�����F�h�2�<C ��Q��/p��A��Y�ЩE��|6�1�Oi�V����4�!c ��������,�8�h�ɎP��4F�!�X�q�a����h4a�*@	Fq̎2j'>�����e&4:�	6�XW��!�H�s�	F�G�o�� �H��I��H�5j!�ө<�jiW`�44�E;d��N��a�&N����DW��f��
�䌇������`P�)긑�o�9�5�%Y�1�N�>p_�8���5!n2�>����r��O�;��Z�;D�i*��6j/���
���Z���Z�A8����{l��t�����*���da!u��c���F��G��sߺs��ވ^�|�ήm��?9�'{����;ts��N�4�����2�B�#3(�	��w�g�2UjU[Ty�`b�+˳=΀�W�ӛI�yb����������7�ޭ;�vn�z{<����G�(Iv4��3����w �e-�C��Ft�и�$��nQ��A��f8W� ��Y*v,` 9B�(�>O틤'�����PLf��d`�`4�*¨��K��1;���y_�����FOakdA�H��%��M�6\o���NK{�JM��A��M~/gꗩ4�W� q����E��Z����r72�f���t�Ɏ�,<�E�|�F���ijK���2*��h񅠈�pR�-�v�V7xt&n� ��¸�~o�?N��<;5s�}0�n��7��i_p��Βħ§���PA��\�/���Ѓ�_�~���D�Ǆ�֣�C:>:ҽ�@��;�v�v��"䂾]&���#�$�1[x�3�\i�����^WѸ��.����(�5Q?A�r�B��i��z�����>T��D��M:�u���>��2d0��Q��x��z*�k��`��� ���O�Bf����[
�@1eњ����\n?�Ng�=�^��15`)[�G6�i����~D{����v��{9|ɲ�Ga��^�DƸ7��b>��t�舧�=z��5ZZ�0VH���q���*^�>T-�B �$>���7�9���'(��$��w��`��(䐣��gN9�t�Ѻ�S���[�0,�ر�O'F-g]r��s��C�lb�爱�Z�f�d�s���Ag6�)9@a[�:k6������� ���A� j�1L��c09��2���˪(z�,��Qx��z��s�e�t���B���h�X�T�Ft94Ȗ�5�<Pa�c~��t����������C��<oЙ3g��5��\~3z~E�����s�vx�?@&� .ڠ�R�P� .@�+�*�g%R�u�8��z��ך;j���j���h2��h��Fk�V�i���AgWW�R���ݹ}�����Yn��p������耾}�ll��3J����2M��[�`�%�j��Ҝ�(j�E"�,F@�0��:%l����%Aű�gub���S��۹e�%a�@!���Կ
��P@K(���>��qrڎ#�gw�b���,R�-�;Y��^�#�������h��P���P�ވ���L�v��Ξ��s��.}�ӟ��ۣ��z���޻t���X�,��~�:
�q�P(� �+��)��}@>~�֣��s>�-�ײ5ǅZlN��?j] �e$#�ٜ�ρǣ8���]�����A�
�C$�M��g"֘(�Fz>D|QI$�S|||�eS2΁n��oՑ��
Ul��l�i`Y|&��t&�h> �kc�2���ҙ-ZNyL�	�eH��A+�c=�C�b�u�aD�G��u�����D�K��^�N�F>�I�y-�xW�	U��ď, ��ÿ�ݺ}�7��іg�p��C�]]��^�Z�z ��K��rU{.��joS���q���W_��H[{�y^����P/��˛�DP'F� �7�N�>�����-z;����g=��d�2�grom��!?wd��QX�=Ĕ:�bK�o�Q�+�r>e����PEĺ�"BD���4v�@|�B{OD�7��M�t9�����)� _�d���x���E�0�95"�<�z�nw*� �=���ei�D
���!<<<��/�
;�K�5�S^wN�	�=TQ�S�`Bg��<��+_�oX������N��逤>�,@FA�&��� �w��_�GI(A0���Z����K`�ϓ�3�IJbƬ ��$���ϔ�_� �O��B������;����E��i@����,��{�3�LAQ}� x3�4]�>ms�r���<8�/F�-�$��ۏ5����t�v#w��l�P�ak5��e�@'�=E�ȴ7��m���
�r�:]�x�6���Rk��[+�^k�'B�B���޴�|,VUŮ�҉�9��U��q�Okk�u��*��k��@)��8�7��R��@+/��?��˂1�(�Y�������l���	�@�O��H� �D�r�
f���� @-U��(i,/�%1j�9�ƄydJۢ��Ӄ�b�pE%�����6��e����tl$�ق8E�9衃=����޹O�ޗ�o�� �m�Ε�	B>����9��+�%��yI����{���W[�ʛ7��#�XM�v$>��-�0f�r$ 0M�[�/��� d#(�]�_Y1�)�p:������=D⟹��C��g�]"��J�V������OG��5OGľ���Wm�j� ����Y�OU�W�����b���Ԟ�m@DW�\�d�g<�&#Ze0x8�v���<��dN�Z�Ʀl(YdJZ"�!�Z1���c\fT�Yi���?������kQ*��+o���K�?���ݦ�^��Ɍj�AP|��jϯ8U�]�^���}�|6�W_{�����������o~J����xᒈ5��ƛҗ���3�d3Sjݠ% z�%��4�6#�ຑ���� �����b�E��3GkK��K����j����I+ͶԖ�����}z��C��ݥ������_Y^�׃;���N���W��mR�A����!f����Uyn��7��}* 	T;PIB�T��O�V@ $�aO��u�o�'kf=M��?\!jdf?Id��p}o�(�-�.����x��T9R� ��Ky>��	�~D�{G����%z���i�����G���ӵK�i���C��C�u�"���;����k$�95aG����D�f������ J%�{A�J����.64��H���uD�,�%0��J�$���N<lK�7�H��5q�a
a����#��&J-�=@�v�38_��s�" >����5
4�7�:8ReM���:�.��zu�"�cϹ�UȺ�D�eDM�r��@|F��U�o��?���.Jtp&=#�JiT���z�*���]Q�J���N��ਦ�'R�М�/>����'?��l�v(Vm����;���?�g�W�����A2(ø��d��|U���_�~��dC�(�V'�줨�"P��/�:�l���{H����H�F�.�1U�>1�&�e���c�,�g���F��<yz���՚&B+��t��b��*2�m���e�r���!P��RX��ў��=�~�<b�/�m�H�Ԏ +8���M;NC�� 0��Uy�$��"_�4x��wc>?�p�;��L�cu*"k#�,c�����Ц�x>F����D�����W^�����~�s��i�=
r9R*:���e^�I��*�^{w��5�[tΈ2`%�8��yУJy���e�@u�;J��5���� �|`�]��Ė� S���Wz߾v0Ca�7
�,�#�e@f1���`�|����'�Q����߃>�i�>��S�U��i�|o\��2O�<cG�t�eM�l��Rx��&d?��\�"^������n�^�
�`���k��R_���~�#����t��u�'�e�ֲ���&	��1��ڠw�v�^���y#@��xO� 	D��v\�X��`)$* B���R�m2�P$L���O�N+QA?��w�)m���dۍ:|�t �� ��R�!iރ��)P3f���~~`�4�r��L����*p�LS"U�g���~��<���۬g}Q�Ŭ	��3)'����7rh�zHp"?����t����Z{M�3�'�-�;Z�~���`O���5��H�>���1�)�co���]YZ����t����w?���x��_:/�$þ��=�Ml&���5��B�x3��x>Oq<O�V�(�/ͳPK5˃�'T�%�d#	�.=�0Z �*v`/z:2�k�&�yTIk��@�A�o�!��@�؞|��<H�a��@�a���7�I
�O�U~�sި�����/Y���ujR�Z�(� ժt����aZ'�QkP���?�W�NR�c܇�UK>�?p��vD��� �������v�nާ+��2��y���׾KG׏���c������}�>�a��F�v���X�:k��������3���|G�k��x�t�����<��-y^�QB�"���d"]@rZ�[��YF@tM�̛w5U(�f�L�Mߺ�:���p2��Ԑ��ʨO��j�SUnD+��a��'���1A�2�KgΊ��d<d�j&�-��IH$�Aw�
dlb}�>a࿈�L��fF/0�C^��e2N�%]W��-T�1k�Pxcq��}U����5�R�o���B�.ѨX���)K�g��*�Y�D��6��v���<�W�i��-mn�R�h<�ͭ-�x�=�������x@{�Gt�A���9ڸx��z�y�fP�hkC�3�����'�AZ��7�L�T�*`GĲ�L��h�k�i���'��	�����Q{����.��2�8{�,���k"DR�=��O�s������w�[(8��͊l�Z���JIqb�( Oi�sEjE�a�S���x��:�� Ǡ�����`3��������6�g����d7��fl٣	o�X V��'pݠ�� Jc'�Jj�I��L'Ȕ�T�WD�����������t�cs�����{��C��6��)m���v�y�ͤ�4R�ɿg�/�����V�0��Ϳ��R��t���;1 (����Kr�����S��E�����Ef\'(�.AK��0ಀV�m
"��
	��5�D��R$��!z��䚼�7t^��@�.�j��F[d�{���
�Zַ̎����ܢf"G%;>2���9g{�]��c�*G�T�@O5�����@�Cu0�M=�"U=�KW�:�tL�aL�R���ϓ�^g)7<��o��DZ_%��@AM�38>�$� D�<�|���؂�g��6, H>������b��o4&�������Y	dBJ2��O�9�\JRC�W.�יe9�}��C����n�K�S��3��xe84۫N��z͢�zW�+6v�Gx�:#�R�uJaM3�I$�W�X`L�MLa>�d^�t�y�E��l��6����{<�n:z}Z���Г�&��g��%R�Ш���QwZu�q~�^g�e���!�e��a���hb������ ~U�/).k2���H�ߡq6F]ӆ�xOj��A�\�@�/�0*s"}���E�T������Ӳ�g����7��i��o���62�n6Ȃʒp��Z�`�B��p�gBzڞ��>�'�e�-@m��8�~x�D��!ݻ}�ja����l[���
��oH���� � |�� QCއ�w�x(a8�?l�L"�:�e��VJ|�!��/ޗ��W�]��f��5�uj4j�K0����9��^��Y��T*%�	���$IU.�
��%ѪD{�0E�����lB���ب���{�xP�O��T��.�z93��a�Wh�Ҕ�7G��BT�:zz��j6��� �4���1�BL�<PܻRo�[]�
o�Pu��$�u��#޴y�`H��\(w��%Ze֩6�r��Dp�3�cgpf�"������]����Ktx�G��ɾH���*��6/Q	����<��m?�Z�R�2��-�Yd�J�*u���������>R'���gh�w��,�ٞ�3RK3���D�� �Q��B���"C��)@kI�K]���^]ڢ[������c�F
bT�$ �lf���j���cN5���}�;�[�E��Ν;t��U�\Y�c��JLhcYI�^���2�VK�&�N�u����ߐyc��r⻟�>`��`���ķ�� ͑żX�L��jQ��o��';Q#qZ�ׅj��ֻϋ�Ȑ�4$�H㚦ә8gK�6-��R�^��#ެ�'�ݽ{�ꭺdBj���~�th4�+Tc�����h����WW�yF����ؤ����"�1 =%ȉy�2o���5�>l�J�"����sh�>o�]���K0���d;a��r�h'Ѯ6�T��`���KN�d",�s�΄bo��6��%(צJ��9Rp�o�:� �)�1��x�n�^�0��@�ӊ!�I9�d7�d�^�$N�����{w��������Ml�`�:�LjR h11�+5�-ˆ� ���6��O?e 6��Dct����� �����t��ej�:C�6$�OBO-ɬLT2�V����G��8~<����4eP���k�i}y�:� �*�҅cM�f`�7��������/�l%NNy�s6��JD�VҞ!�H @az8����iP���čR�G���o���Z����ZҠ���3�BY-oȪ��}��x�"7.�͒D�Q�Tk���x/�$}���@k*����L�j�Tk�"�"��3��%"�hJ-�N/�t�"�;{V�ήu�.Oi��Cď�v��&E�G�(m�N(� �WPR��MM��ZuJ�� ��4�\u���ؕ���d��Z�3
���7�ΫD�^+ ��X�*)�yv^���y���y0I��>�-c"�s(�IDypHپr�9YS0��Pe_앃�<�_��k�)fjj�����4�A�m�,0�IǨ2jdK�V��h��c{�"g�W���Bk���C��ߣ��L=F~I�N$5��®�}#�`����  ��IDAT������^��^Y٠�v���O�~u I(W��!�aʑ֩�^I�X�^��e4���pNB���������t�Rօ��$�D�%(�AI���P���[Z�0�YW��yb�*���?��Y'e��%�3�!U0�a�6}&2*�]���� ��S���/r9kR'Q�8!���i�9��g���}����I� ps�]޼�?�JV�;eQ���RV6J-��^ X����"sXjWh�~�]�֢��nH�����E���k/S�U�1���UfPO��t&<eL���(PF���4f'(E��F_�����t3�Y�taI��U tI8f�<&c�^[x(ŗW��7�]�2���&�ܢ�N�	N3Z*�S�Q|�AZ�Q����:q�S��a�&��@�Z�j\��z�JKT6�����M�[�2D���k4�R���vK�}�xsyC"=��4a�Њ�t?�X7�0Ȟ���Ԑ���n~�)���~!��H�(���駟I��W^{�V�6�U����V�q��Vv4����#��ۥ��g����6��cZ]_�o|�]�?����:{�";�$�͈�Oو��A�ֱ��A�05Wٲ��N�yl�%�9�Ss��tNO�?����G��6�ʥK�� ��)iV�M�AC]"T�V;�<�k��ߛ� ����`��w��^588��6��r�`�\� 2m�Z���E��,���MU��Ʒ	m��	; )�������Fo�atU�7���������=�쉀F�l%պM����F�M�Dd���R�<ݥ6xg����5�56��ls�!�s���d��M�ܬQ�g[d�mߣ���gt��=���u�f0��?�� �$����a.��AI����I�=�i R�E���:K�Kb��܅����[g�6��+{�<?�v��zـ7k��Df��Z�
J���$-�I%x����S��H��߰�K5E��P��G����_��F65�{W�ze8�v^*Ӕ�EGИ�O~�������� !����^�Ƒ-E��jg��P�i�Ǆ:pjN7T�q�q�bi!�$�R�n�m՜�ϟ��/�͎Ԓ"�,!���ӏh @>}��$��q�T�:T� �b�����^������˗$�;���L(�un�>�I.8���Jwc}�wPq�@�7T�a�s��4K��O���Җ�"�d>2��x�n`�-��ˊ
Q�Î���h6`nUz�E����RSs����'/���l�ޓ]��y��T�"NEEU���X�����jq�f�T��A��ҙ�}����ٽ=������"�<o�9����NRB0��1��UyM�RTyI2�;P������=����>�R��PAl6�i<d+Ş,8R.�x����S,j��.
<�+���(��<�f�Xy:/;���ͯ孁9O��́p�����k��x���P'k�Vu����9��g���o�f��W��e�s6���s&�A�^��1�w��3C%�P����b��HB�L�E���*�|2j�m���� ��C:�t@��A �ӱ *�(�r�n�9J��K�2�5��֕��r�\F����J	pH�A��$Kn�6~�{�^�ޠ
�$� ����7���;2L^�E|~��N����g�=d�Kڌ�Ou�)� ��Dt��[WdA���].�BOa�#{XP�|�%��&[a��U��-&��[�U/��/5>�b' �Q<�6���ҭ�oQ�+ɖ-�[�]�&��vuY3�`� �a/�ZD������e�P��&Z��������Q���u�r������G�U��W��u!�jx6�ؓ�dܳg�B�Q��l�i$�CXH�e�Cl��jY�}����mȉ#��f��ed�X{�d�E��o~>�n��@��Z�?iV4�������sA�_j�EV��R�͋�Ov��\�E4:�ŹB�o��B���h�Q��/)��^��K�t�;�Q�@�C�֙���\D���Z;O���E �*���ر���g��v�Vؘ�b,ࡕ�G�D+�h@
��Ͻ��F�ZSDD@�
N��*Ol��YY���}�ώ֌�fE�~JB��KfP�ĸδ��Ԋ�]�,�vPPDFu_R/��xtt@�1��\���}q��x �Q)2�Uv�5���1�X���t��Z�8G�ÿ�Z*P?��#z��C��6�ڴ��J��]͒����������^Y�>ij 1�
��]m��4�� �4R����l���bk��z����x���ޏ�KZ@���_�-�N!2���K�4����Gs�6����&<?�P���ñ�6�q�%�{D�Ǉ4�o�
`�BB6�G��������]j�Ml ��wޠك����Ќ�����
�!����a������:]~�*;�3[[r�x�X0���R4&�jI�u�9i���u�s�#w��j(B(h� 
�4�FM�pzB��D*q�=tF%���^mkt��9u��JЂPC7N����S�6P���/��	%��j�X	W�W#㊉5D���%�iM �� M���I�������"
2]��{$�Bc~H.I�
P-B�T�I��iw mh8�c��P����3��ڵ�~�8?�VQ�F��T�9����}�VS��_��JH��>�x��j�h쑌/��%Q�tVKJ%NCk���V<��i;�L,)
���M�c�ɞ!k���:��T�y���4��dR���������͚�M��}L����Aթ�ʃ� � >w�PU-z��
9	�9�"0�,��1z�i�Fa.K ��W_}���g4��+��R�)��b���1�:@��@�ם۷h��a�xH>�K��;�#�;���}y�3�q#��l�\VC���;��EQ��[�⅛���1Q���Dx,dD=@}
C��o�,�A,qt]�+e����^�����ň�Sv_����^`֢�	e�x��=?��?Y�[�(ju�b��I3�b��y����e���(ì�(���@�KS����ߤ����y`>o A �1�Q
���`̆º(����7�P�PR�9�IG��cG�]j�O�^��:��Ж&��p��}*��B��im}�v�蚫����g"�p�^z�FjK}�/���%��g��`6lޟ���H��Km6�K�>k�Kֆ)�=�߄�R���$0̞W��e,�z����H�!g�v�=J�>���ޤ�î\��s�����h}e�mtC�Q��IҖ[v���$���t4]�&���r��t�i�{i����[��T��Onj�/^�`>\$�Hf����=_nǊϿ؇��"Q���G6��d7d��3��H(f���ء�� ���e��J�`���7[~�E�.;���<���Lh�89(�m��o��e*��������v�#�h���
C�����#��A�Ā�!`������_�H/]�Hw�4N'��q9S�R��H}4�����+��$���ϞK�VWV%+)Ž��#����|uY�OL��w��fAt����;��pJ>���-�v�D��I��@�(AV�ݪ�E�[�]��������Vi�n�6�L	�_��gs�V�U��@�b���d�҄����ٸ!�2��""m86�u
G]N���Q�G��}��n��Jпjͪ�L�	-�.�6�ڨ�YD1
��Ht��7E"Z8��F�(Z$�:���ԟ,8Yį��HJ&��[�P8-"L�7��� (\�MmB;�&���,�u�2���@��H��Ԗ�UH�5q�M��e?�D������߽� `L��}��/ySb08aG��֬/�wP��b�8�ڣG7�Z�X���Uz�͠�{��&�F�DI���W�lty�4ªPѯo4ѥ���%�P��L@���߁����!�8h��C�,/ӭ;����*m��H���p@�V�X	����g'<(�����ԛB�3嵋(���uC�Bu�P�[���N�XL��:M{]�O��2�j���|�u��)"�5�OPl�<n!2C6Afs��q����S��[��`�"O1��ݽ=Zf�{�7%�l�����9j ��6���V�� >6(+P�EOι
�@�t��.�tT�}ggJ >0�(1�@N�|.�V8q2��3(�q���M���C�+�
�>�+Y� �NNc����2?�3���x@�	���w�J6ϫ�;���}�����׆�H�Z��L��
2��RFY�Qm<l��zE�d�����uY���"w�k�ԕ�-v�	{u<׶p�sPH�B�=5G��P�X�PD]�{�s3��)Dy��M�mj�<?�"��u�����t��eQL��P�NҮ�=��1ĳ�d�5`�|������Q�Z��r�EIv8�P��D�L���~���0�E���eIC�B��\6��_�K�pl��>�DK�峣�1,f1�Ή���RfZ���	���g��'��rd�{�Jd1P�]�O��d�UF�ԕGY�0xF��3���
J�A��@6@!�R�K�gp@B�S��a�Fj� ��V�Q��Pa��*�bV��;�8&!P��
����������n˱q2���S��&����`��3��>JUzl��Q� ���;��'����\,�;y1��-�M�kBI� t��yC���'����&�h�lݖÅ�s�* �i��/Q]Gݺ ���p�����#���m::8�Ҧ�[�ի7hsy�*�:�*�	YI��֬�����G�q�m2@6@�}'1_��k �b�)5�M��ܢ�n}���Q{�%�&�S�m��M��)�ڐ<C��1߰�=E�ZfF����P�-��A!:�ۗņ��s����I3^z.sz堓�'[��b	�в��r^X̅E� 
�>�V���b%M����A����/�ӌ���dFvH�,Z��i�D<� ����jLOD�wL��dL�L�&א�g�	=i�(cF�T�����{/ݠ|�{t<���%�v�����	��X������Z!�@���yC�Uz�Cc�3Ġxg�	�#vH�Ѣ�
]�X�=�Ƅ�{�P����st��z4>�����'wU#d���d�ϒ�6�lF	��:�&�9��@ԝt���#�U���&��9���\�]��J��q, ��)Q͌ޜ^�vEj�-����:��F���@�bť���(��°`�rQ#o�2�T�^>ӝ7b��QX�E2��c�v�T��� T1\6Dd\�"���DK���1��Q�s�s)�q3@(:����H�y���줊l&E��G&�k�i ��s tmdk���hC�Z@�O�	�=��G���})'����m�v�79�}��v���P��݃}��18ښ��<�pn"(3�쌅�6fǶ?ѐ��e����#��.�Iy�J#6� ���j�,�#>�i��m��󏥇���C	fŖ��p��� m�=O<˒5�Wi'��[�}����o�!��6���a'���w�O~����l�Wj-����28-Qo<̔�Q/[�qI&�4�wD���A}d�𼣒(n�6�sy^Ȯc|A�m������;�����ң3����D���_���%�z��G��W�	Ts0?�Û�ؔ�Vw:x�ё�t��Y�r��8e�u����m��2�2�~�����K���������J��͂�G��_���xAhs9�����C8XI���_�,��&�꘥���x�7��(Ǿ��HJ
މ�w�%�+��b�प�Ve��[�X�#�4ŶǶ���r���px�/)٦P�>��f��E���V����fҏ�� �{�iO$(�[CMa����;
ء�7I�R�s�G�|�}���M�&R�椈�u>�5J�/�yS�z��`�:�QX�|.�����PmVg���l��j	5Ӕ�?���A�x�n�<;^��
�"A�{vW�->=oNu}>����?�Wv��ɗ]R���6�i�'��ic�9��B�Tu|�\F
A�Th�e
MXH��e�/�z5_ʮ����4PTU�D{����5�D�i>_�?8��'���2|I����ױ��sa�%�`������R�KEEb��S_a`T%�`#�/,���+6�ϝ�`�#kw��!؄G���cm�UDlz�GF���_)�����k1�.[J���-�&v�Jd�@���ڶV:E*hBZJ�khv�vA�h���P�s�2Z��|&�zkI
Hf���%����򾣣#��>�R�M�\������0f$�UdL#�L�V${��#�����K�nÙp��Ao(����Hm`E|�a0�E�MJi�.���~�}����������Z#�o�fU����� 0������(Cl������#�����"WU���\����T�f&t��b1��Z��Zb�Û��NY�24D�GsE�|�*C���6�Y���c/`P~�Nԇ��+%��mq!����oM��h���@2u���xC��M~H#Լ��eDB����I�Ѵ��dQ����ҋ������e��	]<{N��R���>�s�>߾-���ަ�q�>޾C��XjLDJ?R~6|4u����Ue�׊�|��W<���Z���N�7����;h��.�P�,�K��D��3͵/OR+�:S��S��CC���	�z<��6���F�;"Wm��<�e����R)Τ�5�;�����{����N�T�<����D��,F��6[�P��CD��Y/�H6_ݕ�zBůR�g,���"/�@a&�d옰��+(�^��B� E;��-И�q�}��.kU�sG0���^��0���f�4�����e%�̧R���������q�5C8�$�%}9a$C��
�^��星�1?�~ȆtP9�=�V��q�����o�k��g~H�T�'P��ߠ8�D�;���L
�.���vHoB�������/�q
��~� �"�O�;ӡ�A܍k��?����&��;���G��]��/߿CW�^���_�o&_��7�-���H樴l@�%�G�21��J���C�nKP &���f�J������V��� ��+W����ݻ�h��h��¯-/Kdsww��~zS@ �ya���f�0�j;�&���]������]�G�&I\�qo���-P yL���GMɤ"�	9n�4���B��p�֣:)Y�5uo�x��{l]Y��y��VV���!�Rgp����eY߳�����ٯ������bd�����G�$ Z��/6GǇ���$������fSUH�s�{���H����XhQTkV�&%��k�O��J�GT����A���A���C:�j�СJ���K�>R�k_��SZ<ӹ�>������O;wn�卶�Gᙈ��(w{a�B�����}8)��J�O9�� ��";�e	E�	�Fh՞��`PVme���F�����	�����~��y���{�����Y ��9
�@!��EbO��f��ڤ��(�H�]X-PI�k�$"֢���;�k�%)�I${����ȘA��e�!���}�~�_�U���R@`���hH{�ވ��i�}I� �"C�~�x�U���8�{�� �����?�����Z >�V��w�1��;M�'C�:i�Q�:|P��r�2ds�	�c�;��C�f�qL�.n�> �I�22g>D��2+Qq����I#�
���ǧ"��l<�a2� 4_�$B<p�y�q&��P ���YѶ��$�CXD��bYb��W��%��U�+P���ڬ,��������w��R����:����}�#���b�� ,4	�?{�:"��J���M��3�Ł�T��_Pk�`Y!�����B(q��{]���ݺy�������ݛY�^�a'����{�} I��"�єRء9��_a��A����';�OfȢAɒAsI��@�`�魺�k��/���}���y��� $���ꪺ�7���?�����wXB�h�%�a%Chde�U�p�,��T��j�;q�AT���O�2u��?99%qY��4���)�JCH[J��ّ�^-zP?%�_�E����ŒaS�o5������ʼ�aAy�F�/��SYv�(Ǿ�KK߸�t%�	�Ud��khl}<�(͌gFIKt�tt2�@e����C���b�h�LA�@흯����z�@Q��",W��
��rt�\＝��M-r��J��,�N�H'ە�W����~�T�����8�D��{m�v��+Н%����Y%(S���4PR��N�bX��Ɂ��H�����&�BN�3f?��N�"u���)��Ϲæ���#�@�t�Nf�� �Vl��m�r��$�V���e�wQM�-���9~V��}TN���Gξ�׈Q�b�l.l�K��jM��ܩ�k��kF��0�	�$�9�v��
��q�>�W t��
��%����a�����.�Ϩ�S�rF�6�fn�ش��,7DJ�\��}��m:>]g
��ֽ���ѢA��ؒj�����\�ȩ[d�!��-���VK!��nf'��b�`!@�95�ذ���3�)3�F������cy���ڢ���,"R�_����_���������7�o}�;d8 ³D=�x!;��\^ې�ޚ��F� jG�� 
��(xk�|8��k�56g^!��ˣ���O7�E��1���p�x�5��	��b�]�VA�1.6>���E��"Å�߼~]�cF��`u���jm�'�k�(D*����z>&ݩ�>L��VΩ�iʸ�G�˾�5VJW�rc�����%�?�B-Tcf��G�)���dxX�g�&�9�����N��t��i�U;���\�=�K�m���|�2�m6S�O�}��T��ߤ�Y�o6g��E��=#&HA,�	���h���ޏ��|"��X6њh�O�ht���BJT�~����nGp}#[|��jt��$��uz?��-s�xL:�^��*��q����)d���jBoL�*aA?��v�W@`�V�>�a(*}2��#��PP^�KE5�W*�[����Op|�?�q��!I��p�A������gL��
��6�H n�)���hu�9;� ԗ�V|�j}u��Q��PmH���B6PB���@���U
�v�e1<��`��>/ ����a+�ɂ|�y1�R6� A8�*��`��/�L�� =�.�u�:�Nx��5��Ԗ��HF���:����y`�A��T���h�.��i�k�i�c���AӠp�<1f!VQ�3jT�`�C@�\���%�Ђ}�b��H4; ��}�.�`-3)��՞�?p����xc��> �D�p����!�/]���m�{j��yK%J�<`��P�����6�;p1(g¼�fA�L�_#�g�X��c�>�G���LdK���x����#�2�'�>��>Cd�{�LB0Ϟ�E��β�Χ����	�,�Ǒ�v��xm�g�o4W��88>fCpD�&�VU�y��P�E�����ٗp��TV��'Pn�K��(L2�O=>���ʏ��D�4�|���T,]��=b=jXu
 �м��pl�mD�6[@Q�/����A7�rJԋ�B|a0I�@��(�~FW��M�@�ޑ�>#�\�.��4~}�y�/w9	ӸEG`�ZZ�:�[;۔!/ԩ�l�5_����L��!k� X��mm�3#����.ΙN�;]�o't��G��|�ZF���"]�F�r�VO!�z@58=4n^�r��:2c{ft`��bl�Q�	��qV�ᴎ������P���bͳso"�x6&<O���U�"����~�T�'�����`���g3C�����E����φ���K����եr����s�I}	@16�H������Qu�ᵿ(����~f�z�a�r��C���x:�Hz;-���r��3��]ft�ha�?���E?5Џ��_���o��7n�f�G ���)�n?G�P� AkE���CR�[����]���l_�,���<�lv���[�8e~ t�6���������������RR�.w���o�[
�����u����������(r����ƺ���_���~FZ��T1��1ޠG/�f:���
0��Z�u�ܼy��R_��w@�V��H��!��"O�}f�F 2��b�YYf���c�ۖ�9R��V �o��&��#y����?��/��	N���n�̭u3ۉ�7�,:���n'��-��f�3P��;���;�F��L��2A�2
�~TA�상O�Ov���}F[�SE�#�F�1p�z�p��$V1�g:�� �!��蟋�-*�*Q o��a��_ ��_���?$� �� ޜ����KSO]�c̒tּm��+�֧F	�����^ۖΓf+��/� pEV!Mt���j�Ǐ�=����_�v���5~�����"*��Ա�|1�iF�<���9�(�JD����Pb-KW�7?���6��l�\Yf�aM��
 �L�������7�����,t�Vs�~�AhG��(<k� ~�2��ü)U\�J=:�����V�c��q�3��ږ��P�IOmӍ�K��{_����븁�aP�'@�3ݿu�+S�=S<-��3P�Gಠ�sB*h� ����������w�e�s��UG��>���4@��2d�jp�'g�j�.�c����=
�h5��5wB�>wz��K���q�ڿ��G��a��ca^�f��ى1x�5F��߰�2[�ս+[��Y��NQ�p]E�9��˯v>p�����B�m��C���Z�+W7/˕�˲�{=��ؤ2���P���4>0��h�lA���,//�a����O|4�������h��u�]���y?cr�hx(��ܑ�-dL�?Ɍ}h�ָ|&��Di恩r����d��58��1�� ;��<�Èh�����6C��(7�*J�����֗��|���H�
J��0P� ��M�K�;B@����2�.(8 94J]NR+��/�>�X�h��^��7�4[���| ����s\��d��#/l\��_|E��qS��d��)�Y]z��̈́�ʊ��<�罕Z����Y[Z�������)�0Lv�7��hp��9SG�f�d�����>:(�kD6/��5��^~�M�1�  �S����4`��1����Ha�Zt|bW�5V)�D��.i�[C4��S�4��S�Å�p��ܯ~�xD=�o�e��b�ȝ�4l֤�R�k�ǄK����|C��<2�lG�=5�i�<�@+���0�3r	�-3��c��@53�!{������/P�׺}9���Y��)�j"z���̬��l���j����vgNh���G�	D� P�Ⱦɍ��C��V�$�*�����{om�E�֜@�|�*s�m�F�q��{�5ֺ
��nʃ����_��'�����۷9���ܼqE�ɜ5��!rMm�-R�_|N�k(o�����C=
U�(�Up�"��F�Hn��[MZ���{cd�����=i������^��en}� ���;i�X��/�X�n�5SGmZx@��Ц�>ȶS�M�tx�����lo��xr@�V��5O
/Z=`��	'VR�w\\�w����,���Z(�*L�?C�����ߢm�9�ɴ GpR���E.Xߞ�����qQdaNZ<�{��>YZ��6|�Bl�r�T�Ei�����5��>�9�׮�ˊ���?��[��z2R����'�} ��X/�E��1P�y�%�4u<u"Ie*,
����{N�~��?NFV�Ro�U��[�?d�.�{O;.��}��8DmAM6��(.ڋ������o�<mɠ�Q�ٿ磻c뼜!E@VT��),(!��Q\	\V��OrD�X[��ʒG.�sôzwqP҈�r��
|۟�#�e��g���-�aj�
ބg��"/V迏�ց�>��E�������QŪ���iv�6@�}l��0�Q�k��>��5�[��c�T�q�w,�ӑ��S+�{#��P��j���`}<��l�֢?F�Vb,4+��������Y��σ�	�P��h���FC�[�^�p��R�y�7�X@ {�x����P6�U7����2��g����w��`w����GB/���L�"��t����^���ʶp��R)-���
���ˣ�{q}熬��
�;,��g�$��*2�U�'�Y�	4/��O�i����a���3�N�
%t��f�i�ۛr�Ҷ�dA=�۔��L�N���r�ś����:��x)R��Y��U*�V��P ���#����2�97�K
vQ�(B^یV�!��r��j�������ٌ���L��2��܏�g.��U�^�8�7T/!?�E�zK�&��%Q�|��U:�x�be��C��J�8��|!�<+X�Ț¢���d��Al��)A���5���_��=#77/Qmi�u޾��ro���;>��n&�n��6�-&2a�,gO2PNQ�:6��\nmmqr��"�����)u~`Rب{i�6�.n�l�w�!#��G����R��&:�"�lI0�IwX�D��_}��䙍K��C���ƚ��Q5ի�5����k^6R˄ ��L�EF(O�n
&�ܘ�Ϸ�|�(��a� �� Zn���iB?L��	�S��gh�"^�U��ϫ�a"}�'S<&7�����&�@1��5��9�h2k����(���2��ϐ�E_�����6�ȎF�\ui�ܙR!�F�i�o�����xD�uj�"[:^�L��%�Lkd8��������go���eC6~Y�5ѿQ���H������P)����?������("��Ì�0jnº��t"2�`oE<�skaƺO�<��a�f�	[Y$dE7�(���[��/~�g��_�ݓ#��?�#���9i�yjTl��#��h��}���h*�g{�V�N�,���[=7�G�{o^�Խ�`[PUA[�B�n����Y���?���|�����˜�-�wޡ��?���� 04-�>b1V �R ���'��n��݇<C���#��VY�F�2�9��0�����f[� ��ǒeFe��^�0��c�q�YY�2o*PCYú~v�5�e�Q�� ��y%&b�c/��� ������Cu��(�a3`,C�M���h����=f�o߾��>�=�Gz>@��\�����
=2�Y҄@�GK�ʼ�\ӽV�
��ˌ�sq�KG0�\ �צ��(
ĉ���l�PH	�L	�-�nݒ��>E�X�Pԥ2��1|����uX5F.U�u{���|Sf�<��{[����ɼ��e�VY���E\�4KX(#�ꅿ����9��FUʠُp%dUPs6'�K���< l��ӝZ;�3���B��T�<Z�T�j�� 	�����'��� ��ӄ���y}ix�U{rq�2��(�D�b:��}�aP�E���ݑ�xB��)�C�Pm�ړq&��X��X�"����`�`v$(�ɩ@��lO� F�W�a�G�@�(ج�u�݀zb�@
Oef�M�Ps
�$�9En�{�xe/�cd�(7�R����:�]b�-7�<@q`K��E���G�V�����Ѻ'mZ�0��(o0:y��6*��9������f��[�
���5��.ɕ�+�I�5��8�ou��΁���-qS=�P�i��g'�6��uZ`L��`fg�'*n��u�mӾ#y�ӱx����X�V7���u۵뗘S.d�C�EXC�HmL
u�NW,�W0� �*�#����n�]K7D(�t��D�)�Y!O;2O!_l\�a��!%t@: �.z����(�����9%�[tB����f��T>�B(������4rsc��y: ��:�\9���DϠ��t���3�F�p8�0�=�r�'�������<�yYn\��l#d�߽����{W�=ٓ��T\<md2n��N%Qu8Ƀѱtf5RTu���Ց=�{D����{dC���s��鹫{�T7�8�IҖ�z��z���#u��@����(vo쉅L�~��+;��o�"פ'/]�I��l+
���k���tj�TBd?�U 
�d�U�T�\G���s��D�2\&�l�?�#wV+Zf�����j�:��������ưI���@ڮ��Չ+�(>���wQ�_[	\?�M[���r� ��]o����99V��Į `�0';i �F�NP�PL��l]�!�"���0~8:���{r��LN2�Be\k�v�,l �;��ݹwW���-���3@2O���r�t~�V̹D! ]o]�S/����mnȯ��/�7�~S�y�PA١4{�RLF���7������#�$F��/A�A6f{cCn+؜�뮯�p6Q��!C@���|��~���ү�m��gG'�G��'�y��P �q���Ĥ`g��:C������A��2>;�0�Q����kT�
 ��l͘����5y����g_�S���%`Avp:��׾�5n|_�җ._���d��A#F��p�°)f
�f�i�k=�G���@ǯ� E�� �q���
X����EVS��}Rs��d}r��r��܄�P�=F*���3�N��_$iԵ�I��i����-���zĵ����X��,��}����M:i�t��ظQ�C��\�Kcl@)��th[]�ƷG����5�( x1Sۜ%t��o��D�~CӔm���6%v�V������zhI��P@��gg{K�}F�!p�NW�S+v��Q���<�lN�V�b/�	��=�m�,�fv�u:��soy�D%�b���]���&2�͠����:F��ŵ"ĢlK�I��`���"%V��e��{�IȦ�U_|���@ć�=�V��!��[ ��xMPf@� �*��{�NV�h}x�U�0��U��G�\p������ˊ� 4C���gj�Qg�׍?[��}!�;��F3�_�5�Cז�9��
����a�2�K���e6��x�Z>_x��2m`1����#�ް�#�uA��M�f���&L+e0t�2 ���|��N��ϊZ���S�,��֘>1�wQ�T||��/ܦ���`�eHi�g��rK!��`eL)� jz�X;�q��|d�B�0��'3�a�yj@����P�{+�y����zk8ֹХO��{� �*��ǡ�BftP����M���p`m�"k��^��ݕi1���+�g��o,�^��E<�_?�aBd�Q�MA/��(t,X�;�e),K�ToV�a�M��"��ߖ)�]*�|��`ˈMj�A�)o��,�N{���hqI?��<��5U�+�ތ�*d��1�񠱘P�;5C���LQJ�w9R� �ǵ��D;^9��e�(>��M��$.E>�ЯF'�>��e3nHs����SyS�����ɩ<Z�d`�7JԹ��m1B��{_��\�[r|�/u���.�9�ո�o8@q6*͒M�M�a�V�����Y����B�˂5��X�Jù���e:��@_->��k�=��D,�\��A��u�9��-����z��);-�Q1*��|,�e�0�;ڠ���E��	����qk����s����#UJ*#�#��F ����9�N��O�L~k9�>[P��+���,��\�wr6��(�����ѲA���:�ۗ(�	
3��A��x*r��+�''�7ߐ�v�T�3Ԇ�3��T��l9��B���j�y�=b���X���ynO�@_j��� ͙?���Q8���Z�Ny|t 
f�g��!��F�tDU�Ȩ��8�e���`��fڅZ�n�^�)?����Ͻ�ڨ��ǒtZ2R�A�d0��ߐ_��_�W�=C岿��W����`�
*|�2���8 4���!�0'���3�$A�����3#g�jC�cI��H��?8�7gX7A�H]�c�
7E5��9l>��d�BI;�L��c�"EU����:���Su*������ ���/E�Of������Z<s^B�l� ex�eE�kntQ��BX[@�櫟v"6�f�H��f��:>ΖS��:V'Ǽ֝�Kw����:\�&�+dY���Wf%�ӪC@��Z��%E�#�G�M"c �����z�5���:����:���� �Y�SٸZ�@�Wk���v�3�7�b�d�"�Td�?9���c�"i��K)�*@gm(B6���%9W�ss,% Aq5A��Q���9�܁�?QT�re�y�rl��]��AZ4��賚Yp<�y@
}�$�6BF�$}4>n\���������>���9�G��S{نUf��:����?(+&W�7bzilc��G�v"��/�9�N|���D�j��U%Q�K�,����-d	k�R	[��|/������-�'bmFI�>��FhI��@���6hM�OG�	AS�l+��Tm��(k¹����u�:��e#!2�ч5�����
�2�aP�*�~�|Vjkϲt�k��R-��W���	@YB�(��}�3����#���{b�ĢUv�,�,������,�EUl#�7��~��D�M�a�I�w���-0�|<��i7�Ò=::d}fث�^J�6]���b��3��ڔg��I ?�~�7�6}k}�J�����v�hp���!��c^sW�\1��1�eE� �J<.�YI��p��6Y�&���`ѩ<�%���8��klᒞQ�}�����v$+��Am��Ϭ��Oi�}��w�P=rjh�Qs8	{��3��{���/m]�IuO�i���#�;[���?>�{��i-6�ZY7��L-c��E(1�(12��Wp�t<@�;���}�t�v`x�)3L�$�DN's���r�՗T�t�����C���N�lf��Jo�#�~GNOX��j��ڲ���(2y�\x�Q;U�Ӡ�r���(��k8��t��T��!A�T���	���:>X�P_������1�1rk��!d��H�l����dnHٖ��P#v���,N>����
բM�W�lY������~���ء�7�M�u�EfTF����މ��c��͘�ٯ	٭���=w"��̛z�83 	�ǂ�sf�Ii�54�賁|
�� I��o�{�j�������c���������s���ޒ���A���t@�	����h��`���� �h0d������}V��I��5������������'b5���@a�5�u����#d�Ԙ���<>�'*���!(9Gd����\�ڑ���_��믭��g��[
�u�R�?����d�I|�W�W~���+7e���o~K��ﰎ`0�������G4�B)��t}P];�?�+�?�i�,>?�Ղj�d�/X�6_`���E�_�㚮�_��@Ѩ�|�ۤ�,&�]��OO�*f:1��,C�katq�]X�{7��{oΆ��lmo��xA;�X�ȱOa�O��S�fa��yQ���}��>����U��\w � _
J�(��: ����9E(���l��}F4������� �
�(nĜ�d������"G͎)��ё2��(2�`�p����Ӫ�Q¦k˺��N=�؋��=ؕ�o+X��t���lPȘA	Y&�;��S�M��������P_�[WxQ�,#��,a�����i����˥J�!��0g�M�"�ߑ�� Nɖ�����9��П��h���:w�V��<h�"��q�J����]]���5�6�)�[B �� �G�5�	fy����(�̳Otn�,��C��)q�6kxFP$��(B4��1�JC\%�˶9Oh�skE�C���Jlp�lϓ��/L��F�s�wt�d	���(�1���Ļ�>�7�;�][��u�#ؖyP�� V�0�(�MCb�奟�}e�6��>�(ŀ]������p��]R|/��z�X�]���^��![�7m�Ĭ]d��Ƕ`��g�s�{ແ~&�h��9���A�e�<���(	*˱���f���U�n��'�w�@ad������~��w�H�ӗ�C��d�`1���XH�P�݃�E;v�0g`��꓃�	R��U{}:8�GЕ�H��>�gß}�ֳ<���{�!����9m�m�%�6���D��%�eZq}�^z�?�T����4L�(Jt^��GQ=�z��|�"�## �N-x��L�����-cQ����̟J	(��k�h?+��A�;�j)�PT�¯�Qp�-�]_S)�#4O-�������Q�	�Eߘ!�+��w��k���y�hO��
����HÅlmj�!��{�+B��������ߗ�޸-��~Q����+�=�~�Yy��PN��H7���}_�����a>e�xQ(�T����8�P���-����"s�_[��$k=�Kd�,�m��t��@�mEw	����g��D��#a�Y�ٻ��$L��=�� ֯�F${
f���f��f��|C��
���&&l�Wa֬�)rw�R+BƓj@LMN`��!��.������N�|Z��͜jQFGR�K���Jg�0�D��C�ʾ�U`y�ִ�r�l���V�?�Bp|�z6)'dx41�E��6�������t"���1��. ��������=�z�k~�CM�9��ho_��Dv�W�*�,���h�H*�N0���j���}� �s�!���&���a��T�����/��_�W����fooO����}�v�\�~]������ܐ��C��p>���$�K{�+��]��4�)3�V׆͚j� <��W�&�����߸|�& c��wx _��7�{o}_�������������ߒK�w��x��}�H�3����XL8�!��@0=KO�Oe��!�T�/]�\�(~����%Z B���\�	�᠘�������l���[��_#}}��G�m� �]��
�͖���3�9�ǝ�l��<>;S�����6:K�E�����i!��X�M�s����G�3�X�1*�>�EA"U}���\S ��	�0l_��:����l�Q��`O���b��Ru�0?1�&���h��t���᱌h�̛<l��rOk���F�3ʔ�,�:P
�(��Ȼ���4��8W}
;:�����f�B'�Ꙡ�Tz��ی������q����ێH�$?I���1��K���`^=�Х�S�T{D�$��8�z`ص�^�)P�Tԏ��"� ^��lv-3�	f�ĩ��5�%�͎�^�w�r!�k�I9�s�X?Ŵ�ЊC� k��t��^ C�� 5�����`�)r�W��ۨ�!+o5�^%%c��_@��lP��-W��]�)��h������)L=��8��MoDK��ӓ�nKzs��[0�E0�^���t��&��Y�Z4��KA����K�|��_�{�=�� �e�BM6���N���g6^��X���n5i�?�}��<�w���Q1�'	J��ȝ�l��Rq^����A�������,����*Y)�ll���2�J���t��U���5�� _��Q%������W��� q9D��A`U��fE[L}�
����=���q���Z�&�Â�<�V ;c_z�E������B<H�8`}4r�����[��'�v�h�ZEMb�9�<0�"��H��Ԯ����g�֊g�ʄ�\�!�h�k��JA�=��AF��l�#3gqs~ 4S��Uf0dLcKݯ
^�5�E���D��b����w'ǲ��`(���Q�o�Җ,�����W��wO�Nd��D\8A�_Ɩ5���""�
����q��ڻoʵ�-���3t8�������X��zC�>~$��X�|�!�V9^P�@ӱ]@6�[
��bK{O�Q��#p��E�l[��͎��ƍ�K\�!3PF⼨8�4)��[��#��pOn�=Wd#����Ȧ�~Ǣ�B�s
y�>S�w��V���R��s���ҋR�w����o��lJ~nA=�Tu�p:�Ǒ;Λl�sw:c��n��Z�J �E�Z��!�@�T��iH��Q_�t�x�P�����.M^^�0;��f�������/e�͇�\����>zU ��g:�R��ח���������95��р-"���&ʒ�z��	zԷ��]ifjX�)��B�!��FO� ƆY4�s��g��?c��K������%�ss�R��B�n��K�벵֓��1��^K:��u�x�X`�9.�(-E�M��&l��63Ȅ�Ư��p6�7������Q:�:^���/��";�2Y���o}W��w�N *݆�(0�Z�|�c���PK}נ׍zPHM�$��9x�@7�y�Rm3����i�6�s@�dO�Q�S�T����2�/A}���n�m�j�Y/q=:fsup�H�t�>R[1�8=�~��l*8����p�v�N���LH�`��V�~-Mn<	ِ�TQه3�����c��`��AU���ޡ㈱��Y#Y�[�lǕsO�&҆��J�2�XXN�[b�Y�esQ
�r+jr�X��(�u�:h�&���I�suG�?kV�TY�8�Ck��/�N�dc�K���
��+��-v���A=
��Tg�?�C���^B��ׅ&^��K���'	���s���5d:`�8��L�vy&��RU2�����iJ�ҏt�����-�X��<�w]��aT_�H��hbZ�2sDr�#ã*���3UF�v��ym�������_~����ρ���R9krs�0y{� F&*��K��iZ{z!� !]�8�*	~m��Ư7Nmސ�!�a>88����RhASp�P6�)���|��7��P���6p�ݐ���N`��Tm��d\�����5��F����lhD���sf�eحQ��`��6��"F��}��\�]��2��d�co /ѽ�I�wQ�0b���STxF��.�'����i��#�f4x���LMT~_��Veg��Bv�������	2�` hAn�������1Y�kϘ������v��_12��韄6����)og��}�nmn�k��&�����
q�Δ�Y���X[�;.�n\���� L��f�5FS��>����ِ�>�8Z��U}��'��p�~�2>��p�UE�=�YW{�0E>�a
B��cٜ��
6��Xa��r�<ڻJ�������y����ޓ�:�͍���ى��my��{�?ɸaj�s�0R��GB��~���Q��x?;��N%U�y睾�v�9y��-���%?��k�w��EyQ���o���=�$F�%����3$�O�I���7�x��w�R:Y�e�JP��x���5��^4��\�Ş��_�Q�\�9�O���]Y�xF� ��B!K�^ޖ~�ͺ/�nno��x ��r������l�7�,��"�1�#5bhʽu��\�n����j����S:qԕ�.�M�셈�54�^fR%���G�]�����2_c�| ���a���ܱ�g1�&g���<Ċ����)¿m�O�|��@�|�=�l�8����@jf]*����A�Q.]�*�=�����}��8ըSE/���{�xoO����r"?��;��E��@=���є�>�H?�SR�P0���Ã=��1w� `6��x�{z~<��΋���ߕ_U@����P>�M &����J�~G����G�`�
��ֵKr���:��t#��5�14�e���ݽ+��/�9{�������ll�˥�W��s�ȃo}� �֕����g�X���{�˟~��2���TMG#i�;Ct	s����Y�-���^ǳi�g�7��>����NH�a�g��j�:�,7��m��������$�_|���}ub���_~�e�q�ګu���:Fi�Ik�l�T�V,Cԏ6"fZO����c9�#��#N����~�I����|pW��*͚����QL���H��C���R�t�+s0��e+1VF��A�G���l��q����N�
�
c;8���t��"w��k�
�h�B�
��?gOHe��-��>����M��Q�����Π��H��Q���ۘ}#'��������~�*3�ś�[2O�ل��r�����C<�Ŕ(���1�,M�7j����P2��i�(���$ws�ǁc�g�g�b��ާ��S�WZ{�A���&����WF�p��}�
A;���lJXp�c���f��iQW��ߺ"f�Q���B�!�ʯ��Y60��d1&�u���	��܏�P�����03�(�� }��_�=�yҋ׌q�,�gZQ���L���h�zV�`R�������o�D4	�)3/Kō�	 �b6(g�
{�ҭ>z[ ;f��N��j��F����,�̌#��Y�o�BY��U̠w����v�g��Md��LU��`��݋TA�֥��F9.���$��-�lN�E�Ga��-���H^�U�������7�I[� _�o�m��3䢶_=�fֳ�O��!x@�2�Բr � �� �����P���h���~��g>#��p�E<�L�Q@��{}C&r@�-�j�W����B.�\ߜ3� g�i�Ts^���/!;h�%�ʹ`��)�/ԭ?�2/�S�=�O��ɷ�V��d�>�r��h�'=��Vą��t%�$�Rb��{kr�v�}�`��>|(C���κ$�B��ǻwY��{t �&D:���O�؛��&�޶)#x?]��"��Ajx��YW7�F!g�3���y�����ɷ�/Wn�Yo�ݣ���M���}ɠ؊쇃���Q<�{�p�F�~��dg���]/��K�&��kf�B�a�AT�� ���ϭT��ܟ��Nҕ���m�֥Ӳ��<��=�)ե���[�ov���Xf*M1���,z�g ��}9�s,�س������y�ҟU8��I���!��h��T�~N�{�0D��t�-j4�@��Usx�t��&��,C�L�Ų��������$�!�~� ��B���?nth�lG�-Mht;���yp<!����a�`�ݗ��&�_P�,��ٷ�ZR�!��z�]֯o�\�d�������H���(�.��T�߃R���U@��ޑ��dd��hw� F����B�ʚ�V.o���ܿw�t��hh���TG���ʣ�2�Z����@��ے���w�ǆ�ܻ/��S��R��_���p��N~�{o(�<�Z�[���7����?+�F*��U��*%]�
���;_����y#��ѩl4;���T1ԏf��G�-j��/Ȍ�c\�>?�{��r�H5z&A�|��d^������n���{lŁ�JD%��C�{it�rtv"�O�����ҵ���zGN��D�R��L7 S��bSL��4�x���yC���e�O�wcK
�B`��tc�3�7�r<(���2Kts�]��$F��Εə�n��x��fr|r,_�˯K�ە��#���]F�m>H�i�}�Ɇ퉣��[T*��5h����1�p1�b�&Ao�6�=NLd(� ����E��R�;*33n#�rq�RB���uc��O�u�G�L7�X6�6�E�7o<��%�g	� ����tWPT3�J��E�g��F��՞���˺��3uP�yL���D67Zf�V�����t��;�O�=����8|.D�����)��*�dg��*Bι�z�>�R	�:���z����Z�L*�ܓ�ha2�F�g�o+�.�/����&�
	A�j�r�آ/̬dn��!��I�/��9�+;�db�
�6�h~���u�ƴ�@��@�����e�U�8Jh`O���f�j�rW��#s1��v<�m��c�<}P�Uۚ���*�G;Ƃ�F���sR=�-��Q���`L�E����E8���ᒨ�1$��L+�{k�����L��_K�%ꥵt�j�mϢ`f4�Zf02�
Zǅ}D��*�#R�3��u�(@����=�q��!�፠[�bp���Xo+����kH�i&�J�2��E]:|��oz��c�K{� c���+l){v��>� i�;I�o# ��y�����g��z ���{aOJ�P�}H���qT��^y=e���i/�$�+������Q�������<�<s�8_t����>�٬f`Z�ӄ2[�x8���"�0�����S�(���w������r����{�#���Rz�PR��-�9zh�S.�<7G�@.t�s&��8���9 ;��!p���~K��u�S��;��|�2��8��-xP�X� ��8s�wn�3�t�e��|yʞ)c.�vW�V�������h5,�t���ǫ�93��E��:o'���y�+��[rY��aEchDg@ac�T)�B�� ��r:0���k$���j��9���HFQF�-Av��"rj�=۬�s���s�|�}٨�����¨���H;� LVF��Z��/bVfR3��X�.6�����%��"Ԝx�Kd� �6�j�>1��[���Pk�R�+9V�-���U��GU\pd��B�u�z�B=�����e�5b�ѡ1Cm[��"�N�ק��2�kEVj�	ĉ<̖�������J���]�Jw���CC&
ֱ.������t��g�UcX�CHfq�S=ㄺԣ}��:��0��ݡ�4�ȣ�9��X�<���$�S:�{��r�_g:w�T>8~,~���H7����������/��/ʿ���O)V��o|M����L�c_�kDw���:�s<s��`��j_-0�l3Z���r��X������*�rt| P�`��mZ-I��Y�< �������E4g�����)23�9��ڢ�n�
������}��2׵��R!��>m�|�fV��b*G����1�����l�2��k�;9ҬE�K\��|{���tC��d��Z�:c4�d��0��8R0�Nu� 8C���i�d#����� �L����R�цy�9�s2K,[��ޑ���2C���7Б�C�-D�rW��z�B�A�H�O�jn��ˌBh	TJR��m��fÌa����k�� ��jA�>h�cP$eA��u�;��V���K5pt�A�G#3�C����_~�rxr$��ݥ�o��u�n���[6�݂���{�O����O��|P���[ �uE��"����{\�,�|�!#��ʲ��{��>���8%�0��k�b�dy�YL��ܔS��8]�9u�����b)oi�Oc�7rQ����a�R@HH��`g�d'Jq�k��O��uQ`�ٷ!m.E,��O��`����T��7�#O��j��b�v��Z]޾$�'���u�Z��ߐM�7��k��\Q�:�<��2�l�E^��u����	�{���h�/	R��LLQ�/ʌvN?Ճ�(�p�P^'�Nь��_�\�Fɇ=��[��:�(���d
`����`t"�R'g<��dh=P&�����</E��\y�RG1A��Tm�P��{lF�����x�ߞ�N<�B�
��9����Y��{-挢@�����CV���C-���x�A\���C*�o��-�m�'�]-�?K�<ŉ�|Y��+�P��E��\��e�擃�}(�.��y2X?��Q{�#��v�0������?�zm��QTъO���CPB2!�2�e}�L����x"��5�މZ�ɩ�f
�Z�@4�(�Pg4�E�uv���:�"�����J��_����pbA��litR��O���D��Ȣ�i�0J)o5����M�@7�/2`�y6~��t�P�V�_=�"@�ͣ"(F�ò��v?]�xv"w�t#u\c6�V���=��ʇ�1b�^B�aͪ�w�l�c6�d�NiÅ7�yFyɐ�Z����0?z���'F�0��%�ў$uů�_�g���vTs�����0P���M0F48 >���	����,@Q� ��s�S-�/֏�W�S:dMg��B��kB+�13_-u��T;44P=��ۼ��x�1A�8��j�ht�,&�J.��?J
��;�F����C}�PEx*kk]O��YkQ4�Es���W�o���-�{{�����+��s�{]>�w��R�O� �AOs�O$�*��u$of2k�����smC�ݱ�(��C�������O�#7�G
N�q/���O�����%�[;Tx$��ypO����ʝ����e��k�k_�\�&9�S֛Y��&j��d�υ�����9kn!b���{z"�$�㣩l�.I�w��#�����x~<&�DT���Pn�����Ȳ#��C�3�F]��Kc�#�����^�&o˾�[m�s9L�����;�53sB `�Ǹp1���Z̴
�l�ki�N$��u"q�?��'��܍�Yn�rҘ���UIMdg2�Mme2��r�c0(�T!n%MFR!�2���tp"g�SRQ�����]���:�g\�9�/$K1�2��u ������"���)����𰏹0Z�Wȿ�_{�.U+���1�^Iσu�����h,-h=5%7o\#5h��1��^�@�,�bs����,3��C�]��ѣ�lu�Q1*Sd���D��l�~\�J���r�E"y0��/3�	����*V]^d��ǖYq��$(*�V�X��s-���+��U�ӌg`��:YRQ��ep]y8�TEj�>��)ɀ2�m�O�Z�L���%��ԁf�YAs��;��2��k�W�
��=��ꡣ�ŏ��k�Z?��ʤ���5�Yܢ����c �<�Q�>�h����S�%Ĥj}ٿ �_`=��?�%(/d��KW:]Z�QN��Vh5�0g)����t�j�JF5ϝ�8c�FI����2"�'&��,0���yQ��H	\sk�^$y媗�m���ꘀ:��0�o� 	�'[��
��F1��c�g�+�s?e�b����H^����~,���$�����P�4/[Ʉ�x���-I���wvv�"����t�	l"��XX���@X���T(6�H�b�?�����C��Ϣh4�8���U��~TO+s�|_�S���S��Ow�/:G$&��E��~Ȋ�$��9K���]^�f)��`vc�BX��3(�;�*�`��dp�|�EQex�:�T��,���� LI�A��Bm���@���ü�A-$��")'���$,(�4�9-*UE#æeA��V@tQB��a��ǳ4���3�x�P,-2��9?T" Z@ϥE��hB�#�ͽ���.G�@)V2鶠���.�g��F!�b
ў�W�e��QFaDQ�Р\4i� =��,�����l�m���2Z䁗������� >
�b��0��I��R&m-u�3��Qi$�[A4�=��u6X��G(�����9�Mv*����$M?S�)9�>������@O?�@'-��ͥ_A5Rl�:vCZ�
�b���P74�E��z�2�?�$��əܽ{_>x�C�\���B[W����6�m"ۇ{�#%,̩e!�3�1hn��Ĺχ��uzH2��h8�{hɽ�G
��ı��QGѓ���{�X�
h��&C�`����#�"3�4 �,,�,PZܒBc�b63��� �ޗ��[W��;��ZoMַ���7��Gȝ�G���AM�j: �`�u8u�v��
���|��7��
�v�$�i��b��+���V9U�[�i<�g>a�ut:9\���2=x������BY�"�^+'}p���A������Jr�/�����_����M�O6t�?�!���`�/�| ��>��R� =_O���x�/ǃC* ����.�3�jjv�q�q��~�@Sy<_
u|ŉ�@`E�Y1��7�gy�Áaz���E��z�W��ſ�Kg4������~몼��M��]�ƹ�C��`�i�1�ע#V����AZ\��h6��Ԝ"a1A'Ug�=S%t%8����u��G{�c
�II�Ei}ͩ-X�O+.1M�h�����c��"���1I��$ڗ5���9e�>�'^	����]��8����}1�C�����R����O�<�]�Z�k�^1G?I3��a4	�8?u��ӈ�q�/-�@�)ӆ~�!�P������޿�H�v
�S�hT�}�'G�[�3?x�@ں��5�Aq=�Ѳ	���p�#½��J�!d��A���Cf�\�����uK�ܶ6�6��Ȫ��\Q��j�d�,��g�j!h�[���MAi��F.�
��%tCC�Vj�H8��⹢v���Ġ.~2�Q��>����x��
�b	�E�P@ܴ4N�ݢ.VV��0H�ʠG�
Z)|���n��7�*� l���QAHc.�O�����F֖���S��\8S$��b���~�t �����_���Ja;Q\����#�I�[Q��x�%����	Q��X��!2"��QE;(7}ώ-�H��(��7��S��t!7������#V��pp��D�5��v������G�y٦ߤ�&꩖z���-���\���w�٬��h2'����(��`#wL�V[�%ռZɇ����FJ�)T�4��{C� ���hD	%�騨Š� c��MG*7c�"�eV�EK'���m�qn����,�2�5��:��׆:U�^�$��A&D�#k�n������ǉ��8�i�=�����U����ܰ�����Z�שi��jމ���!vѥ¢�Qlmq�շl3��@W��~��&D̂kD�`�^0�MC��D��(��s�t��������YVf�g�pP*���#C!���-]@eƜ�-H���-�~_6�]�a����/�W?c]^N��{��2�tã�Mv87�	� ���
Y�X�N�_l����aD��X��0#�Ɔ�uF����Ha�&����%y���%�߰�P?'�Sbu�p����]������'�ʫ������ϰoO��8I7���ѾQ;��;6�Ķa���P�wM��kW���+m5e�`�8ZȰ8���z���i��`.?�@݌}?0�I�孾<�6BE�r��s�Sb5���@��5b�Z9�(��3k�TPؼڐ�m9����������5{�hud9�IC��Vdvs�Nd������l�KA_:��-�G���]b6�z!R�t�H%�O��dh���6��.ˠg�'!�A�*��1b��@�_��դ�z�5fđ!NRoM��b�Kr��
k�co�`5��IHIcB{�
E�+����p%M`I,
O��1�	��{s9�<`�n�Ƙ%�x�����ݒ
K�u����P�p��`���y��\��3ۊ3c�E�^d[��:9��Iz���	�
Z�<������\T�wp�´�E|��U���D*��^.�e%�z���9���s��%�YT�za�.J��A*�#d�kO�I�#�J��<�G�
V&�5q���[�����$S`�����|����S�[�`���x���_ ^�@����)v G�="�p��l�q?�_�J\&s?c���0��\�M��`[��ֆ�L���L���JىKa�	A@��4Z����KG�s�<�� �DB���V��[���Z,�D��.�q{�7���H\�`k�\�\Q���Se4�Xm~$%��=������	���Z���.v��]�;PJ����U ��'�	42u��>��X00U��t �B��S�Л�)c�׮3ߪ����D?(�,�=�:/��2p�\V'Sm`�K��.�J�\T+�_��E��e?���o�jO;�F��B���znD�p�N�+¦�[�?J-2 �h@�>�<*�F�Ol�0c=wd�(-A@�5Iqf�8u�u��n>3���u9uP'�� ��%�ŊN�l6�FIIa������U��.����h�m��Z$�PBBW��Sձ�a<C��L'Ǥw]Z�V#֔,m3�>�qկ��ÄCq�[c�[�������U"��-6eIF5�.z����7�a��+�"7:O��'EYB
�7'�m�Kf�2�N�"�F��2���S�5�{&)�
�Q��zǤp���@&
9�*gcu����}�ރ�E<c��.ynoD���U���n��o"U��<��#@gP/�_HIg��ۖ�W��50�u55a|n`��> �Ffl-��M�'�8"_��bݬP������Hs]@〜� :F/��Q��6��X��f�� ��k�y�͎lt�r��W?���A拭!<�� �"
����%Db8�p+��=���t`^.��Y]�s���Hd�s�;DAe�E��ߗ�Ҽ�v�P`��� ;`6�Sd�@Il�r� 
q
�ڗ���K�ȳ�{QzW��a4��呌�)�c 0J/��VX�Y����@q�em�T~�9�ش�Ukq`�}�~�b,��U@�I��:� �SgzO�P�Ou}�l�zres��߆^k��������C�ĩ�#��ڌ�.g��7(H4�G�H�X�|�pQz��L�ia��y���L_����{p+/�2�ř�+n ��#���������88�C��w$�s���d��Ց���؏�3yx<��l��(	Y�	݀�������N��� X/��l���{�q:��ff��Y<��q�'E\:�19+mG�en3\D&�#��V3���lv��1N�ii��q�)1���^��穗֡X����#%���y����~K�yq���X��s��rg�!��@h�U!�=
�Q���Qꖇ,|��[�[�ߘ���v�������aY<�4����M���t /n+P���pR�Hi^��ٲ2��,z���xM�ZC�ݎ�O!�>TA'�i�b���H���
�޲$v�Z���jl�w�d{Pal��Jy�@��p���v<����u�ߣ���d��A�jq^)���؛3ğE�w��,qu ��N!��$���[[L*@ 1/�O��i��������.�f
@w�w�������������s9�m ��W6
k���f����^�r�J�G�#c�%���]��i_�!8�`���[j�١�=��X�z���R���t�Cߤ" �z݃��9��{} ���.:������G�fF_��E��ψ<�YaJ��& ���m��yе��H�iC c��c�/(&��^|�T>�4b�t�G��s\�$�P,c��Ep���̍g��ƶ�y�+ߺ�.in9�P{�+���hJWu.+ixv���#�S��9� t�X@u�R(�-)��If�F�P��Tg"�&�ȇ��@��DA� �h�)':I�vJ>;c�z?���`Ԁ!��Y�����xC��/��@	����u�����h���43�e�هȝ{S�T �??��
"����/�\Y�Ι�s�6H�Ȭ:ZQ��{V(�(�*8l���ڣ��fe]Jp��k-��ں��)@CftĨ�&���+�f��i��XWŒ���\>\(
7�[%��=7�ڏ;1Gl�l�]�����@6t���G-�H�>~x¶K�̸��r�{���>�����c����]����tvA��Z�iS��T�GcA�_9F5_��I[�e�)'�X��$fk�R:A��I���[�Ӝ�,�DD���@�lD�#�	:���n�u}*��<� N�:'�� @��8tu����xb�m���+r�g��_��������+ �Es��/0.kg�3��&P��pH̼,�����71}�;�݉�p�}�k�Y��e�q���c�ell�n�gSf����ќ9I�
���p0=�ÃcI��'M�N��XS�j*ũޗ΍��;����'�m N�`TzfnNU�L�
�c���̊e�dq�z֜{s�YE�p���N�8�rl�8w������cG--��	�ϳ�R��G���#y�we�d�>���Xz�>��h�7a���dEx�,�ty=���k@1�'ZX��)��e��Ү�xR�A��`�2��'ڿ��,L�0*Wa�9���E�gl""�Y�Nw=;X����: '�(*_��j2��v(l3�mYG�}kR�8�~�m��|�&�E��mn� `�V�{h��ѱ�K�Ҥ�6.��l���X�Y��џfPxαs����} D^�E>�U�~| T� q�tϝ�g�q���VՎNC5��2� �d�v+�@UA�J�t�D��d��e�>����(=������Ǽ�� �+�ZP ��}{�%8���|[��2��V���CrM���Vf�|ұB[��k�"�hmn/���2A%��S���})����$-��!{wzp"K��M�{�$[��9Qxsxh��0d�c�����D� �m���_���n`�b~��S� Sx��%���l��?}�G���E��2C��G���\n�Oпi�E|��{
q�<� �柕.<��,�&r�`�h4��r6�	j���}�
 &=�W��lZflM��W/ߐg��"�Syy�����C9>H� �!fp�(
�Q? ���mǿ�س1�w�r��&[�X<<�{G����.��]=���������'Ku[m9�{:L��wr&�NC�C��}'���t���ono^�+�;r��M2�>��Q4���}�n�q)�Pfbb�|(�ɉ��!���<D��V������à�$8݁U*�1�OII'��(�W\��Ksu�g.�э"F*8&.���h4
�()�欹�H���3����S۟�f���?��� 9-|#�I��4�ɉ^e��̤����\	�0�8a{Z1QQ�B'FLи�8�� k�r!5Ŝ$��fl���h��F-��_Hm�������T�#� .�k��/����}U����j#P�QÑ[�a�[s�����ꥷ���]�Eg���=c�U�p���7��K�`H��i+��D%d�
����P7�( �%�E�ch��?/,s�R�gI��V��0����i�Me�0p��o����^�g^�-7^{N������!�����N(��-	Y �>F���䖟IB��Ö9U~�T�AP��;��N�ӽ�O���~��:��4��E��\?d[�k�s3�=C]t"��B<6`	�g�Ŕu�}=�����I�Ϧ�����>8���u�zWT�@��3�6�z���(qZQ*�r�)̧)0���g��7&s_1kq.
�oY�����R :�,�`���t"uF�� ud�v�/rcs]N�Q�Je�ҳd�yNI]�R*T}�eY�N���
*�fyY;�,b���ۣ��������z4����J|��Q�kMi��Ki�3G�6s��JD�,�)��\�<G8.J��8�p�̕F��"a��|��	:�I���Riڻa�gY]u���֪�T96�w�K��[+�� rI���j��:�6,V7�5&��k��O:�O>������u��\. B��\�y���!
�	~����BXW�ڪ��ڊ���P>k��X��u�6�״׌I�j���N�g��G�e(U�r�	.������Uƾ��>A�h�9���!n+0o���L�,hIe�`*�)}��(���p�*�=,�{�b�3�з5��X�>�XZ����=j��.Gf��VO1Z-�	���q�Q����"P�d2jscS�W�qG��P���k2�������TQ������Z�A\��`��� ���i���PSȖn�x["{��G��|tn�)D��?99������0�V����c���PF/��5t���q��_���;�������L�Q�
��)�#��&�P�k�hOP)D�2�(vj�\&���{��0��$��Hzi���PZ�"�#��`�Dd.(��$��ܾ��(m��Nts��g7w����j�2��~?V���'�:@����Ng~:�h��9�?���ǖ���\�~o����#I�$J-��-۽�nc0��o��0�� ��a ��1ڽXj�v���[��v�%��s"�̬b��D����(V��{of~�}�ŉ8q"�Ne3��L�{�������:�?���in5b}��o�{M~�_��𝿖�����	m�8A��čGκ+3w�	6'}q:��*�:��j���v����r�,��;.m�4�^z�΍A��՘�{�8��W��Gڥ���0ЊY�T�7��|GFa/�JA+!��?��D 0g��/�\�{=�� ��%�:a���h9/����8d5}w W|�v��@Am*�U�n�3��>|�E� b<u(~�����Ξ<|�99y.�j�7���~m��{���b:1ꮾ���o���t��o�������ܗL��&/Ag1W�~k�P����������b�"��+s�����)ͩ��166��P��ei�12V FQC��7E��$� ĺ�Q��VTsQ� �y�T�<�d�1G�P��f&yKϾݒ�{�e��[�;���b��)W
��z  <��z�u�Y���f��	z~Ȟ��ZhkOlk��X��"b딨�Wq���[���Ԋ��1Cf,
�x�-��u-�"��Zl��x�L͆�Úga?蘫L&h$<�����'��u�
B��8��Z7��J ټe-�N�^>c�*﷔J�����,�����I�>��s�[�	�	�0�a����0n���%���P�4��3��z5b'�}�h	3ǽn��h�r%�9��E��A�O����ٹ���w��599=�'=Tg�$����2�������3{�hOE]���g��Q?��Y@ r�b��h�1��&�]ϊQ�?� S��\r�\� �<�yk�_ٙѻ��a^�Y��� *�����,pD��W���={����<�y��>����*������P�6x_⭎0�k�]���{���o� a,��@��H��z��[yy?��5��p��8b�Z�CW�����m1�����!���f��B�
�����~�:m���&�|�b�Cڤ�� !\Tm���z��Fm��|���]]�ӆ�R� ���[N��#�-��������<�=��6L6�X0c�o�H���ŋ�WP���e�4��./�F��gx�!��j�+��Kc�q�4O��E��~2�R�.��A�u:��y=�9��D�%�4x|���Ļw��3�T�k *Q�P�m���'+�&9Q�䌽
qχ������QQVL��RV����0����ҿ��m:~	YB�U5d-CaT��L�Ŕ�O�s�ɇ��w������!3h�@���ahI�\=��UK`W��������A��ݓ'��?:}!E;��l�$�hO0����e�B�Q�H�"�m�YJ�;��^�Qw$_���L�/��Ѯd�h,�g�������ӱd��s1"C�/R����%��3iwSv�^��4z��
2Gj��n�׎�ˇ�w�g��-_pEp,#Ft�`�2���i�����*M�A)-C��4D��A�c�ׁ��c!��L}�ʐ�* m��"n��聅�F]z��#���/��IJ��gi��l��2:6�EOH	��((�zV/��5LY��	hWQ)Ȓ������o�uX��n��;��Ŭ���0.������@����0��/9XF�0\�/�c�7s�R��ʟ�ɟ�7��U�7���$/���y�)�:� pg�����+}L��  ��Vyd�^������/�
�pŔ�6e����`Kv�#���p5]��"4��Z�2�QYG&Y�4Xf����s\����
9KUG���-D
���9�F-�BinURD�`-K.�#���J���~�������ݛҹ�#[7���;�E��Yf�(J�9�e��Ed�F�?�3��,��/r��V�zh1��#3�t(ڤC���K�}��sp����b^9"��ⳑ��k�p�\��r�^X�g����t\���[��M�F�b��kY��d� �Ε��ĨH�Δ��2�~�PǅՎ�
²�bąw�����Z��z(�j�J�

��2�Wi�cÈ�!h�1�[�{�:�?r�F���_}Ԛ�2�2PX����y�oVl�t$��~������-9~�D��c��:�VOL�DP�RO�4u*_C�la�@��(��t4��� ��H���e�y!3%� �&Z��ƿ�˯�@!'��, ��g�{�Vt�����uK�U}ðT����!Qۍ&[-߄��>�^RP� ��]���k`�у�b�+2[XI�5�:�j���b`XP�xށR�r�Q��`>_�����{���]�2�S��썶��ݗDv^U��b������}.�A�ꇞ�l ��cԬ���*P訓_�&�� #�]C�2�C%�Ԃ9a�E�_��&Z�N,��i��tYչ�> ,�.���iE�L@3�v�<.�T�[7l]��L������AKmb���Qמmr�5���3c�k3��@�.B�7������.�2����ʨ;d�e6���|JFX �X�n/�*��z�y�&�z�Lc>��M�ԩ�����P~=����,�7��T���;��[�{!m��0�r�g�_wu�S�?�����b���((�f�G�3�X��)f)���+h{�P������=uB6�t��Zd�X0���g���6�O� R�W��sy�|��Z�\����nh��[���[D��4��ee���w���Ek���H�ƾ��TA��>��R�5ؑ����nt�:*pSl��h�˰�+�/4�:mu�Od}6���ܒ8ܣn�_�����7:��\��M��H���\z8�zm�E��ۜf3�}h�-�'b���׬D�Z�Vi�؜���)b��U�b
N�t�m��y�p ���PzN��Š�X $��FE�(�E�#f)�[{�y�U�ARJĢ�e�rz����S�J������g�W��x-P���g�!��Z.:0����@gff�Gt<{
TGm�o-T�m�M �V�O쥖w�� ��PG��!I�X�)���"�qb�Ǭ�u�>��3�n�3���}y��l�����v�'�͘�,�����g$3���:lfP�L���5��:F��PE��Z;#�(�b}.�S�'�v
$P�g�4�&a�����%��G��_��\m���>E�W�qJ`��R��D���[��g���;o~���V)����F�Z�s9Y��2^���B��TN+Y�9]��u�h�����t`��r�W �m�*!�*[3EpZ�G�>@���n�tI�ՕV�"#־e�hut!�㫒B[Q��:�,�ֲ^�չ�(U�*�TF]`��Ap�o:�/�@��
�Г&3*(l0I}E�$���n�%���bY`ot飠�-:�(�u��!��ӹ��/d6�CZ��#�>V�ӛ�D�{�Ba�<���jD�U���Pڽ�lom����ܻ}D[�`B���P:��/Աl�k��;2�1����ud�Ϊ�YM�����u�������eR�`�<-^�\��r�c`DE���.hc��
(�e4nfCV/���#v`YO���֯fxD��{m���C}��{QxF47p�,�ٱ�1ƅg��j�۴R�����9��٤Z�.����������˲q�v�K��(:�2�ᳮ��O��7~/�H[e�Ô��??}!'���bc�K�=E�;���-�Ay�gm|�FR��z����K��=�� ���P\-��7�W_�Q���n�M �ͽ��>v���+�$H�baR�:�V�׻����jU���yB+��q-�y>�I��YJ�8�W��e=�K�b��}��,��[��;�_�%x�����������tՏU������XΎ�X�*(K\�����N��jo�eW��PÑ���QU��v��6th��Z��-,�0�O�F
�Y�a�\����-
����W��(!���U@��mV�g?�Ez��[�P��Y����io���N���G�wo�X^���M�1u�@�Ihr���A�C�:"�Qd����N���9�>F	�i��׿*��?�;�=KP ����hŢS2+�����#9�g�rBL�57�3�����Y9Rp�?;>�V��;�����J���e99���L��7ޔ�N��>��]�[�\PMI'�nfp�Q��~8�PH�]57�X�k��P�qO�g/��@���x��� �P��vZ�����j���c
N6�x��DtQ�����v�	�g�^�O:[d ,��H󀿐2+5Ls^�x����}�;� �*�%fQ�/˖662���olp�V0HÀ�y����V	6j��x���Gp���ǌLو�~W��(���Dv�����_�t8�k�H�
g Tȸ � #��(0xu~ J:Tc~��jKfp23�:�L/�;?��L�m�|M�F�g�(`�b+���ņ��@��K]N�;����*���u�^r5�7������m+XZ�9�f
P؝u�����7x刱GR�v--EN1��>�TV�bQ+߶l��2��9�Z�&]sm4Nl�:F�ww�����$"E0_��y� :�q�d����T͎e�و�| �?�M�6%��@�F�@MK,��³��Ba<֝^뤛4t����=�
�J��
�by�Q����Y�4��¤��:�ec�w��?�٪���Z)�kx\���=�d��Fx�y_a���\-�t�세����>k5`�	i ����+t�-#����-G7�8�z:ۜ���S����-�h8����E6}K�(tz}�ޓNb����C���fQZ�0Ȍg�]B`  ������H����k*��ň�Su\@Ion�!�Q��m5�Y�\��N��v�Ktl�ՙ���)�Fnǟ~P��JWP�z��]�}�c��d������/��Fkf#�DkJ���+()+�;j\��18��9�(@	_���&䟤}6����)%����<8�	�A�WҐ��}�=�Ww�Մ<������(�&#��o�U�	3�r����.���Kg
H���Ȃ�O'�����'"󂭙�hV_�i�����pL �>��`�����s��k�DA`��R�D�J��	
��Z3x��l��%R�ٕ�=h
�ՠ"Z��4�!�VHx6��\ѐ�l�#��g�lo��ْ���ؓF�+�-��#S���*�Z��l��Jx��G�)�Y��^/��{�:�l[���;7e��;���B���E�j���;�*��g�裤V
R\�w]����6���rc��b���;Ū�>�����f�rv.�������Go���T�kO^yp�=éz�����@��A�֖�B��Jt�O��������C��fW'�jo��G��S-r:KN�n�E(dG�Ȣ��pʕ�Z�؜�ӦQ�-��9(��Z�n:���H��}ف�����%��!js�ա^�(�K9�gҞ��t�ej�J���,d������6�.����e�̠�%�N_擙@�!_�\�:>��dʚ����*���y��n��G�̜:7h*�Npv~@����aҁ��~p�L���+��O����#� ���[�T�+_���[o�%�O.&rv~
fGv�{p@i⎎8��SW̗2y�Lv�
$Q���q`�z�ȢYIUDX^��?/�T8 ���OPd
��G3�d��t��##���,:d��:e�O茚�2�h~�7g��雟\�,���dE#x�%�΂s��;wM�B���]u~�H�d�>���yO><�|1���P���W������pvz�{ �3�׏�Y"�u����|"o������Y3`�S��$��3�k�
ڦ@���&r��m�������`�z(���0��h����G��{����8y.�~Wf������ύ9W($�*(���v�b>�	��1̃�(�7�j"�p��ȿ׉��YU��\?PR�f��� ��GϞ������>p��������}F�����<�,;ky��ɤ�ɣb,�^TuД����M
�%d�=��DM=����Ѫ٫ɯ��	��S�(�|?�*����USq���X��Bfd����0�g�k�,��E}F5Ц���0bˤ�_O�ܳ-���r���56g�5�_a���|�2d2��V����9/��Qx-�Β�<E�Yݶ����B�W�y>=9�s���/u�\�%e=f[�_'1�_�WL:y��!���xv)a.tJx���Q�X-7�@��U=]�m��c����@Q�c�#�>�h�ۦ�pI�s���;|�p�E�Z���ڹo*���qm���ە����D)�(��V��5����OA���,��4��~�
�Ť�[m����P�;T�T��{�C"�ώV���P��0���-��zJ#�I�I���U�����}׌u��k s�F>�f�+z����A���ֿ��*x�(�ͯ ��r�~y`
~��p�m=�"pƅ:���ۋ!f+ [,�Z��Ԣ׉E�t֥�q�����X��@HT�'����(�@GcT`7��.��e[�5���@�X9�[�`���e�h�)@����n��v��mr��Tw�RWǄ�C0��@+r�;��|J�k"�y�E��)+�	>�>Z]��ɡ4Ժ�Iy�"�bko[^z�%
�<�xF���=���!H��`�ur+@��jI�����w���B�/m�l�%��k��VB�ѱ��\?{$S��P~��,�7�)w�޶2��CK�k���& ���l�+��㺍�t�
J��v�*E�EF�a}��[���ݗd��o�x9'�8SG}���8涓R�$Յ3��M��ʩ>T�@-������B��sH��ϓ�R�<����<oI��*�#]8��\�?{�eJ~�H�}]��%8�mF��Ɔ��Fݑ.�d�F�b&�م�W���I�]�jmL������ܸE·��}��˷��u����K�@{�J�sQKhM�-r����Y�@0��.\ϡ:�w���_�qI����l��Ѷ�v����]:R�Ι|�Ï��g�ud
Jؙ��Ӊt��xЖ�[C�nֲyz�^�8�+u��͎�j���I%�J9W ސ�Du@�u-�������YfLB �ꀚ���i[�T���0�mn��-'E6�	~��KQ�4�Ћ�6~��#��XW FߋL�|���^OvC���9��da":��'��r��Υ��'Sy�G?��dN5�;
$�{mY�Wr���f�^9��g���g

u��k�;�y�[B4�����|Vpto�<�Wt���= �Ӳ�}*pa �QL�Q��:��k�ʫ^�5������LHsD�w����m�b#AV1H�[�flmT��0�ac	A���G�G�hF���n[+���bM3���3�?���ˢ۠"���XpeU���mR#���f�tG�G}9�)EH֣XVmݠs�,�i��v��@H��A�Mp���/�!'e]E�����7`SU�䛖~���B2���2��'��Z�ؘ�,.Me�s�jN�l_f�,5�DQI�93�����~J�װ�~�W+��2��}Q,$�A�'m}�2U�|*��RӉ���Ԗ��:s���Z�d	F�D�_,C�^{W&p�=`)�Pj`6��%	����������Z-*�L�գw��B&�e Pڐ&�P��v�`kM�i��ƟT�+�%JZ^DQ�a.�/�q�lB�v0r]���J�(BV�s������!��Zm���A.C`�o�z���i��u6�/-��+�q!v��4"�,�k�l��ǡ!}@����&n�Rnى����)#]4�׆XOpJ<Cj�Y;�ʨ���@��iGY.�E��{��Aʤ�"�Gn��x�-o���yso���;��I�����U���j�R{ZU��_�9�:{C�R�������A�D:jS��[���\�V���ԁ_ʰ=��t[��fr^�d�:�"���6/W2Cp�z0�lo�� ����9��
�\�����ŗ�,i��W���Ԩa�_���
=��o���/5����q	�_�#lĻ@��A��0���n(%�|?	���ғ�/Q]C���"�Dз����u�{鮜��ɻo�/��sٞ��Hd��`4�Ɂ^�B�7��;-+��6Z
�����&seJ�\Y�~4Y�եCY�%i�?�GO?�?�PNǧ���ߔ7�M���?�Սo�L(*[u�|q\j;�Û��e��&����jxA`�ۢB>^�Bw�mBl�}��M�_����P3��TCBT���HvH����?aVb��X߳�%��3��$��T���.['xsN�������3��G���'�ҁ��������O���_e����HO���o�;�넼��/;���P� J|Q�A Ml��ng(��D�7�2W�[�H�ǂ!e�{k$�nߐ���|��Cu6�rxp(g:1�z�R���~�j��Lf^��w+���,cs��x�A�C��h.��RF�>4���Ӳ�w����#��K����>�c4����ҿ�1Z����W����a�;�ɽ~WV
:vG#�\�ñ�Z%m��E;��椟%ܶ��+��[����tlQ3�FBS�زy���PxH̴�FȼF1�׾QZ�xP�#gQ����k����L�;Ib���t�����
/3J#�/2G tc���\N��ˏ�C5�C���UӢ1dTL7H͗�$�ꐞNƺ~��t��tō�n�g��w3���h�4Z �\ǭt���t��"c~>z��V�X�(������?����DF�)=ڻ��a{F���Ϝ*������a�,���~������*��, �
��L�Ɯa��#�kY�i��}0���[R��yW��:�Ye����1H��s����5�̦���u$��|�$�	0�Gu_O�j�Z�����!�H�UUK��鷲1Ve���e �ʷ�"���/eŁAE&�������AŸ4a�A��Ȭ��q�]D�������>�hQ���.�k�#��F0o���V�� z4�8Ѯ��/���<{�\��������B=�g!0����=���N92@�¾6Z�`��%�ϻ��k}����v�I���B�N4����<�;�������Ƙͧm�Ԯ8MP(_��o��#�/L� ������T8@V����P�"�.Ue�pK�/�8Z��:�}�!ۈϓ�甶�xzc�����G>fI"�1�̕&He���H=�^&�(
�)ঈ!Ĵ�vJA��*���yD�����)]�-�pSFn���RWR5��;��"��j�+���(��04po	D��]V���G�95ı�"^�Uz1^zI󞜯r���Ų�� �����×�f/���D�������j�Q���V8��13�V�2�4�K��
��cWZ����h�"u�������O~]V�,��~y�3>}k,}��aNK������R����Mq���])GQUnTx���\��^��.?�n�񇍆��Xf���%����������啻d�`_�����sY�^�1u���V*��9DIHP�K���̰�kC�#��;WLqrq&O����gO�rz�_w�ߓ����k�&�AYC�/�W���=�R����N��<~�X��S�}�Ҷk>�#u|O�r���e5Y������'r��m���+������ʓ��{t[���TA
"L�EF�HA_�ߑ�u��ό��������:��^��tx��ܸ}$m FL �H[�\����͘�/�}A��]u��yB��P�����s�|�n*k�lM��G�D�P {_ŏ�zK>|�!�)�~[�-Υ�u��i�,�p�/l� �����	l�jF
�r%�x�yp�5/M����/�MkP\�ow�n�����TR�0���� �;j�t|�
4�N�����0ֲ��&>B*:�Qp4�#ˍj��7���s��,�{�Nu��S,t�ȘÁW�mm�B�h�8:�Jc��d�9U� ��*D�j*Ut�zS7�'��r�ȑQ� ������C�w*�W�� ���MV:���*2�S�{D�q�HF{�|�0Rc������=:�x>{�y���lK���|�Km�J���Ǿ@x��Q�xz,;��L�Z#����CJ+D�Z��K}�'ϞJok(�f�� �� U"S��\�e��a��R�7}���	 ����E��ZM���� �=���Ns�Q�LR@����vc����2�w �V,/Ƨ��7�����JҜ:1���C��X��TM�m]
�����
��1A+�T�U!Q�e�:�L$��Z�������̡
��8�u1�OhH�����s|�v\
�� 
���tEи�%D0����X,��T�n��v������c�'�Z^I{-�29�1��GK�B�⁎��k��VP��@/r�BX�0S��,:BQe��5��$c>��tG=7�d%DR��B/�I���<YS�Y/X߈(2Uh����J�E�ò����	��0�Me/���E�1���S���b	A������\2*WpD��B\@ )��9�N��쑘�Tb�/z S����h;^!P"gH�D��ȯs듘��H;2�^խU�� �ˀG��"2��)>_��dw�g�Aԙ#�Ct�k"6�q��`q��xN�	_>F���^D\��~f=�� ����,�:�s��u�D���G�:ǈt���V��F���VT���R|^:�$�t��W�&g

?~~!Qw 7ﾬ{϶��/�'�~*�~�G2Q0��� �l����Ee��@���I�,��Kn5�A��������\���Juԁ�'ĥ�����V��@o^�j��/�ݮ�hvu-<��*\�'i�_$�_�� ����-�}�6�ɠ�q��\vvvx�-�à�M�� l'���n$����Gr�oT�LߋF��m��^��O������L�����gL6��5�~�K"HϖEŕ�@�1(�~ �G
9`�b�Į��
T�B��GG4���Bv���9�� �o���?���c��r�i��ή���>BVt϶:�:��,��\�N��#�l����d��������'/�.��K_��7�D��mo����DAڠC:� �Œ"5菆�+�Do�'O��Y�� v�1PGp�U@��#��<�g?����ψ\�?Z��6�O��;�3}O�d�^*ݐGM�]=o�0��m	�Mq;��������i)�UJMp�3��Z�T4x�BA��'��
�z��S��yM�5�@���ŸX,*%R���7�N_�؎ �`�Qw�.��<	U�Jw��p⢴��ep��.�
�Ѳ�[��q\QC�*�zf��r�ĵ�g-��0M�w3��I�ح3k�J�p�����J�&�s��5��A����H��[��)�������gj���.{�!�1"��C�v6�Z9qap���~ꞥ.��< �6���d��oHG�T�Ex�~��ҟoI�=��^<'m5��a$2!8�p�2�H kB A�Vϑ����k��DU@��FW)�����*���Hr�-"�litb}��J�n,[�wd��CIn�E<���n"�1�2���^ �֥m� 5%�������0
�+!`��kP��H�I\5��cQQ�i�Foy����8=�5�
�����$��})����ld�����f���a�-4\Xn}K-U�`@G�ҁ�����f˺?;�W1A,�Oˤ�:py���L?�L_���g�nd�<ӹ(һݖѺ�cm�YS�����C�Ih�ڿ�:Ơ�jY촪���� �p��#EFE����f��}��q��ռl��_�W���8���~��Ak��m��C5@�/��SV�m<����nʪn�A@n��!2�p=��ZQA�ځ�`�S4"7|��>�[�1/�l{V�G�ll��Pz��J�s��Uka�"w{�T���K�M�[b=|l@�
��+�0x�ѯ	0z��_L5ľ|�r@犬��U�p�-�5�	����*��'E6
��ql�\��t��F�jg�s�}NP���{q������PZ�{:/S��O�7�E��{��K�����<?{&+(Z��~ #+����r��O��_�Y�����ؐ-а�#<�b	�S�+|���}�]�%,��xBs�>k�Ǿ"��
��=�2�I�"jR1���z3���@Q%�
��z77��?��)6�B@��7+� B�moO����H�{�}���˲��|�ým�0֘WYW�%��i{cz�"�/1�"/��Y@�lr*�T�=�/�ѣeq�{�/�տ��^� = @*�G�o�#�8�ȥq��*��_��:*�����o� �L���%�c��	v�rrrʨDa� )����\^�N�O�⅀ʉ���E7n����tw8����\�T'f�˗�$��.�߸#��O�?���@��ؾq�%����3�~+Y���P� U�ԥ�S�N�:'��G?��T��B�ܽ�M
ZHU�h��m�Y���Ï�Z���ȝ[7e��3)w{���Y9d#�*_.�]F������tSA���P���ʣ�ɶ.(�b����Y�uz����X�1�/���Z��X�xc�0�9`#S1Y�PMhTظ&x�0h%�1RXT�t�B$��^ӂh #�F�58Ȼ�������,/6��廒�2��t����i����щU�.B� ��iL!1#epc�N��1���+�:	��G�yg�8ǉm�؃�n���D��D�>~�Ƭ�ǉ��?�P���!��L/$���5Vw��$N����
!��;��-=�p�*���S0��g�,��p}'�g�އ����F�����X�$
�a�Q��*6U!�2�q�^`�����ci8��q /e {�+�&�sF�%��\��d��sǲ8�������5�/���� k�E�tv�d�w�I��=y�^�d=e�&�&lѲ��-k�1���9Qn���γ �ɢT8�=DN�M�ԥ��Il��6A�"?�)�Q4�E��t6-AQ��L���Nj�}e��A�%���f<e=��`J��_���\%���F�@s���lZ͢S�G�.D��a�FXe�<=l,bs^鬄́_{����{���	8����5��`�Q�U�����҈��,뭧28��"��)[�$>W�l}�+m2��J�ٍ�C9<ؗ��=���l;A�5����K����;.m���AA��� �2�686�
h!�S�:��L�Q���;�c��2|�&��/m�Fn�.)2R�B*��e����;H�\�	4P��Y���j?ۨ���޳bb�K�X�`�F�5�� 
�V0s���0ϯ���\Di{�� ���(�^�m8Pz�]AmfYn��Z���IIP�#Ѐ!҂�2��u�z6���N}5���mH �@-�:c��o��]v�6��M�ʗ�ݗ����Ȼ?��<y��T�v�2W{�|1c����i�L��T�b��"N��[���Y�EQT#�ܨ�o���i���\ \�]�V������	�j�.[x��8ֵ��&9|Ί�]}�gl���f�P�֘�~R�U����y�i��v��FP�ӏ���6�n��W�D6�$�7~�y���,9��d��)�9Mn���%��Mէ6Ӓ~x�Y\(|�2W95�?� ��ɉ�X-��+/�����Ƀ7^� �t0�����/��U`J­��Vg}/�6�b���o���Ļ�L�A�ΤK���1Yg��/���נ�mq�`H$�R_���#n��������Zd��hoʝ���������k'ƹFf�4]d:ԘuՉx��=��׿&o�ސ�'O�#u����}pC
u��޸!g�Yá����T�~����@C�im8�w|����]n�ڧc� ��Jw ;�Eߒ-���}@���;�dW��'3���"�����RCry�����o����2h`�F�g�O�����l�ي�р����l���qݞ�r�e�&s��Zϭ ��KK?��k�D/�GP�Bq����$y�@��{p�	�À�e$Bq�x���
dG�	@K�c������˺�`��}Eà�V��/D�cW�2R��*��-�<C"QMw�2���$�98�n�j��T��4h�,�/��c��3b�r:��r>����Q��[?y������@�!���;2<��8m����@O�*[-�ܔd�*��c[v{�ឭ���W�u5���{l��5���,�:0>���K:.��vF�r5��>�H����	Md��:���[��Q�@���CQ5��8�*�=𬉉��ldg��"�1�ZI�i��4����9��f� l��vj�޽���7^��-�h-d���Ƴ4ʈ^�*[̡Nr�(gˊۓ���)o��48^#�4Y�1�5�Ft�Ԅ�$(%�Ao�E.��@i+�YY�(D�I���\�U"���3��{l>�Y�ۢw萊�h}�Lt%����)�1�υ�<�̳�I�V�5��*�:�^�8��&��]�r�QĞ���� ٸ��rV:n9��n�ʛ����n�>K�ɷ�q�w�
���]P�l����K�J�ĸc���zB�廇{��z {�1)�C�Ǡ�9p��zT=E������q0��Wy�ۅw8Xu�T2}�9'U��9���&m`�To,��y�&��m~h{��~���T�@���vr� ��3�Y��kYÄ��:$`2@R�m�ʠU���4Tj�<�k�iT��ʏ�a�>t%�[,S��^���g�{�wǶ��9�𞘢=��q� ��l,�O\S��9��!�  9u�/��/뺏�;���������������'l4v����x5��|F!'�\�ҍ[��?eD�����rR��j���+2Jޑ�$��~Q��0�� � (��0�粯>�}�eU��
&ERW=��}���P7I;�`bfk��t��06P�0U}s�x^�!�e��a��%%N��
1�vO���,g+��|O����ͯU�y�=�Ay���������'cI�	�,�L�.a��8�/��g�X����S����S�/X��ʃ��������ޖ��7��&D��G)@c��y�*���bk��Q7M6no0
����<} �n@\���BK>�-r������&���D�����o����'g�V�N�"�6�~K���~����-y��?�w?�P�O/ȋ?_�eK��͇��&q�Zʏ?|G֐��ʩ)��V ���ڀ>8�e}�F�ғ�� T�Q��WnW���Yc�����ν�2u���D���#j��wn��\1U���q��ܳd��W������	=X���Φ��l�7�d��s��??=7�5@���`oO.�괨ӻ�3�ϊe��EԱEb���ް�0�7ˏX�F��P����B[՛���>�?���)�:V�]C�5�z&�-ꠣ/�p�SFCMn�z�!+�⦖m2�#�#��8���e]3�[A�,W�3��a�9Ѯ�&�`�$��a����⹱��4��������G�Ѱ/���Q��)jm6+�8?���N�^*xQ�8Q0��1��%��:��T���w\� �W'5_�L7[l�͇�3�H�>���ܾsGnPH��wb���*���V��Sy��<�x��@	#�b ;M��\	F��Q�λ�d;m�ή��嘇��J!��y�.��m�ƈ/�� }P�{g���MoR7�yA�8v�)�ِy��Ν��O�$����l�\�c�Rs�l�,e�+܅��b�%+�M����#ZЗ@k�(�7ӯzl��8_�~Y�����M�k��djuV4z�l�0���m���k��Ҁ�a$\�g��Yl�>1E>l�A�ې�]�gS�"\w"oZ�ˣ�Q������8;P�=c�ݸC���H����;'s)�ֻ(x_�f�=��al6*�f��RG��ʽ'��������}�X��2���H�voH��la�U��_�~�.��^�BJ�,5�>�I��di�f	�D�V�IQ܆� �T�*�`��Rf(8P]�.U�̜�Z�#��D�@V(<�+6�^��&�)%j�-&�t?ˆ%�t�s�Y䴆�~�߄d�uG����Y��w�	~NK��|X�{��S"��S�

���_dK��g(��~#��pbf��'�3���O��ј��kfA.���|��L�w_![fwwK�~����פ�23m���X����Y���Jn�8�Ӈ�_�Θ˿����@]6���c��T��k��IHk�Wj����X.n��W_Y��s�x�t6|U����o?G��Y 2/#gNY�-)�}���V�\E�����ee�b���g��o��D,	s b`w͖q҉
�Z��G'/�}E���/�����?``��ɉ�8?a}!X`?�s<*ݦā�7��ԗ��G~v��J���7!Y�o����������~��V'���ra�<7�"�۹�ў��GP��6����q�q���{�ҵL!x��f!�6U�Rx�H�!EL��>�Mn� D�#���`O�2�	�jL������b�V�
⎬�"��R�y��|�♌��\���a{([
8[:��<~��\�kDτa��D�Թ~z�\Vӱ��Z@��p O���'��	�/VpK�"a�0�l��hK�
$��j *=��
ܶ�Mte�P�;�cꪔ�b�bwP%�:,C4r�M1��*X��^Υ�f�+����m����]�xL���mdn6����ߣ� �nT���r24�Щ�֮¬��x3��̓�Ün�m��ٿ��3}�Ǥ�ZДR`�Ѵ��Ç��c�7ӎX�	M�*��s�q�,��裟5����.���@�P���K��-�����~h��Ru��|��">	k�R \D�ڔ}`Cod��$6��l�#VPs5J-��>�^c�kK���B`�k������P��d���ܠEb3�&&< �Ǐ�3��C���E���	�@ʚ;dx���b�ۢr�>� \Y]�O.����D�׃�MB`�$�#��8"�I�2y�x<[�c�̉�}��$����o<���]y�8��� M�?�qn5�X�Y^8��/˳Fr
�g����P	e�B��Q\scϫ��x���+\�B�w�!�#g"4�2*W�tV����מ%��������=��@�������;p�A�aay��`�Mn�E���k%l��c~�a�v�%=ҺWbk�O:�]�B��0���1�@7�W��e(�V�'�Z:�!~�+0�Y������:�v�2�{��uv��쥣�t�@<����+uJS�=�L���br=f3L5�@�VΛ�0F$�rm#�P����x�ڿ5e�� 2<�Q2h���\��֋e�p���d�<r��	��·e�ː--�u�Prj��! k���#r0�k=,�)��ǈ�����#˒�.�§�� q&w��z��˘%K����ĤL���3��2��2&6.�'�3̋((W��������t�R�J�ҡ�0�������Bv���Qf�3-�+����E@D}�M������b	���R�	�Њ��	�T���/�I{�����Ac|��԰7A��,f���>�,�r�����3�ԭ���	�r֟G�_��+ �_G �$JPu��] ���9%���.�L�2�T�J�M�k؇�j7�迻2��>��s �������Bҽ����.gky~�T}�)�<I;���X��gr<~.��9�]3UQ�>�G-�>����	��b�|-����?�c��߅,�5��V�����/����O�=��aY��>�e���|�}Ο��2\����`��y�Ne`��z�����S�O� Ҳ�Q8E�s}���K��cAB�N;��ѓm��,�	�=�u�I)$��n����g���Gg�x����,Ʋ�1��d3��N<����o?��K��u�sn�U
RЎ�T#6O�{o�X�2��F�Č�'y#�c��� ��_P��k�*e����|��a@v�P@	c��Le=_��%f��YDˉ�2�#i�X�#�w��B~�u�{z����Ÿ3�A2�$�Hbu5�u(�4��C�$c-Q"�B/=PO��LY
X R\D��0�p����7�Ag�] ��RY�(ԏ����_ޤ>i��`��Ҹf������EPG�HJ�p(���hl���Md�L�d��0۝=YK餺�'�~��ξ| �F���b��
��m5t+	�
����|�a�\x��li
�h,��$m[�n�k��  n+H�*�N���T�j�QP��y?���Qi4��|�l�8�����gP?}�Ҽ�"g���"�2�_���l���S&B#�\9o"�o���4�VޖV��M1b!�n�"sd��TZ���69�q�ȭNA���[r�՗e��P����b3���kőIu@ yYͿ�tl �������J�����=*��C���tҽ|����"S���v�fe48S`���Ȕ��T�C�HȰXK���!�����T���OQ�S�*�,(Θgl�[��?�obϮe1�*8~]�U�]�,�/q�Z|���@�G�1��5-�yL����$w��J2�}�	����
�Dտ��"���6!-�٪���zP�U��8���Z��[{C�zB�R:_�4'u3��y �В*^_el܎A��Y�U/D(�:�sg�a(�,��}#�2E�fK��6�sH�ĝ�y�O�E,��d�ל}6q�� �*`�	;E�xY��U��n|�W��-!��9Я���D��HCkyiYz�Sکp���=A�.m$s�[�g�'!��Ao�v��=C�)���ɫlcP��e&�y���|*<ޠs�R�+Q?e��b����Lԯ۟�ɍ�=9>9V۟��h$�^G��T>�81���,����n��γS�l4�G�BF�Y� ������Za
�ܸ!�ސ���|A��jw(���)��m����8�>`/t��	ŭЮ{K�T��d	yk��=������T�C��P��TJO�+Y����Zh�ӧ���Y�[XSU ��߮y��w.-�O\)��kB�a��0Oկ�Sf�.��f�(��c�$k������L�SOL��!���6�n��~��r�֑>���t�$���O3К�b\!���<�O�	\�B�֢��+5/���ްEN���N��C����srz�P&�����)��Bb�G�����h��Oa�;=)t�%;����#�$�tC�~��U�픵��K$�� �'�	�@UE��J��x%�^��}�M�%����}WP����ˍ�@nn�˪��:c��b�@j���[Y�M@Ai�,�Blã=��f�z�T��-���UF ��ے�"�m~� �b�R�EU���9Ij�d�����:N��+H��ftҟ�_��h�GM"�}t�z���,���Y3�b�{����{�5G��Q�Ks��_7�܂�
T� N���a[m��Y�wϸd�V�9�@3�&�spM��4�Mj%QljEd�}�!I�{��M�%j��F"�@��럋�^u��عAF���pK���EY��D�tp����:&=y��	ŕ��Y�h76�����S6��s��d:�=��`�k�BN��:��5���[���*c�����Wl��`��q�ϗ��B�Cީ�-z��}���x��!q���3*��Ejb0!�6�x���X����f�6iz��İ���8!ռ�c��r[�O�'2�9��ޒ[����oo�Yv!3��AJ
u��*�K^��pe�[}SCڨv��(����.��cS�<���UZ�0�:��ȇȤ�Ϭ�׸�S}�=�;���Ķ���Ԟ����r|uX��8����]8�̍��dJ�5�3�22G�ψ�`B��\?g\5\�K��	M!�Uۍ��X��%-4�ֹ
� i;�8���c��s�E��-�uҕ�H#+|+�@�4��%�&@0�^�&j3�Fܸc�u1��Ǐ�Ç�?��2�J�U��{�&r��{�<�^}.$d�b��JO���F[���7��N|�E��"�k9�||,X��(V]pob�Z�5sDL�%dJW~-��I�̐ؔ.=3G�r��qe�OL�ɋ����A�����2#Ehw� ��������UQQ�J�چ5�w�5~
I����Y�X�������UG�D܎؁�j��6��Ʃ�kI���@��*�z)�p�wnw�	��fA+�Ȧ���������/��~� �� �\V�vpx$@-�����R�������L6�13��u�{]�>O�s�9��4/uhEr�XHo0ར��u����A��`��j�x|���B�i�����u�A�ʎ~��[2G��Nl�w��uLp��&ml(Uڃ�s_%���b6�����3�e��2�'c>~�,�]8c��KŲ���E(�f�߫Q&�(�`���}c?m,���q}��r�#�Lg�����	�T೒��j고u�懇T�Q&4g��Վ�_m�A��sSZ-�Ag0�^(�̀^�\U��c���#D٢�I���`c���6�NXzrrB��΅:�]\ �_h@�x���E!����h ���C�&�d[�5�%�ʛ�f�{���ۓ���9���d5���?��n�믿� )��~��٥tU��L���L��J�����i�`+�	����Zqr鎒x<U~�=���vϣ�����S�����a�oJ�.%l��ȋ�����]�62��d����J��vq��J��l1�Rѝ[", �u�yCo�bc���+�h��L�.�ثpB#�čS��⨬DJ�5{*ė�_6lǛl'/lD�I�[�+�L
#7RJ]��L��*��إqRq�)��N�1�LM�zn�9��M�*>Sվ^�l��e��?���� ~}��+Btr���XT�oi�'KݸP�\���PN/&�����l#�&��4E`qd����W��mK�g��qgKI�=�PP�!1��t�����x19��?��4m�Mljhv��t �:�ؠ���5|��d�?���	kvI��f1ysJ���(�egc�0E�%}���7��LmD��Sv�,�~����P� )K

C%QG7g�hP�t[w�2�����Gj#f�tx.P�a,[�M�Z��6�M��EGF��ߣ����eUGf9�S�C@�Ðm!P0
O���F�q�ʖ��̥���M�F���Oyf$����_ƺ���I�����_�d_��D<��4N�_a5UA��kẺ�Z�D^�� XB��\�MY���#R��p��Ź֠F!ȃ���?j����C M�۬ij��dO�\���XG��5a	�g����^8���}	�A�)��9�<������Z2;��/�ƌi��7d�1��yp�V���݆
�����$��Y��[0�g�!���`�m4��EW���g�2P,�:�V���15�l"�[a���K}�I�ş ��@rT�hyݘ�u��3,��"U��/����j-�d,���*!�Ş�?�5�`I��҂3 ���(�zy�5�u&/��(�Е6�%1*2�aJ�S� J��?��ud�+�;���$(��Z�@�5�/�?����ɱ���̏L��-'+����:h����/溗����M,�
jw���^R��(%�&D����x���<}������t�YB�i�e��!�����QF�t��1տo)HA�
.����Ko�G�a����n�7Őp�l�g�I�/m��G�_f�&:n����_o<]t�Џ20L���
zZ���jU`3P�=�
jr�}��!�
�QV�8�CǦ�<H���X�u����`lo�Ǟ��/\���D�[�� 
���z�;u`��~�� 	{O���6'��JT����!��j1���˴�y������h�0 ?x��t3���f�\�s �Yo�Q���H|Њ�2+3f[�Z�WR738FqR���nH����űܻyW��ڛ�;t�ߺ'O���x:��:���H^{�u�VP��w~*gj�"d�-YMW
�������uw^ ����mD��CP�Q(d���AM�؄ڐf�����.�g �n�Q��S/M�=�tt�Ö��c�Ԁ?è-�=�y!3p��P#�\jР�p�(6�B�t�^�r�u���8y!�/�)�.q<�?d#�-�w:���QX+�r�u�S��+��KS��'X�X����*\ !�HKh�n̅��H�����}<E�E+�����в���h^��}ZV+r�����h�^GfE��k-e$���t����H$2� `�J��O_����k@��t�����y*��=�'ǤO���s}f7n*X;��f9�����E��Rs��^W�q"?��]J5��m
�ܟۦ�����Y�:�s����O�ѣ�&c���(Q�Y]k��{�y���;T���1�w#?za�<u���&��t!!�Xl
]7���:m�n�K����Ȅ�1�^[2Pyt�[
!PD�ĺGo��bAV,_T4�@�TB�7E\����7Q�9x��?�� ֶĞ�p�\,�z!�oNւ%e︜�3M�.�ÜsP�<ԵA�wa��t�:��Jʨ�ky�Y��k�C'q��)�����iΞ�-�r�W�J
��A	��O�}:�|?�#��������J��Fwt���,m���w o� �{T�G���a�E�a�)��Y�Ly�6I*�խefJ��S�G�J4�z����ߍJ3h�ly�Yd?�gϟ��\��n��}��R��Summ�5k�I����~��(\�vl��US�Bm_ڪw~�AM4P*�s�2��a�<h�~�N-�g6Y �$d=}���:�;�� �@[�8q\�{���V�(��jB����#���h{-i+d��J���`�����?+`�op±w��� aGBS�ԅ�X�M���΀�Ii�c�[3Q �|��g!]��9�u�0�n�B��T�ڸ�`[�}�'�B�j���ٙ��uz������˔�_1��&7�@�z]�b���u��;b)N�2�ik�{�����5h;;V�1�-���B�����n�T�}[-�U YMd����&��]R+e�Sƀ��XM%��qc�Y��m�S���i���]{\���/��fm�5�fu��9��<��j7,�.V��=�m��Q9+���=X��e&|W��J8�)$W]�)�2ȋ���hY�aV�2�ƴ2߲�޸vo~�� �����I@����G����%��/s��w�#
i���]:��њb!h��U�e0(�������x"+G@)hv�N�\.��r���\��L�n*t✺x7:����]���{oK/����&��U^�w��niY��N�j >}*��~�����e��=��}Y��t��ԙ^d:�V�������m-fiL�w�؆�����Ջ��d:����ʦ�mt���%-j��Q�� �V����L:��<x����O��=ܖ������ngK���bF�5��1�I�t��ݒ��&�?�G}(Ӌ3�1..&�C����cf	�8��܄��(
�O������m�!K�؆�߹<)�Elꆯn�#���!t�Yx�&e�K�
�P!�Vո���1KR���ڃ�el+C��A/�s
 {~rF����gdF[�r6����#��׾΍�ɳc9WЈh'(�	���6rx�H�t��D%��<d���^��������ӤHd�:�P_w��g�Di
����9���Z2_-���GR�<�����-�\�Pè�f��d;?�5I��g�"����LPBUE�=E��Bç�GX����
��A���|n�l�o��_K��n]���쭙�)d-%&�5ܕ��-���/��7��f����`�#w\K:Q�zj��&o;�{�	N���4��[D���N�#�ѷ�ΦO�3��᱁�B�~���,���בX05��1�C�/���J��L�0 ���.6֐:d�ٚ�^��'����X�m��"���!��t�WQW�|�1rD�HG��H�G���QT�ҲV����{�ơ�7szm!=�����Ƚų��Y����d ��P@h���8����bY�]A���-x���}԰	��g�6N(b��S���|~1%(ƿ�E����`�M�<��2c�T��_�϶��Ε�]�*p�XH�& �U���."�Xz�{���K
�%Tn#�s�r��Ly9���{݆���^��Ȱ�9�4gy�� 
�BB;��EMBV�,k0��
��l˨�������W�����Qe��^���,kW��	��U�_�G
����<��{���Em��~�k[�]����Ne��Y.׺g���)��{U&�b�{�fjĝ?�	A���_ �����
f��$��r�[� "6��-L�T�/����}�_���0��]�
�^PI*�$b���]dj�����1��(<FO����%�]�o U��j��p�����=J_e����5>�)���^��4d��$��V`�%��6��E�Sޑ�HM1�*f�[TJ�b���W���A;�>�x?f�00���zµ���>�`[��v�v��p$��;B��pF/���#C�Ňh"3�܎s�6[��:t#.&��?{�B^\��:R+��Oe�Y�c(�ko����&b��s�A�i+����)�_Hvr!�|�˲�P�
��p�/�������ߒ'�\Cu6��q��i_\șOБZ��M�2��n�A�:Q糩̲��)�����l��Z$4��58�gQ(B�
3p⩒�Q0���T8=� ���i������ݻ��p�-:`Q{�袵�Ё�tӎL�1i���SΕ��H�	��}-�sp]�G�B 6D�������y��&FS4Q����(op&���u���xm- aF��)��W�jQ9���+*��M�M����F�N��x�$2vgԴ�k ���Ao ��{��Ǐ9�Qc�,0�£�]ʤ�&4��vv:}9�9�[;�w�/������K�zQ֑��Al�	�m$�2�~n��C�4Bs�%ۤ�w�%�p�M[��9���ӍMd�@�����$�U��4���7��	)�S�[�4p��'~fJZ,қ�34e�@�`d��ڄ�LF;��>ʲ�v��)x��N���4� ��	
�O�����^����S�4D�8	}
-n|f�3�q��ĉ�����X��hFj0>�o
f�L��ׅ��,�uaB�EU��P�H�)�ԙ��ڴ:���E�,|>d��M��UB�<@P0'���]]�6V�S�^��k_[�������^YT+���{���	F��y��W����x��E)�:F�khR���V0�B����*��H�y�b����dsDYMش��t,CRxT�h�Ą,D�&��B[ȕ�V/K�8i�5�奠�牯�2*B��)��V&��\�܄Wa1��U?�K�鯏B�h����\>� ��z��l;�,k�I�LC�vR�#���� 8й�6�r#k���I�|�H��[z^e�f��g�͚%��31?�{޼��������F/���䰇ː��6��d�y�����d�'��Ez�4Z��p�f����@�K�P���枑q䟻���[�
K� �辨�dFF�8Ǐ�ʂ#˾�bk���w� �����%
�D���B��Nh������Ҋ%Xf�c�wTF�6�wf�,�X�W�!�: ,�թ�"[��3ɬe)��ߤ���,O��M��llm�"���ǯ��� ��G�M�>v�r�S�!~@(m{\���`���xss T���s�dH�r� >��Ύ��>:>� PX�"H���ς����)���P�l�_����g)��75jo���:����)ؖ�����I��:��"n���(��~Bek\�;3v������/v�H/��{C&��2��i���M��E�v2�>����t2���c�t�Ye��D��ɍ���eW/��~�����W�+ߛ��ȢG6I�҆��;����T�^q�%��僖	�����E�c�P�hΓf�k|j�4�;M:e���c��8Q�i�ڛEZ� B��,�8�1�OG��n2@��C�H�j��{���;�\���+�p�N(]����D��;�i����	x67��4>	mU��B�����v�e;D�$����L jԴ��$����(#��.�ac�;!�w�c���z��l��h:�Ҡۓ��
�4[��{���bt�d��N�!ݽsG��N��4R�O[T��?Υ3���٨Ʉ#�{���a�ZTՄ꘯lEu���)��-"���f��7N ��M��,d�_�_@�������U�W\,�5��������0�M�' ��)����dl�z���� 4�9��B !����R@�חz88��EK
�2��#����엿๶�9ۤ	Ϲ���Ê6"���{���73d�[Q�T�`�!49�	t=Q�Mb���P-uASP3QE}Ѣ���e���S|���B�<(2Ȣ�Oq"�vp�۪�B�9S��-Od:����t�C���h�φ7�����7#='  (ڱ�$��6-\h\M�[0���6l�2����� �ƐR��%���X ��zޕ����dw�,f+kY��o�S[�%��K��P7�``�A�B��Ld�Ul���PM�Ǹ�Bڃ@���]�( �6��"�7ZRc³}�1�����{P[�M5�Q���M�r�L�H�#��>�LU2�`x"�&��s��4�g�Q��Rj/�͓���LB'�S�����l�^��i���Ѹs`p��2C!�edD�}XE�!�ML3ۢ�zܕ��J�,��F��m	�8��"C�A�̒�*Ǻזg�9����r�]�t�@�(<����yQ]�7�3��&�cGT:RC����2*��:�$�i��%��L��p�&�>V���~/	/���Ϝ9��C\J��qy�$Z��Z/��Y��st9{ntq|³�̔���<�l j�!j��@ך��3
�ו�3e�G�T�޻e6��+\��F�"=z�:��G)��{4z#��S�g���%�>�Kb�����t4a�Ֆ޸دp�h��z�ȂL�rl+r䄦�B�E).��cd�[Ͷ�ٯF�s��7d/; 6W�������ў��t*��B����-�����Kdo�R~�T���b�����DC� �H�#$��>�$!		��ƬF�eQ���L��z*ɣP/A��J�,<'Œ����i?aQȏ�8���'����?�I��V�"�d~�eOQ��}Mf0�|`O��9c�EQ����4�^�f���Z�����6����u�%X�|~z,CX�'��Kx|ޛЧ�d�|X��1�_�F:���R�Z���:�L��ѱ�(��E=�F���9��9cC3��<Q&��&U9'}��X�D���'cvvwz�Ƌ��o}����nĀ*g�������={������;oQo�%�f��)����A[�J:-��ꀁjy��Od8ͬ5;m�kq�t��Vʙ�"E�U�"m$�rpogْf�O�fƧ�x �p:�k?��'3�����
	���Vsq���Y��T�g}��y(����=�l��?��#���HqlBD�P�|�U-".���#�FwƮھI�A�r��J����?�ͧ}U��/�;2џ�������҅5�Q�>#���+J�}���t����e }�3��nn�`�*Z�IA-j�Z��_=�"�^l,x��Xd�Q����|:�w�G��hcg���dxT�3�!朴zh���e�{�.u��Ԯ��q��6;�[��&@
h���P��FM�P��lhd�|�FF��q���+��p�s��C����/?��c\�g�@)��?�Ġ�|SvZ�'��=���׮Q���3���Fh�E	�,�^w�2c�\K�*LSZ����q������	=)��&����	N�F�-~���V H!I
���G]���9�#��%X�3S�-�рϝ̴/�Qj�y.FQB��:D!:j���Ζ�O'�&)E�-ɍS��
E��g�/�(͍>�77��mK��6z��"��^lhj�_���ʏD�l�Fy%kl����:���M�ӫZ�j�jE�wK�6��lduذ���$�+��Ч��*K�W�uY�CZP��ttE�^���J�Բ��7��74�I(O����RNf@/2H��B[�Miǵ�y震���_�Һ�=���Y���;�2�.��iݼ�ǐY��ԃ�����{�s�9�d�*2W�x}$"u:E�zJ�f�dO-����5�oE҅�K(�b�M�������/�6��4\�؆�b7�>0�u��*xxr�o �i�[�}�-B��;��A�gS9G�2G���,��_�P{��v��B~"�!����g�>S� xVس)��4D�y��l����R6(�"��m��$���x�]�,������yp��V?eP
140�f	[�Z�_|Q�ͦ��{PHO�NE�����}2����HK�"UF��TD�^g���ëv/� [�Y2]�߂��+R�@|U��%ZT�E�O��
m���'�U����2��s�������j��.�j�Z*�5�!q1�_��2�o��{3�����B~@QH��m�.\k=�r�}Vn��_-�� (Ty��j��^�0:	�S����]����z>��	�찐P3��Y��	0(d��p��"Ȇ!ci]�DnчM���8��m>׷_z�����Cz���F޾���GG�߽C/�x�~�{�C�3O��%��{z����AER-57����%��?�Svzr����B����\��1�p"b6pR��+���ױ`'N�h����AA�i�.�����Ќ��K���i�gP���*	��h�����޹�>m�Z��J�&R#���!�08�ġiv2>��#��^���Ds��w��p�
��Ķ��A�k�Q�}ZPT�Du"g�$ef}&�bO(P �W�^��Qx����T�� @"��Z���t\08 u�!U�M��zk�Do��o*�O�S�1V��DhQ3��u���@F�7���&��̣�怮<s]���;�нh:��k�ݒ��+�����p��bvttL��ޢ��)���,����g@�t�-Қ-� �:�\�������Û ~L�ɒz-�kh;�Q�`���~���M�S:>:�[g��j6���ui���(���yF����MZ�{;BWL$#=�5M��'�5B{*T��e�H�.��b ��sH�k{�0���P?�q�V+5v�:W���ӕv�D6�ZA��}�-���@!Y�eQ����"����
~^>�e�[�8!0��Ơ�/�%�hр��Lĉ��Q���� �omR��)t%�V�ڐy\��#"�p��A�"���MgǴ8����7 �mi�r��ƶm�����r0*x�D�lC�����%�5�iC���u5v�U��ǡǖW'�����DĦ�ڈU| �9mP`�ׁ� ���IQ�J3���%0��b E���<c���\�7��IM8�ظrZ͖���
̕�X����q�~��E4"I�E�e�(0Y�`4���-ӕ}/�lKR������
�S��#�(\&�Z��"!�9��$���;dJ#n�Y��ڰZ�
�YvBƆ�|Y.l��r}��',�\�%%���喙�/ہ��/Lb�;�!*�A�fԠPCo���d�`��pj_>O��n<�Li��Nv(Q�>Oj��>h�q�/�)�d�Eam	�2��Odu�$��hH�T��0�"���n�6��f;�n��lb�-���� ^�l���d��BB�mޣ@=<<��`C�������g��%�i��;�C���X��Τ������'}�@����/��dk�)�Z�)�Z^��(4c�!�K��j�]�:�0[-V�O�Y��#�U��u5��B�^�Y��"Ē�Nu�yC�B���u��YP�c��O}W�P�ѝ����:�rNh#z��VT��oJ�~wg��޸.j�'��{�?�_~��gKuxXN&�/Ɣ�Z:��۔B¾�He��Tw��.C��ů����~�ӿ���Mz��Gt�N��N���=7أ�z�u�moR���T��L�qw�4hu�B��7^z\J�jUҡ@3M't��#���� �E=�����m��z6�v���7oޤ�z�N
v�;��a!u>���G0FcM4@e�w��i� #���͞�b:�6��.j||�Ǹ!P��y͜-L��l8�;w>!��_��u�]�8N��hxvN���\�Wq�~�Y(1l/��a�>i%�o�¾�2���E�Q�8}�Vep�Cm�:�����2+�c�XF�񨔳�����uS!ϸ0'�"j�N�g�J�I'��|6��ع�{�g g��[7�����e��t���v�Ƴt��3���4hި���������@��>��fO�����9�` �Q��`V�uNs�ۻ�ܵ4%ӝg�re�����ތz�Wo�B�"�Ġ���gI7o�#Q\�-E�4g��	UWQ΍�6���>z��d&ˍڌq���ÞS�&]o�@�В@B�H��n���-J^z@2r�"A{O�Dd��.����I���,k�m����7�%i�BU߭w`%nAR0)���2@)��䵹�:4�`C?�5[Po�Ҝ<�y���O�Rc�K4�  ��IDAT��.E�Xj1�$����*�KО��)�i�V�u��Ϙ�T��zH�/)a{qz���'��g��-m�lSsg��[Ɋ�񊯿M݌��9�ѓ����hO�[��M)��]��(���6N&��
/9�wv>	&F��T�����?Į��J�Tx���P������BV���yN�	M�Y/
�V'>��:Y�_�J�,�YT_���	$T�R&�^��x���|���s"���hOq��̿�<0�h��œT�+����7��/�Z��V��Y�Ƞ:*BL%`����¦�� /�7Jј�r������^��u{
V<���J�r�5_�p}�J`R�/�j�x�"�	��.X �i���
����G��)����p_����jcph��B9���y���.~S�z�7QI�0V���}�_Tz&��PD������|���K�Kڄ$��`"5�uT�m}v��+`�K�Z�/B��٠��[���-��x�kw��٠f��k��j�(�h���=��'4��$�z�P�C_�B�Ұ�����~�֣�y�M\Ŏ)�E��X�BU��� ]�������g`���TO�����:8��fw����~<vM���h����>-����q@X�����|?ys����r	}Ǔ����W���/��ָ�样��p A�muR}vHg��FRa'����ub����"���	� CD�pN����-��v<����o����ݷޡ��!e3��Ly9N����c�Iz����{Tw��ٱ���ؘ��Aw�٣�z��zԥ���8��L�v�4�^��g����Oӕ�˟�;��﷩����+�Ԭ�2�v�v)��:A��ĳ�0�Z8$ e4���KZ�x<�̲C���X��t���2jgM�z��@c�K��]��tK�X �h��E%;�h"��gt�/�`d>�]�4�� U�$mx�a�tQ-�Ҷ8*3u�F��'�_�6O=@#DE���ћP@U\t��9#d��}�(�+sV.�Ћ˲T��4�Y B�ӝf������	fl�J�-�|wh��6? �c�Y�oR�W�ѕ�+����#�=2�'�g�0]M��o�B�~[����B��ء�
6VvP;҃(����o�`oO
���c~�[�����Y紳�E{�M��N��`�E��gv�_{I6M����p�
UV�J�?�ds\ϤW(��`$y�)����)������I���(�9�6�t��UP-:����f���B�I��M���U#*������|�����{2'����j�!s'�����a�֜��pJ�gl�/��V�S��g�j��P`�u�@�3��f1e�9��3*��-��;���9b-`��F�bԢĦ�)��9;G5��������%E�sj-4�L(f�b���ߤb�C�-�-k�R����o�-L����(##����2�n΀�ѡ�l+x��$
R�6)�L��OT��ʊ�u�š
�`d�U������,	ufP�^n ���s[��(��R�i�l9hR��i�_y4�h��B83)���h��������mG��0�NO�ώ^7nS/���Ɗ��$�����e� "ĽD�q`�=�Є��zu���S a)�0;,k$�2�AzWe�|Q����uG��s�IA�Z{�'8�j�P��Ш��g�}��FQ˒�r����*[�/l���O �_��t.�XW�Wj�>���$�����DB��B=>~�dw.��.ү���*�B���E�+,�)� ��I��P�0��>{�ȬXR�����6m�:�b�m��m���P�}@�:�fG��Q���U[�R�-��kd�\�R�er'��R˲%Rߝ+M�����{﷓Sm9ዲ��Q�B�l-vCڋV3��jׅ{�p�|�u�dTِ�<����y����SgC}�\�.��㼲�.��k�6�c�s��*� �� m���-�ڎO���T��_���"����*�)��X2%�Ղ��B�-]v�Z�X�E'�f�}P��&�.8"5����fLcvj�8��ݤ��/�
v��d����f7�F�iԠw����ɤ�V"��T�d3:a9�Ms���nK�_����Nf#� ��6=��O�����o���������;���������N'�(��ݛB�CT|���/ӫ��6�u=��%�'"�wB�X��`"ʉ{^�!<Y����#�:{%˗�o8��1I%��)�4�>dф �	;�˔�Ev�x
��kF��ȯ]��Cvz��Ҳ�� g�����+���'o�2'e���Q�)dd�U��=PF�H��+@hBAJ��糞eޗb'"�O�Q��,"�k��!���g�HU�3�2<�2�������`����t<�긆:wo���i�өD��'���)��R�^nIS�0m��0$Җe8��i����h97�Dz&���5q�ƙI����ޢ7o�M�<�2�\9�ͫW$s܁�3���7�_��ݣg�o�v�~y�=	�x�sh�r���76e�μn�"&d4>%��Hx��f��>�/�OQ�D+��S��d�C�[fl�6�7�8�D�}���3�Ի:�����ŘH��` 
���g���"{�ZC��!nw�Wu�qd.�V 	���3	Ȩ����J7kP�lE�^WG<�!�kQ�l�ڎ��%Q�6�}�A>?��ل���ZܸA�CG3�imr�85Q�C/A|���J!�ζSkM��&� A����cG��}��}�s( �]�lPv�C����ƒ?�T�}���̄ �єϱb�dP@$�#5�i��r�h4��2�J]D�h �B��[�DVn�-�A*�)DF�$��
���{Y�P�yt:Z�h��4�k�	$�h��k�7�՜?M��mola�|�d�ߢE:U��4�����6�?|��s~&W^z�����'`��s�ߜ���������
S�ٻל*R�Y��F��xp�|�ITE�?�*4���P�Vq�_���ӏSX�T�g�mgS(�u��q	uI������Wt�+PX�e=���[]��]�,>v\�*[����$�	@��}S�g"��g�����H�@�b�3���@�^�wEy�~'���>��F���D-
-&����]C�2׽m���
�����+¾ �I�7��%����u�C�z| Ծ%	�V�G��D�4t:��W���;s�KVg�o�'2E\*}����__�;�g�e�կ����~��خ'���u�K�B����6P;X!k�t�@�e��b���z� ��ka-_��<�2Z���jH�����բ���(�Ţ�n��nd� 
�ja�/���Wt�(c����r*��Ĝ���3���a�,���|��$z& ��9u7[��[P�,#*#�'f"�;�ܬL�	`�1�B�ؔ�jdE$��ӏ�����{l�:����;W鍗�A/��2m����&~����}49����?Џn��&yJ�ɔv��{���������G�I��Cj��ɋ`�4[���2h��>r�5>�G�m��N��D%[���4n�|����h��\i_��SLQ~g&�Uu�p���!��7������.Wg��9g�	�D�cjM�}�t��c]�ٚ���PT*uZW�.H��QT�K�Z�]�c�Y?G�m�g�}a����8�̀jY�:(��\zQl�5���x���@��C�
mR4�FCt�����N�臿�I���:n�9�q5�/��n!MU4(�UfU3(Bƪ��ɹPX ϼ�g�|M�&�H��ZӘ�m�{�����(�9}�����J]I�����։4����&u�ʅ�r��-����of)$��Η���573��N����z��=�C��GP�])�;b�3��	�0t����䈔�\���h��p���EY2���>O���:�F��-ߐ:�|�	�ԙ]
QY�S%��&[Cy��~D^
��j���¢�oU�sR'*5�����������`�W�f�h���m�6�tο��|�%�ۖ�T8S~:���@]���D���!�k�]d�%+����߷E�6��pAێF��h|��2ϳx����~[=Z��4j�5QwJ��j*j�%�a� ����$���n��g3��-�ݕ��?5P�[V�g��gvAH���b��+�1E�f�;8����A��@:��
	�8��Yt]��)Zdt::E�^$L3^S�nv�4�h�Ӣ>��<�9p��y4�Ç���q�F��_���m�I���r�����u;��Q�&H�|M��V:z�����NҺ�=�e./I5�)^�]����O��Or���lT�]�{��#��:��s|� ��=.��]��g\��>�yk��E�x���9�O=�S���M��йTj9�X�d�e������)������v@E	���P/�0���~�V���}�eM�C�*"'�%L;�5LZ��"}��o�Q�%��$VY��T2͍�@O&��Hk��|8gP]xVI�l���Ŧ�@]���ť��%��:�c�
����q_�������r!�%Dks̅0.]�L�3w6��Q�t���e��-�?�����x����r�я0�>]"i/Q�H�˔���{9ެ۽.�T�F4�WEQ�r�p��)�U;��#$�}**z�
4�w �X_-��R4�'�=�#�������ڼbY-�Nv��r8cgc�N�=�G�\��#��bg���C����9�ŭw�_W4�D�����ј���P�Apq:��%�h�i�Q3d;�ޠ�y^�ϗ);�^�t(A[�缘Q�4�A��gr)}^
ˮ�X�3�~c�6I�K��8��;?�k�Om�ƪ�{G����1�lf�,�ᜨ�B\&*Y��]X�0x��Z�����Q~�꼊~t�����?�c��A�^7��:0�Wo���?�M�����\@��kG���
N�J����VpP,����Q:�6�C+�6hm�����37�ν{t>��3]М�g�c3dG��К��|�s���`��(�j{Mujm	�Z[,��2ǘW�N��R�A26��5tw����烺|�;Vr�M�{[[t���ϾM�]FZS,s�ml������M���7���#�oCv�����ӲF�����`ۨ���I�������\�d���20i
��>\�� �	I*��G+������_���=T^��s��`5+r�@�Y��acZw�/���	3*�/Ҿ���z=��^c��Z���m�τ���wi��!n\�E\�b��h
hY ����VO(�s>O2�9y���T���͘Җf	㆓�ZQ�9���(�2ЉD"�V9�Ք�O���X�y�����٤b�Ѵ�s�ߐ>��L!>�IP~�x����z/x���.���+oj�0����j�dkq�0���/�����H��2�β�Z���n�6n�4���r

�8���N<�1�1f���);�<�6�}Q����{tm��|*���V���@����?��ݮ����I6;��_9�o|�d>�'bG�F��(���ſ2'�2�%�әk^Q��[��t����X>	��A%=����D� �~����tk�؜<�%��+��Jav!|ծ�+��]�娍�s�ߔ/y�x�K~�|\]1��T���r2 �z5�5��@�̍�%J��6�a�e�T���|=����&ۀ�����T}���p���ůb2���j�*�g� �6�'(�����;�:nUz���|�6(�"�E��@�ui2�,Wu_�Y�g����L.y<�=1�[W�LajĐ��/��:W ��윾e}�T�֯&��qQ�X�DfHcr�Eh�<'�bW�CP�&���Uҩ�Ї��Q/Y��t�P�DF3�'�!��؏��"�a����A�B+p���@{4Q>h��`{@�?�92��� �. ���!u"��W��֟��x�����m$=��ݎH�ϥO�ҽ�e���I��ЕB�v�@Y�FN4�iE5��(��u�b����-d%1�P�W�a:a'�n�L� �A�."�������ۿC��.gg�Î�!�bҖ���#����X(�Oue68�a��`ŏW�R�"dDUq0�+�i��QK�Fy|�ts�I
�|v�N��шnO�3�� 1
�D� ��:��A��=+���ٙdsQ�% ܞ}h<bA:-7� d�D4�s� ��1m%M:ll��s/Q>]�B+�i�cHOK�)D/��?�?���9�x���L�|��c�/���F(�5�W�͂��s�N�%����B)q=�lG;[�\9���{�c6� &ϟ�(>�7B�d�����eu�����hY�`���jd����
�ʍ^|�\Uh5KΠ4�"��P�:�)ͦZLg��ߐ���~�s��ߔ������rE�gC:>J�o<[���L� b��b�3��?s�B�F�Z�>ڛj��10ʥ�4���ET%:A��)� Qh\gs��#�k&Xd��=;��6�>��qF�b�4�¯���*�a�s�V u~��G(u~�9��Da>��$�r�2��F��@�@Vp�� c`5)��tLӳsJ6��s}�6��ӊ��d�m����yN�V��=����*��Q� *�PȤ㱸2ͨO�NW��b� ��zu,V�@�Kd�<�����H�N�֞��N�@���Va�i[ſF�<���ER�ڌ���kG7´%��3�ҩ�Z"�n���o�z���c���B�G�K7gS	�-`d�����z�6�%�%ָ)��������RH���oQ��<_'��ޅ�D�M�v���6��/��lxDG����4c�8��d x�y�dٞ�"iR�Pq,��=��??��bd�b6�^E�1�s	 ���5�Y��]x���z��O���W�����(�vB��[v����=�<�ɯ�x�5�X\�ٹ�W`]� ���j��Ay����"�F!�����
́DX4qm]'ߔiD�S�V��4��[��촏�f�
e�D��"\Ee���:x��Z���5��W��0*�M �B}��y  _)G�j��>���4zW�cBYB��9Z�X2��]&?7DI���u�kH�Գ`E�����X��s�m�(���Aq=mX\%5����ϭ����,P&��܀&��a iQ�������g���.�$�η'g"/=� J��e+�2@���l��T��'�Fz/����أ��$mvJ����M�4e���۞��[�]���	m ���LfpP�:�����i4��I+�eGa�fA*V��,7���(�{ɕ���|�5��h7%�$*��
��Ð�m��D��4E�L�	@���r"}�<4�D|�{Q�����}���A-K0��X��������p6�E+�N�h�{E
b:Nk(�l��J�g��;�Ҙ|Sd�uE�D�P�
�N� �s.52N$��(� �rT(8Kۉ�Տ�yA ��Ȉ��#�r
p�5nd9o�f�D*�	|dj��uy3����ϯ�����M��*N�ԡMN��Gl�N������W�1���+��PҬ�̅�Z� �PWc�0d�*��l"�6���=D3[��6���<_��I�]$ԼfJD"��H#<�������&��r&�Y�ԲW����$�k��mo��� ���k��n�їP 8}x�#o�GOhr2���o�	z @o������guA�v[��Ɔ�Mh\2�OD`g�E�'�)�Y���m���fO"�=]�n*���~IE�����)�j�ԟ1 L�YƵ��f���C*�Ѣ˹�:�eu[&[���r���,$�'F��H�i�Y�����#�$���j4g�Ք��x{@�F$��%�s�-��\y�lg<�9��>~p�d�<w|�3T
��o�@�&	��#�N�gR#5�hY� ��@��5��|�� �YlS�^SD��^�QԎ��ծ��|����}�l�>��7c��NT�2��X�Ȃ��<���
}d�o	8Ys�R@ ���)������
0�6;��D�D}U�d���n�[|
�=�wR�h���.MO�t��u�w��⍯��hz=���<ݽ{�~��Gw�� ��#�߈��� ����
�VX�e�}�G͹��eB欚#X���W����z(��q�P�@Y�����G����E��Ϫ�S���-l{���䲷�5�yEQο�
�<.��m�eo���>�;i��d�$&L.�N�s�.�\RѬ�̟8>�P��kW��Y.R�/�M#�@D�������<_i}e�b4a�,�*�
#2�錮|\6����S��m���
�b��DS�JP[�I�& *[6�X�f�<��鏵=�I�� ���.�f*k�vUB��Q-��_N��u��Qf����o�e�=�+r�Ϛ^�I1��ٟ�,D�>�s.�,~U��W���,}����KD��@Fa)B.�;9>;����w��ס|5�E�P�av2��D��@%ҽK)�r���Z9�_�[��(d����|��ь4Z�B��I@�З�����3�B��R���1I����c�t6�k�������Ƌߠgwi��{�ӿ���5׾3hv�o�鄍�;����t��w�N�4V� �eZ+1���uV�����0���E�����Q�[P�3�~B�)G�V o^>#+c����Kd��#�օ�^������� �}!��iTBpqJ�e'�����!"z�"�/6�6�İ�&����f^P#�(ʎyRF��
��b��7QELgDMtp�&Tӏ���6hx>���}���¬к�L�xB��']�!��ҙ�n�X�!��g�[�}�]�j�Z��n��z��s�����{���P��@7Њ� ��4I]~���)敃Cz���y-6$ˋ6�N��Ql��KJg`���8��hxJ����N<���H�B����)ktg��"*#�w#6������6;����ܜ&��׋ftci��5�b�Z��_�����{�扷M%����qqH0VZ���gG%2`>_H�^�ס��6��.MQ�ʶ�ی���u��B#�v��f�4�eK�KE�k�I��g�9�E��g��є�_u��f����8�`�yz>$:�I���n�z�[4��{ۅ��@N�,p�e�P�ɨQ��*�& A���HM���|�z�z�B�H���lp�?ST���u��>�;;;+�X��������lk�F�8���>�ɘ��<g �\�w��m��?�r�����3���67��t�<#jC���ui�~��W�4A�W��&�Zw:>���n�����" t��,�K������Xt������Y��S]�G��C��vS����H5���/��"_�ہeQ�M z��5A�����_����_iyN*m�g�����Z���\��'����^Rh��ᱦ$Ï�'���:���y���Un���ʜ� �O	S�y��Z��������>���^����l����	u��r<ò��K�����0��,Q�F�5�Pj�T�X���g�<��K�V\4S��S�mB6P�+�����~���j�U���T	
҃V|E�֕V?n�S����T�ι��i��<�d+���ѴP��L�h��@:��3�w�}H>�O'�FiBw�mE��=dS�ؠD�#q�(8��Py���~dߗ���֧�? M1���H�#��mS�jR
Zg�Nht ������o��鈮~���OD-���t����t���t6h,�2>}^ �<�}^(;,S��F���Dp$r��`�9�Z�����6�j�t�XQ��6H�;�@-�X�X󿃍Mz��s�^d���d���CJ	Ag�E&��(�|�|�(hSHn��6�^��7(h��Ь��F}o��S�w�2�렆2�K�����]�آ^�c��B���N�71����z<ACeUj� :Q�M'�D`�6Q"�A�[�F�lD�}�k�}sj�j�Q].�`�ˊ�Oa��&=�_Pkʛ�d1���^��^�&]�ٗ앬'�~꽨���K�p���l9��n�r��(�ȈM]��ep�Bi��(��-5��׷�h>�Q*��
���6Ns�J����� �$�J�f�Ȣ�Q����-��t��ZS}�����y�!%W-��M������D�b�u�k]cl� 0ԠE�����:��4�x�
�Z��4hm��̈́Пࠬ��2wZیy�9�@�P�;��Y��Z��'�b�Y�
jZ��A�uT���܂Z�x�~N�ql;O�ҫ��6dA)(�n��h.��a��g�ՌKUƬ� NavA�~��,�&��P����C9͕����=u�q-���'8Z+��YI�@�a�E�DC�W(˹:krϼn�����$ڷ,|jNE!���pF-�����/���t|�����[�·�������|<�b�hпJ�ЃG�R_�gߔ eC�X
n�W�Lk���jC
����0y�y�;4���ʹ/����c$5�5��ąZ��%$W����[��l�P\o;��3p_���&�	�߇M	���ML��TOt�.�eu��qa|��_��2�����ˆ�U�ǭ��Uα���ڋ>�!��5Y�j�@�_��]��V��RցDLC;���k6O�����݉H@��yl�QU#�_d*�k�L�Y 3��i4ʌ`��K-t�6Z�H�x�}��������6��5^TTm�TA4���F���{����c>��Po��0O/�r�\�l����g+��l��Bw��Y��Z����n��+�؛�����e��h!����L�F1�L�.�h��J��g����9���i��F�_9ۙ(<� �U%�t���k��
v# � �����k�����xb��2tH�JϷ��D�iU����樷+R6f�=�ߥ��w�}���P�������o����GD������w�q[���.M=��#�4:��e��E�vE�T��lJ�u��X���(�>����Qmc)ZD勡0���FC���'�Oú\��E�;��u��Fq#2Q'J���dN4�u�@�}���+�gE����§dyNAB���C�R�۲1aGY��_JH��/�p��<��B��$k�\�!ĿL��4�.����4B&[�4��Ȋ��h_lF��EV=���M違��b�.�G�*�p�:��Ծz1����Ճ+�ܦ4�NE$	G�Ք�̚�#�����|����Db�BB��+��L�5��G'�P�l
-��N9�~^x�E���Y7;mo����񡑬�7o�Q�Eh����F+mul{Ц�;4ss����ظt:|���ktx%�*݅�t�QN3%��U�CZ˹��!2�6���lS�ǯ��D�,Ҁy�A���P(�-�5���^ԋ�i_1C�2ݱW**��Mߤ�^��'5,�n�hI>�)9��2 ��%�л����4p��,���(�g񿍥��4.$�;���QQ�h�V�rȢ�5p�U�W����$�A"�NZ���tc��"�>Ҭ{�LUT&Qx�V�
'P���sUэ�����MPi�ꀠ������>��JuM�V6D����mt6h�`��|�l_'�b���.Q�����mXD�^B-H���/��%Mg#q$��DR�)m��&����#�a�e�?b��
;@�-��NE��E�w���������=�r�� "BTQ��P�"�UMYT?�J�<WՈ;lޗ���;�%��D�j���*O����^vl{�O�g��k/Í����N��쾷x�Ӷ@b#�W\��A�,�}6�"ʹ���r�82 i>���A�#:��"v!��u" z-ʄn"�g�ꡨ�Ό� ,*����x�P?S�_QT���gca{����З���^�G��f<)���܃%z:����6CqU�H:?��L�z�y�a
ċJ->WA�`��U��>��ީ��K��ɲ��3܅��7��ʔ@�m�	���=0�qHF%�Mܸ��Ҝ��q���z���ݷ���RcХ&65�͡�v�zh�^H[胎Baj��XZ���!���-G��"
�[�
�ɩۄ�����Dʻ��n;ԣ���օ.N�Vaiy͢z���~��O��>���y�=��O~B�ٌ�n�^{�u������4��ӏ~��ƫ���o���֥n'B�5�hB�i�cP��M���.����0��f8�)�F��J�/�v��
��Ӈt2F��B�S���LJV�WjkT͏�[����4�n���z�^�h/�I�S�hK�@H�WF�ϭ�f���q�1 b茞���I�b����r,;���(IoA� �Qi�Ű�����N
�$Vּ��h� �nJ�*HPks���9A��($�F���ٷn����_/!��S�	�s���]�J�)_�bE���@������v>q�::�8���P�8�Lhc0)��𜿆���%�C�O�y�:�� hl�:tes�^�ƫt��J�-Y�p�*�b2`��˻�1�^(�Bݴ�*,Z��?1�s'k9ڿ�O�W����#ɰ	��]�s�a�9�-�开���Ј�G��jc<Ճz������S�ֶ�h����N�b�f�CZ�>��IJ��W����L�mu���@���8���9�t��%JU����H�q�xQ'�q?_Rʀo���HB��63��Fٔ5��Ճ��E��_3��I��ߌqŽK>ҍ:7uOQ�[����zs`���T(Қg2���:��T��9m��v ��h!s9��r�������<����*�_mL!�[���6#�nN������)�㌶�;�[�)�=x�k;���]���u�A)P
�(pTf�"�'��*�����q<t��D$K^hk��hXƤj�)�t�����)IZ��o0}�P�2.m��	�����)@%g`0��ڿr<aw�H#-g�PC?�)���)n��% хy�l�5x��};��.dW���>�0
8Nk����C�<P&��-�Ót���(���:0�`�����{���c(�@��&%����ބ 'IaJ�V����v9�;�3�D!AfY'�U Gi0�Ő�^ɶXh��@o���6�����7w|�28����e�С�D|Oܲ�6&��W���r�-WҚ���T�}����Rwڠ�s�u� ��KP���z$������eJ��?�E?� �DB}M���K�(��w���n��mv�洳9�M��'�xDBq*x�L��a?����źB��S�#!��1���W��j�G�}Q{�Q�>�y�7p��L1bX�lɶ����:Oes��ߤv����+��|E�\�?����Ճ�%8N��7t��]12_��t��]v�w�?������G��[o����J�bp׮����5���#�(�i��0 *�Ln�~���m����(
���9?�V�=��p"Y�׳&�;]qvÊ�m����|�D���rjG�P?���&�a�IcGn��T�b�@S(��eO��_�cЀ�_�����,9$_(������j�p�p��|iu�*\��	m*0�̴��:/I}Va4H��Ks �3�,�U�1QEcU����Lr�L�Cj��B3c"�]X����|���{�ͦҒ��F�trJwO���*ֺΘ�[��H�� ��4���f�Ц���?��yd�00��s�7D �z��U�����1��s�)Ͳ%M�s��QC7M���7ʈ����+@~��ƙi���	U��_�2mmf�(�n_ߥ��f�̴y�5��]*�cW�N�Z�@s��.AH͏,��`�b�9�S9wQ'���
jJ����cDj2�jmn��`��k�k��Jp�M�i�R���mqBM)�5�Χ�vۼ؛�l�J-ھ�"�t�se���� Ƽ��&N��[0��Ӧb���Vہ��BF��mQ��v��5U�@�ؼ����Z	yB�`��-�f�c� PՕݰ^)Қ��Zu�c+�3��G��@da���,�d�eN������&���V��B��}���	�������c��ϳtJ��sͶ��m�s8���V�kc���%�c�u1�= ���`Z��c͖�~�@�
vօɉ�0~F{��r�֨YڇM�?Ff�B��UY��u�\�@��u�;+f����]i ,�q
B\P/�@�[�'Ou����5�\��ԏ�`Z���*���2�+���jM�`��E�](ޖY�LQХ�'�OW�l^�_i��HZc���tl� ��_C��
�D��U�f���$>)t�Xl\\��Z�Q��%����
(�U�Jl�k���5�Q�,_K��v\y޵@M��:
N3�Q�B�B����*:텽�>����T�\)����V/T�,��QU��z�,��L����*C��9����G��䈦�1-؟�N&��g�kWh�v��Po�a�)�?�a㤬)4w{�T�1i:��^��)0����*�����2%𲡍�(87�ڒ�;wn�B���Yt�tF<Y@Cko����Cz4��ə���4�`�roQ`{��l��k�r�:�3���������m]hQB�;�	�ow�w_�-z�[��dв� ���k�A�����n����ߦ��-ڂ��ل26����ߧ%;ۣ���%���hȠ��?�)��=��rA��MJ�1L'sQ�
P�Jy��_u��\��Д�8�BI~�y�����H7��_x��Թ����8��b��	n�$�I���+ͬA��Xο��3}z6G�w�%v-��l�Mh٦%h��Ig����MZ�3��d����<j:��Rۀ�-G���#mv��.��
*��͡,�������5ӂ�w��,�j+jMsRڨ�Y"��Bi)������,�l�QP RZ�V���F�׍	N2h�Ȕ��:[*�S ��j����F>�zi�%�s���S(�b��}����!���쌝�-����@�	5@Ȋ�02���ܢ�Ȱ��+�!0���2"����u�<K��ޅ�.no���u�l�x=����p<�n�pKj�Nf�2�Q���{u8M!�G�uPo��[�z}����(�z0�f4d�M.�:H�2F�g��a9��1S2_P� ּ�� [�ǰH�d�{�޸�P>s�m{F�`���dLM^#+�g3(��|�9</77e'���������\�[��ڤ	_ۄ����?�f�A���"2���m7
�M4������@���¿�>,-H�����V�(l[���P��@� ��s�Nq/�:���=6�� M�1`b�ˀL�Nz������{6xnM�'�dʋt!�Q�H��X*�Ӂ��!<��/�@q!TQ�l1��d�C����;ԅ��Y���m"n�8�������aK�7}m8�;qu�VWM%%O%�о�:d�m�&T&YDo4�H�7.�	eU��S�	߇�~��.ۯt8����$>�z]��r���,���j�5�J�sF7������W�ښ��v"8�s�o��)�U-��1۷Bz3K ��y��1���Ҍ��x��#�3���p�f	�ʽH3����p-�+���DЍ"dqN�|+1	��J���Y��ˤCm����[ ����q�#��0�L�)Bv�Л�T~E������2+_^�zY.��GՇRБ� �r�b�Ω���qC��Rs�$%	��Tc�촭�����ْZ�u�w��e� ��m��|M�r�@�th��g�=��lBS�K�>:������>s��?�]�v@�~G�f�:�-�c�[�����_FZ����*�����[��L�oq}����U�]iK��Iv�����(z3�&;�-v������U~��x���wo��{����)=ZLi)Quv���� ���g��L2+̵v�1�2 e;R�*PdY��HHԋq�6�@�c���Jd?��+�=O�f��7R��A�ԏ�3z�[��ݠ����^z��uT�f쑵�wM���^�\�;�[4��>����>;��>s�nDcvR&1��{��ty�f��,vd��3/6*��� 倩�e%ܱf��h��xiF@^a��H�P"WB��8Dx�lKvn�.�yL�QS2�0�	_����ZKdH�h��e�/�e�5\Cj����`HMf�C_��\{��>��M���)/�WS���acr�ߏ�:]�k#i	��Y(ETS�
���]�"o�95��5���,W��ȳɘ���&hgp���L�7��dA�k����6�X�EZz��~F ,��P�.hײ��ꈊ��TA/H1Pр���|Fm<G�@7�(n0�CPf�`�����k����6�gS��T�7����ӽ��o}@��䟟Oٙ��QV�:���tL(��g���P ��9p&�ё�6҆4M~}���ۣgv��ʀ���j>����FOj~���[T��>a�J2��J�s���`���AZ��mdQ� ^C@�I^)w��6��Ti��/�v��c����y�N�O��5��Ad/���)5���Z~�85^�ΰ�"��\�Qk%�
�\;�$�(x�A���v�F�B��q��	mt�ʅbC����Ȝ�$A�!�(�hd�0>l��0D�*0�
sR��j+d[����|��&��¿����(j��|K���:`a�kY@oY>�8�?���ۆ�Պ�A����u�Js�s쵨]4h��(eg2��;��B�x�Ŷ��s�ՠ�����G�Gt>�(��>��ΡP�c*������h�9�	JB��c�1p��مe���`a!sl�9��o�e+ph��o�BO!SR�F)��RFD6Dd�FKg�P��������A��2����O�B�>�rf�bB��YF�h=��vm��`p{�N$JŒ�@L.�\��:Or����y��=*H����� D0�sQ����{�lI��)�W�%�x_�↰A�f��A�DB��kg
�B�w�
J�I��1x�hy�p�b�º�
�U4"U�I�C- �>3�+�7(,�F�yW��������}%�n����
���q���i�7\[�b6�Q
��_�{��V�ފzklL��$�@M��u�F�ܱ��C]e ��s������<���_�B�.P���i�f����PO�ޠ>����������E��#����m�~��<[2z��b|��������,ؕ����w���#���z������ID�PP����J懨�k ˑ�qȭ����4C�i%�v�X����e��N�3mG��Ie��2w�mT L�9�]^�)]�ߥ���x�MD�m�7����N�'�~�O߾�5z��5���>����torNg>�BS���ёbi|Z�r��/�Q�p��7 �B�҈���g���;�����ّ��3�Ģ�I��٢�dF��I��AOp�_Cf�	gg���{}(S����G��[7i��/@t�6�x1,Eğ씿��oң6h�9���:��N��5�:{I!F���5�6J!N��E�k��K��_U5-��iS\��%�4����h!��=o�&uy����7��ޡ �
��>��x&j�����q�
(��)x��c�x4�Y���yN�'Ԕ@��\�2㽂B����2��JPv����!-�L#��V���]z���`���|�?��}��Xi�+>�8���1)~B]\J	?�Xp�}t�H�*�r��P2�7:��Z&4�Ȣ&b�eoT*6�s�Ɲu�8dA�ܨ}�h�2�P-x!��Ѝ�$j���lm���L�|�v�C[�������ߐqo�X�z]�� 6���g�x�Nn?�z!٨�n?�Ǜ�1�y�mG��N?��Z`�@Q�ˡ^I7J����B`�����gi�c1�u����4>�5l�����s��P�ۣs�9��,��B9�JE7I�^F��Hc��V�B���Q�e�T�h��)�W"&���W�{E�����7��߃��A�E�#�8ϥ�Y�m���*U��e;a#��S^� �NQ��Ji+�JK�q��yFMLaK�WI`$�qo@�8S�?i��cԐyK����H�B#��/|LڧJDxsr\%��a��Ϡ�_�B�i��ɹZ�{F\�[�6\'Y����f�Ć��-��	�MKi @�4{�b4a?
���M�����u��<�z���8��i����Ì�~!�`:���pH3�Љ;r��Y���!�^<y���e�6g�
K�K��:6BOWj ����^Yp$V����8WA�TR�h�JGJ�^�$j ͫ2���\�y��e>�k/f+?�(Q
����k���.i��
4䐹-]~�������w�h�v��`3r���0�������5�^
� �IF:'�0
��ꀷ���c�C�(@{)�/��R�y�h��6�3hj<���wm2�k�^� 8�
��kڼ�9��a�� 2���b���̆K����t����N��A���+���Xԫ%��T�����/R_+rU`+<�O2� 	�)Gӹ��@M5�P�)�}���^G�}�uV�C- �վ+ ��q�X�:F��%m~�ѫx5�gߕL^��Z02x������l��O�yu$Ȫv���#:����1���h���b���nݦ�hB�����a�ϟ�ZW+��S�ӹ+�p�6d�ִ6 !��ly��W�e��c�?�����;_m�P���0�������D�ߣ�N���6�q��@;��t�|���no@���-z�����	�!���p��=q�W"��ʂ��8$�sf�I�L1���F-����N�}�U���O�Mlm8�<�_���is�NO�e����=R�t���%_2� �V�z��_s:��>;�vn���( ����F#�����	�)Ft�yX���� �	��u+"�8-0��m�M���7D�Ņ��v.��X�{���Y�b�Q��F�p��ȳ/3(2t���no�!�۷?0�M���Aiԩ�WV��<�l�/�*#����~;cy�`��q�xC[2��ΚoP��(j�dWV�9y~j�
��U����8v���S1�l�-�B���y ��G�Ґv.4�@vGj����z�:]e`�rw@	��9���掤/!�?7�R�T�C�i�T�#�pZK��jٰ��Rd;�j�����3��9��<_Le�VCJ�\�X<v� �?ap��������#�z�&<��v��<�2�{����tD��ÇC��}������h7������������Pc� ��Ct��^� �M�6���� \D&0% �j;��o18m1�����������f�"�랑��h��j4�A���j
n�8��Y�G�J�(J�㜚
���G���X#6vTh��	�,�+��i��l��9ۂ�t�ƭ!�Qseǅ��+�Z�U
���f�bZ�$7�>?�6�%ۏ�%MǙ �x�n?�|8&��S���m}Q�\]8{�-�f��f��j[�i����u;(sFj�I4V����x)��D�0��a���P^W:X7�أ9
Qdj�u۫ߔ�Л#YE�Jg#4��C3hy�)�:{>����Ul��@=�;P���E�b��!Et3�w�h��~ok@q�C���s���YfIE� �K�\U�u��?*�"r	�ΡY^��l��@Z��)
�.�F�t`(Ǣ�R|ʍFX=#ւs{�0s&<#�8
�&�P�5U ����;=�HpZJP�C��ґ�����{����a����Mgu��)��.k4�/��m�~�sPv�DC��	�\*�J���V�s&%]4B}J� �=M�.V�]���~�O�lH�K3˲�mOXL�F�t�ڳtp�:5yOx��[�:��9g{�k���Ϭ��#�c�4��2�J���{�PxK���Wk�C�,Q��Dp�͇�	�<!*���/��P�ol���U �|/Aam>�P�[�Ǐ�t���;�����^���bՉ��<�/w�F=	>常6�y�����P��,S�&���2��dN��ܧ�!={�k��s�2���g��ڑ��=p6P=KZ���0����`��A׮?+������{@�������S:a?b6��d2�^~���^P7R�:"S���I�C5 XU@*y�_;>�~�G@f�{��>DlÏ����{o�$Y�\���b_r�̬�����g� 8C��(�L��G����4��D-Fh� E�`�����k_r���#�&?��}�����f@���ɬ̈�{�_?�Ǐ��eҽ-u��VKƊ���H��L�h ��%�hKS�hp�i6׍/it%�K}�L~r~�U���@I��buD#'�tC($2;��uZ�?`����.��Ξ<ll* �Hc��l�1����)���k3g�%8�v��Ԭ�:�X T͌��j$�Y��ѴTG��jX��ܕF�-዇�ӿ���nA�CP��h�BPz��:�ꄫ�/K�:&�sD�8d��|H���YX���z^��f��t"&�9��_�Ϡ�i�{���h1��/�B7P'!V�D���U�gE�e�z����'k\��=�S0r��#�tP��bz�:��5�
�\M�[P�<�g0S ?:�lz.mD���̧29�ʫ�3	fKiV�d�1F�lJ."����)G��&h��Z"�H��>�N���a��o�?��ߐ���?}�yrv,#�5�]�c_��uC�qOx#㉨,�$��k���!r�#��ME��7��.�����)@���F1Up�����I�����&�B�`5]�^O�wv���-�P�vp&7w���{����
d��+P�u�̇sy�󯷱!�۷X�
a��>;��E3d���ǜY�/b�H�F.����;2� �e� �5��� � ����D����&дĊ���~S�]P/GT�r+����S��s����4c/bS��`�)�rk�� a�����B�ϩ��5]��5d��V��;��&�L���	Y2
Y����#?XZ��TLs�o���T�0o���	�L��6iA�9�����R)T��T(:�QZ�,�`:����q�.X�\��J���F˪/�����GbY�X��\VB߇�tY� ZsJ��5�R�̸�b�
ez}�)K7�^U�ӡp���]��vG�ܩ���T�ى����l���!��������K�)�u}6�f!]�D����z ����\[��	��{k�YE��jC\����r��^d�F��j �4� �'p}���r�5��{�9�l��M�[qP���%@�5.=�$��C��O����
���s�@#���5h
�Ea`2�eM��
;�"<���i�2��s���|�"�����!"��
!�{��ץ J���H�?GjG��&![�� �,Wp�
Ū�d�[������*�]�(�BAl�d-ʉԛy���5Z���P��Grr:�,���\��[�^v+��԰���,X�
C�7
����U�#�s6���2`�,�M�
��>�\NǓ�����"��j���F�8���\���xe���R��jw��6֍���
���8W���\VJ�W/a��|V��������@nO��g껧�+\��B����HFgci�:rk�4kmc1D��h�a�?�կ�XF�������ݓ��\�ݥ1���ܽ���ݑW���'rx�J�^ʉ�b�2�9���ߗͭ��+�� ,&��i�\G��}��M�2w(����~����r���D���#*�:Ġ�Lu���`�sy18Q#ђ������F����@6u��ڗ��X:e��%�%"�C�xF;֥;]�"ح5	�--z
Y��~5���ۼ!�qK"5<}}�FX�̟�;�M�֍;Қ�Q�,d�lWd*v���%�}��e�vDl�����b7��%'��$�u�w�w$:{%'�Et:
�'.c+���9�mnɶ�cdz�3��LG�5џS��{�*��eLC���v�,��T�I����s�85���,�����X]�޶��i� ���:�v�j�JS�]�PPՖtt��^�$� �E���G��2I��)�DϢ@��z�Ϣn�W�e�v�/��C��!��%w�C��LF��{\}�
��Dh`���u�8�aet]Ss7�A���Pn�"%�n�ے�k���R�2@skAs0Z��IA3���
�WZmڬ$EZ	"F�3���^;��8?��P����4���`%jgu�K�iΌ�|:c�t4�_N<&,ξw�my��{����j$;}R0����2������r�w�D���L�<��^���\f�l�+�D`Чp��(2^��D��I�`o�0��J�2KX���f�(p��ҵ?��1N���u��H�Z:��
�˚0���#�V��;���5����_m�`1?+�!?���x�nWpu�3xW�U/&���f���`��q�&�ZB���	1�2�Eꡲ
w��v�l�]����fb5~�˄P��32��$ԭ�D �k*SF�㸉�Ρ)�$V;��+'�-�:E�Mm��G���-�u�����V�6�|+���6�:�3kl��zK�z�zH�{�r����Z]�! bk�aY!	X_fN�3�>�X	A\n�RE�e�0ٕ�n,Kma�-��<��$���x�ko�4(��Y,�2R{���AT'hF��P���Hؽx �K;^�\�L���~Lb�s���ȹT�U�tL��c�?ye>������{>3QF��]�1׻�B`69X���2|K�+�l_U�{�"���*߫�#��|�ܾ��K�_j��!lm(�8S30�.�����c��F��K�����XB���?�<WQ�,�J�rY�g����W߬Q�,�TA�~�r��^��*$�MI'N��<�I���$���g֭CB�"p��Nu�4K�-�T��i���­�K ����*i�磸g�".k�׮�4�1.�!^�K]T�*�R��e�|��}���W��U�]�Χb��Z~����>�s��U���=ĳ:���:@�<9>����Od>�KG���޾�=It���+�'t���������\�����G�O�w������r�qLo�ޒ~oC^���^	V�h6�'�>aP��[�՞ߤ)m�{���6�4F���n�@��l���><o�MGYMn���J�F�D4�r��q`�@B�"],(P����O�ޭ;�CmQ�FdK����ݕ�,�tr�NF�������dL��:D-�Jy�w仿���Rg���M���鹺�
���*��d#BCm�b��ݔ[m%�?��;����lA`�:�W�^�P��e:�)����28;��8�M
���4G���c�io_��[
vZ2A��f)�}}[���ֆ|��[r I ���L����Tɘ�=  ;E�TfU��t��Q
8&%�� �su~ƣ!�"����t�Q�D�s2��E쁶UoK��\z
N>П/��h"M1	YG�L"X�b�F�Ef�m����C%��2�����d�՞)hk5M1s6S@(W`�Bo�B��ޭ����M�s����Uiaizg�c�$G�M]��q�/VE(��Q��R�Z��NK���7$n5t\r�7�̜Qy�U�1� �=sS^��#�{��ޢ���4߷F�@���~�����)��3�>°ʴX�#����f��N[?_Ǫӕ��=i6ڤf��ύV���u��w����eksS_ےz�&[�4�^(�EV/Bq�L�g�4=|�����JΗL�-������2���
 �`:���=�K��6���$��lN�swW�}뾤���B��i�wdAyH�S )���T�%bR1M$��|f��������M�.SX������8xHL��R]��*���![��t�f0�-���Q#�R �4C�T"m�23!1���&� v�	$���F��@�w�p5�.+�y�y���بB^/W!�����d�v1��;�|z�F�%K�KR�t��W`"�ڵ�pɌ{[7c0/��Ηs�)HJ��>�" ��Zi(�f�f{j�(�����g*,*_1�\��k8ƽ�T��f�2�U1����f���*.@�Z`'��AK�E3�y<�1�|a��	�}����f�Q��?A�
Ԋ0g��"�����@?�c�Tt�u]�k q�a����� #t*���փo��*R>���e��#p���ƍl*��X9�Eၠˮ~����=3%�����H�Kq�,�>����zvpm��um�ܽ�4�{9Q1CG�H"cs�����>��!��+�������y5[��ya%!!�`�8)(��=:�,( ���5ρ����6��8W��
��o�z�X��E�Z���Y��(�s��|GF���Y�D���*��{ �rTf�M���`��&���|D�Qe�\Lg��5[�z��(���p�u��^�+4P��]�kt�^]uտ豪� ��~�`��y��C9?9W�~]�'�7n���M���7}~v�$���J/�K������U	�?�҅%"����>�;o�W�ٕ��5�>} ��<����V�-qW�c�X8x�أ>#��}|�o�u+�W�����x���U�.Xɻ��)B����B'�P,�ӸP�T��	a��|@G0؉�����:xw7nH�ڲS}_6��B�$P�+����yo�|���!�:�V�V��$�@��!kv>������,R�K�c�PG���M�f�+�{�1�����))
UN̺�����Q��	�`������<hl
�~-�$���٠���R�t>�l<W@<#$Ζ��㖴6�4���:ԅ��� ����!Ȃ� u�沐xo[�޺-���t����L!�g�������ň@����ޖ\w�1����E�BdD��S#�<��y���Y�s>���A�k��ѷ�-S8�:Έ܃K�*^6L�?Y�/h��s�W�,���s�B��D|�����L�q��jaSn��;���~������o}M>����vo�xq!GG�-�;7��N��?��_]Ƚ�}M:��������3�I�������ݗl>�_=�	Գ��"îc��� ���n9��-&:�r2����T�v����������("�T/�qvz*-�4��/�=���9���w$8m��/��[��cSfN��"�	^fPPP��s��$�Z&|�Ps�r�mu�����t���q��sމ�Qȉ��q\���cÎM!sF�X�%���z�Q�T��~,t"X���WE�8d����Ӑ���wQ��ZP�⢞4*M�6	�P R`Jh�
�Y�&4�晫�PG�E�c'�Dillv��kQ�(ت��:> ���t�@JnWa5A�`T7�&7�b�S i�v���D&��p�Qψ��5�۝�e���S�X�Y����g�~	{�Cnb4Ij���$����̝L���4l�:�k��7�uޥs�V��U;��J���kC��a�a���-ٲ�q+6g�p���P�h)�؛���-��uu[H���PXm�5{�� ��c�NPF|�[�ϗu���ei��^U�X���Qߊ����;�} �j��.lbN�P��3�?�7Μ��N,�`Ni���D����0�W��|�Kc�E}�_�L��@�����������Ȓ�
�%E�[/�����	���9�/�W��ೊ6`�z��l���ڡm��l3�Lm���BjᲥ�n����@�&���#�Ԁ�P�a�����d�7b		U���u�;�E.� T�2Ѭ�t {O��c���̢]?j=���
��ܹ�J���"���е�(W}W#'�V��
���hmD��q}��������E���ѩ�|q��`]�7���%{7�u�e��k�֠}��Jtnb_�
2|��tF���IVK9w�@+���� ��A,���������>y���T�=zNa�_S�	���Q���D���)]6�����{�5w�J��ï�Q�������DBE�mE�g�2�N���c]�5u!�q�!uJ���+
��<��ZK6�my>��^��FLM������|���ZA�c+tE��E��^�R���)y��aҹ��������<�G'��c.�eb=�P��}�
p��jl��4$Q�TMd�f�c��H�7�>�^���8gw8��+B�
J�c1��͇C�S�D���Miv������hm��۷���+��N���
 B6�ܨ7dc��rc8��|��[
TP���{���&�>�̍�`aNf���Nm]��!+� .d�+�:�R��ϡ@�<�P�$t
�"ֻGHQ��)q��	���7��k�e��꽗~%�"�ҝ��vg�J�Q�#�S��/6���-9|�B�� ��틳����S�,���M�?��ߒFҒ?��?��W��oɖ�+2�5��O�>���ҕ���u �����cnΩjj5����0��5A�L���'r��H:��޻�����x�t�u��hA���3������}O>z�9��&`QX@��ѹ��m��:�8G tm@髧�gX�d�NIFV� ��g�s�\�D����/�,�3��jnn�A��aR�32t�QoP�퍍�]MA�!U�1�U0(y_X�#I�üptfF�"�J���qƬ3J��Pͤ��0[�ld����� �n0EZ�v�Mf(	�@E��e--P�����D�n����D�+�&x5<�md�}-*�ee��SX�ux�,t#��� @D[���Df�\�08=צFiQ�43^��8��c	���F�tZ(Q�.��#9Ab �O���iE���Iqt�U0�Vf`�ҵ���W� �y~�qrY':���Hz��>�j炦~��%�VǉI�O���j��vݣ�ڒ�Dm�s`���zm�;:��u��]���| �¨�f�-�m�YﮊTҭn��|��_����|���AW�r%(/��kW�v"�{�M@#��bEeu ��ѮY;�\�M�U����w��<�����:�:Y�����W��-�hhL�ȕH��`���ym���x���˖	vu�����ܔ;����\���d�v��^������^�kaRX+	�M��i<�*�t(�ի����y-�"�Jx)��1��
\V��X�������.����x�@�8RQ�s岶�D�ρ��w>�C�"���Ӥ9���Ok��2fېxA>�ʭÏ�'�h5��̖R\*w������Lt���+̿F��������D`T���Sy�ѧ�����~F�ӗ��}騽]L}��'�jw�(h�J	c[sm9�\]��FO�Զ��5�f�M���р�}��3����f�z�/OC9:9����r���ϡ!1�!���-�z�=t����1��z����Ʈ��kt���MϝhImz=8��t�������SK����:��D�L
u��SNd��Z)�|FI[(���hy!g�@���?�����.��k��g�'
�������囷���F���Y��zH'`���O�H�ۓ��9?8�;7v�x�����:��+xZ"��Lh��G:��)��q�.�l� �:X�R����?�^�K
_�6jdcXh����R��I"�fM���k�hln�P���\;���mi�ۤi�Ը.��K5�'G��ek��%�Z]N����� 0-Il5~ET�Ɣ�N_͌axe��+���A��YJymg	V?O��+�HM����?VkTJ�r�%��j�W�� r��˖����������-�on�o�w�����;���\�@"�;��<�Y��Aj��x8��s����_˃�у�rv~*��7d[����:�?��c��'G�Q��q�����fD�Q�%/�N��������Lґ�cѓ��Q.Aovtg ��Mз��<~�5��^=��qh=$��x�;��44p)��R� ���u��L����L��4uM5�m9��l6�P7�X�g��#����|N���9d`P\F����-wN'�TR5d����zS�#���7��wR����Vn���+��Ԡ%3�)�'�IY-��V�TQ�4S�h��9�5t�q�Hm�@4Y�����[]��͒Tϭ��9�x�Tus�Y:d'K�H�i �L��/��K1Q �>_�	�p)�zF�(�iάE�~��`'t}H��6�.)#�A��h�9�(�\�\�Ͷ���N#���k�Lzl�Yn�9�8#��Ѻ\�K��R�����5[J��W93�|P(4Jh ��NA�6�|4bm0�Nl�`��hS�p�
�:ǁB>h{D`X�1E�Uv�/���z���P��.��s��Y�g�)(\��Ί�X��"�ul�ڋ.}TQ]�YY}���ĥT��Qz��^��[9��:��Ky4Z{j��_�*�Y�Vcf���]8WAa�v�L@�w��9b?sC�~\�@���a]�����I�Ts��1�����hJ�\{N��*��q��JU�� ���}Pb�H��`�ח����7e�@���֐OƧ28?��|,�N���j�s+���E`p�yA���~�cS2��f�}�4��J �I��`!�<1u��HU���K�"qa�!�z��lp�K�,[`�j��|}�w�L�,� ��_�.hN�ـz��l!��ޑ� ��.�%��5�%3]Uh��l�*)����~��C�9.&g���3����ؒ����z����ֺZ�nGb:�,���%M�={E2J���M��(��c��f�-�˾���.��2�Md>C@��4;M�ygW�o���VV!��������+��J+���������A�?�M��Wj��qI���OKO�-�1Y|��d�mr#�!��f��A@.D�E�w����d�Bh��ꄾ��	2@,D���BqbJ�%�Jl�N&���(��R���u
�r<ɉ�]P�l!a�!a����z���`�ו�w�ݓ�3��������rxv$�R?�դ��ͧ�F�l��`4���PƑ:v�����EV�1/�v�/������빧���搇�r��Aa1cс�:T���YS �W� �;�B�ۗ��t6�%j��ӡ��R�d:� ����ޮ:��X��`-w쾦���T:-�&X�؋��"���j���&c[�}�^Tms�/#�y�Q�����/{pc�|�l:��n4�Z�E�<8>!$�O�	�²k���=]:n��D�^ʦLPh�o���|�9����;��p���9Ǣ�?��fP�8T\ ���Cc�Q	\�ˣG�_k�V�K����?��Ӑ�5�>B�6��������y~z����1�S��NXLb�D�d�v/.F2���O�z���؈�n,��-3\�,#�f6Z�Ay.�M��#���HҀA/eo����^��3̅�����M�&J�P��)A0�0��o�/K�d>4 B'"�l��sT�b��	M Hr�hR�;17 B~ �!��cS__/M�!5C�R���U.-�0�0�@꿠����<�F��2PG3k���5�\�f��?�!�z(ĉB��J�Mz2��( ��7` a0V�H��te�si�{@D [�7�1B[���^^>�F�Wj��)i]�y#� O"eՇ�����a}Ki�� 2X�65EY	%�������s�Q���!ql:[��'-mSG&36>��T�S�E���`ne��D������M�u�7�%[�Fr̼RěM�u��Y�/�@\E��6+�+��g�;)���0µ:MY���B&>S����]&��)����pY��
��
��C�ip���|9q�H]�ш�8���y�㳉 "���@��;p�r���f��3��I��\�l/	�.]�z�2���S�3��ѕ�[K�/:��6��ڳ�X�����g���P,_;d�
 ��4�7e��m�&tnܐ�ђ�/e8��pЕA�-G�G�<x�vi ��q�61cCcE�E��)��HDk���C_�L�fY:�3��`�bw��tڼe5M�9�⾻�:����VK��Fq�q]	l����x+|�Z��@���3������z��������#�S_�����t���Eɗ9�}�uJ,Y4���糹���ɋg�I��m����]��IS�g}�l&�V�(����ln���J��V�%��H�:�7,(=�}�r����.��To˝��ꗟ�D���������������p^��(	��T�.�x�d��A|�ك�jP���Q�Y3�9՘ �%�Qc4T��ƒcuN�\LF��u���(����#�45�j,�������QRcĜ��8Gl5e�i0g��\���B�����[��a���P���'aO�����(�������ѝ�uv?��S5t5y��ߗ��o�`8���ocs��	�]k�u������X������#9��:��:'맠�t���8@ k�\��9ӿ!��C$D�iC�2"�^4j���$@@d:����G�ӟ|���P�L����`p.�sONu<`DS��g������d���Ai�~rM�-�<���ьʚste_Y��aae�F��mП�g�5R�]�9P�(�Mp⮓��<��	��y�����3�i6�FfZ����looS�c :��G����y��}�m���j�vI=��N�n�h%!���[��������������ā g�D���@]� ��ց�n6���6�#�:�X���K�ay�y�	Ai��̚�E��FÑ^��o�:ݳ\2�YۨsFGc�\Lu��`#���TFs�˩�6j�郂���>�}�S��ǈxh*q>��F��&�!�jr����tu�ԇk3a  6ȹ�����qEzyd"B��dh{�E��z���ph�$����@���X��[q]78���,��C��,�Z¹�E2�躟�̤��%�V�,b��
(P����ʞ:�jG:;}������¥�:7fN$Ao`v6��~_?/��GeAZ/"��}E�^�Q�� {�5�h�঎�ܼ�EF����(hKX�˨�8�o"��@�j~���P��ѽ�Kk�g�}��-�Uf�Ք"S��`�V�+r�yJ*>�SA/Bd��AkȖۅ��v�p�<N�8�|�ɜ*����0��>� �w2\xl��sY��i�e0[�	�d��Nl��x���e�õ���TH�Ă�����/�8�%`���Wvւ6AҢ
�I��+2�_e�}�«�Z}��8��{�jtb/.�����2{�=�t�q<Y:�+d�:C��o~���<����`)ݬ�d�tq�2�3�tic+]�`]���yf����UP}�+Vۥ{be���"e�6���/���d�D �t�G2V�0�����D�˱��"{*3��_
V�����^K��M���r�r���O�4���u�xD�}����_�\
�m'gl`��S
�z��9e�պy���U�i�7Y�D<�J�j�8M�J��$j���k��W��}�~��u���]�ses.�A�=pk(��\�g�OS����^G_v6w����A��~Eͬ������J�d���P(���R���C�� ַ�z K���*��������[���O�)88;>S�x��cv�t��^���З!]K}S��\���zӔ��Z踸����F9;;#z��NdC� a�aܲ��NS��8!��BTc54SuBQx����>'M��j�~�h
lR�T�鐱7
���F�L>}�X���R���tjߦ�M�����m��ޭ��7��ё��/������=�!ʏZC(lB9�ݓ�nS�';���@~<�t.�l�veh��)l� �YL�}!�A�ʁ����|��*0l�����z���H���P>�DAǄ�xgwG��ݓ������W/e	!��o�{���Z!���ޒb�,b�Z!zp	#�֜ڄr��x�xR�=qW����y�<��3T�s��-����W_�gm�/tYl@��i\�WM����B��\(�{���ܽ)=�b4�����ߕ�ϟ�@�t� �6��\��{Kvvv������ɧ�>��-������-�I�eI�C���6�fҴz�����n)M��4�Y�`ƢC��	��0s�#;7���o��=yp�Ҥ�A���歮�y��}P�E�C��zF�./R6�E׍e���j+�F����P+��Ů��:�v&�7��9?S����
�1S�	�H�c`��R��/D5 ����]��p�mL^ݷ����<\��ҵ�++�q�UP��rc�))�+j*��w�*��+G�$�
6�{��oX��f1��?.	�
��2km"����^o�F�yЪI1���El�N4��|���"�6"�(�etQ�7=�KmГ�ߒ���79�A���eg���F���PW][�3��X?��9���� ���w>7�jG�K*
�?���z��5z�(�׭L��s�&Y�/k�������"��Ș������ )�k%��.�	m���RI��&�^|hO�u،�h��FfA�� �S�^pX0v!��	SU�ҕ���樮�	ל�2��϶Uu>����.�Ķ]=\W�T�l�d����B �+V��%��;��{[��U��`�5�}x\͜�ȥ�LA0g�t'\�Z�L��Kn�����,���^��BY�V_���N�W��~��ը��V�7�/�#W`�rS4��]�bu�ҧ���_�����=�zSb�PB�J�
TO�'����𸔳a �㔎>2}����<��}S���k2.
����n#b�<�d���ݳ��%���޵��M&3֟�]}��:�r�xK���,w���u���P�͕0��T�{�&�f��
���;ڤ����*_��:m�N��I���A���ޖ��B���*ڹf��g:V���A��f���Ci�|��!H�	��	���N���'`�"p�ą1;�LX�?YЅ��/m!S������^G����Ǝ���}��'2�_�x4V�}$�����=�ҩº/��BG�Ƴ~گ�,������7��՛�0�U�	c��63@_���]�L� ��BjΧcy>��t$n�!��4p���DY �~�����!/�0���9���JPG}�l�:��F�����䎑�A�"������ar���J�֒�]�5y������Od2��qJ�j�;�ޖwP���KWd7L��@��[J�
���%��I�J��2B���Ԙ5�3�������due��:�[�l���x5��r|rD0�k��+89�HO�x�dЩ_�Q�F������F�BoDl̩��pM�9�y�6$pF�Ϧ�/�҉E�h�k�s�/{/U����3�޿\����Ñeo�%w�l����V��"�����Ne� �x�)#�K0:�����D��x!3u������eaS����ol�e<������z�L^)���'?T�����P�����@�?�������'&Ϭ�5�:��D��-i��չ��b��f����,�������{;rSͿ�����2��oEV�ۦ>�����5�d0g�ł��U����o&�ܛXo�[��d��&�oo����D�n��q9�P	� �w�1 ���� �0���>+ȡ+߆N��k�H����[�y/nNBL:�g��3��~
���щIr�Ku>'��͚�A�թ���1�Z�?�<!�+��+=�H�����3���u�-���K�Md����� N�!c8�3ZX���u؋BZ�-:7��1�k�@.O�lK�۔�f_�6�Ҏx��� \<c�ݨgz�KŤz?�D��x�V2qT���:f-�˵ii�wxJ
��^�`�5������U�=̰�(]����jw�jqW/��B쬀��] ��U�D.�1�]���������L�?��B�m��1�`�o�3iyEq�E�/q�k��	���DN��z����lo7HSZ�T$an�N���Y��UR�g��h��(ho��r����w�D.g��/S����ҹ��i��㠪�]���~�ZY�-����<�~�Q
<�v4�K������r�K�#;��5�5�����S��Q�_����lŀ[���W��.t�˘̓�lN����4�yq/aoj���kY#{�	{���O0pn�bm�?�|Ĭ�d�;d��Hc5!x����d��$̦�YaL�X � I�x0?倳˿����`�/=	,���*�uDF�7߃�?���B�>:eun�;V�*��$�2�$��k�]�n�ˣǏyb����4#���e�@!�����P����e2��D��H#���|pn-=B�9��f��:GP+9���,+�]�n)r�F��$3��'���_���c�>�m88Ȧ�}ң�lT����V��D~�֕,�Z��W�0����P�N��W/� 'Pm�M�����)�a��d��:S3���s���@N�TXU��E?C�B�z�i}��l�7������۱S�ӿ�O�g�@���M�ލ[���{�޽we�Ǝ����\~|�R'��)��M�.^� =��z�~G�M���Ey$����Oȷ~�7�.�wnߖ~��l�D?{�_��#B�Ѕ�ڨ0�[�ҡ�ٮ�2�X��Rׅ�k���q>����IJ�-uH!�g�ڭ��#9Q 8�g���K6�<��>)Y��h��oc+�O>��@ ��Qh�0��7`�E����j<y�l�*�h�e���A>c�]w6��=����=�J��,��Y���\_=�5�s޵ӣ@=c?�������ͷ�ޑ�: �KGm�+�;::e��=˙�A���Mz�sJ[P�҅<~��i��Cd������<���}��c��7������Jh�6����&Xp�c���h ?O�=�V�Ȩ?$=�VC���u����VP�ѣy��F���^\��@|����*���tN�l�s�(M�Y\�����PC�FQ\�,㎂��B�ۨ'���
ՙ�X׭�9
�	������3��n-$J�!a?)�t�~�*Wd2��WǄ�T�B#qn��>s�Ŋ\��u�lO`g��j�p��X�RƧs��[E�\Q�O�Jڔ��w�.���uhH�>}�E�aB�
�&:�:����>�d�-�k0��jlܜ�֗��- $�d��&8'Q]�g;�r�.��ǉn�uq�>��������� �s�l�Q�5uu���dԧz�a��&�`
�D��W�{M���S[�ۭ���Lt��꠱G�z�5������O����/	�8Y��!s  t򲊴��b�d�sF�	tP@]H����O�n����6�zS�7NO�O?�W�GAs�L�a3P��쪋 d���MD���7�b���7(��Ҍ,��@��̺R�94��iӲ0��,[T4T>��}p]G�Z�]+�]�+�йG��f�`v�r����>�^�Y�(�`�TP+�멲�"{�����=����Ҳ��ٱ���*3�����+�� �M\�4��f����
�A�0��p5�[ʪ���
͋�o[p�������&�r<�ZC�K�W����@���|$�F������k��2#��v�5�7��O�A�(ͯ	B�Mk��fK��Y&�yf"Z�˔���!�:�5��\P�5�oc�F��:J(�t�{o�����'G��PHٷR��XTkY�
ȹ���`�5O9p����>��U%"�Ct�`�~��P�����?2�}�����z}6�J$�"藎7�1\��Ҟ�>��˫��x�^�G����3��#�iI����u����<�
B�MH>��bLߠ���;2�H\ ��@�'�ba\"k!2����|@��Ǐ�15QY���Q����	�f7�#M�� Y���<p8���#u$�:H�ަ"�.��������,�ITX�/8�h�=ן&���T�&�5,�qOlaB0 dK��x����?�P�}�]i��������}$�z[~�ߖ�;{�@�����h|~dt���:��T�� a�0������׿!�) ��I�����ܻ_�
���Uc����4ÐAR�:���N�F�I9�Wc�.i�4��8��/BQ��T��g�	l5�5�Ej�U�T [���}�q�.��p$�G�N6�����/8U�_H�A\]-�_4��+�i5��lL �rQ����
��Ϳ
Hs
���V0O�݉ �Q��E��}�ʪ��@��E�.�\:>�����w%y��(4oLԂY_�/���d�
���i��\Τծ������fg�}�j�u�/�5邟g���#�;/�P�/��M���x�s	%��X�����@>��ǲMH�,��Z���Թb��O��b�`d�o�>��W:��=5kNOհ�e�]���j:���%�Z#pm#���o���_���<]����%�hu��e5��UZ�����.+�Cs�K״׽�G_/�4��h�\k�h3Z�p�l^^�sسG�#(v�Ae���kH��qz*� xvv!�+=�8������f�4xv�#�-�y��M,i8�s�-�(u�Mi* \곛�3ڐ��,Q(�m� ���ot>��O��v�%p�'
�uM��X��,���4Ci��(��֡>���2��A���hʞ����B��R�/Zl$
C�[|�kP�%�l��f,�V���i1wX6�v@ʞ��T�p��0���^�}���6}��D�s�Hzy�2� �#��(,t������<<�P��Ⱦ���;RKޕ�^S>}�R��� ϬS��:o2>+���GeW&��%���,�� �1Z2��g��a��~���ދ�t�L���H�P���gU�\�����1�,��i��Z��G/?3��Wk�Cq�ټ�6�*ps �J�OD����m$�@X�ʊ�J׊���Z�4�G'6����3DV���
(y����:\���g����[-��c���� �+��ҕ��6$G���u�j�g���� ���VA�Y��D��b7�� Va-Skz1R`(��{�O'��S�B@�(]"ˏdD���k�0�:�"�����mKG���F��q�.�������z����#x_��T�b�4}6o5r�>���Fk/\;|;�m�{�:a.�e�]�$�{���<x����z��)���]ޏpW�X���.\�Rߒƿ֟'2������'���u��HF�]p�vk���������qtY�]������>!��ݗ����'u��7�-h�lOŚ�w��<����mI��l�w��Ł���we�ͥ�]{'*�l���rBT�&z�O�n�!����x�4�����N9hd ������D�Z<�.~d�5���~_0kCe�X��C9��e�V
�1̠���~h�^o2R��t;���H>=z%����Gr���P�ђ��O~������}���� ����P>|��<:xA�T�����ДV8eN�>��Nrl���=���@�����=i���r��-�<��9wD6�FT}� e%�:+��6�'[�p:�DTe��O�Fp�@�wԹ7�'��KMH���Cͺ����g�F��������ݷߖ���>4O?������Q�\�W�	�G��,�&�ƲQ~!�w�P�7Q��U�;�L���\5W���AV���{	�@�d�(��d����M�	�=(��̄�C���˯�U��ߗ����4�^9�+�)@"`���fИu8Pygg��z�A�g�(HbF#(�(8
�KtC�����X�A��5f����ڛ�h���B�}�f˹ձ:5@J�����Q��7wpz&��-n��S�z�u�j-S������>D���C��?AvKqf5\yd4�T�|܄�fKZ}'�B6n��x9emb����;*8ͼ�M�6���[I�+�!�!S�8X��F�Z;���πsk��.(�c�9ON���:�Fj����6ډ��-�N�E�sy�s��TgF�oƖ��	�b}V� �
"�j�DEW�#I�K�
��[]	;�	M����	Pk<���P�t�K���{j�nt$��::�z�z3��f�vHW�d:���Bm�H'Y*a�.m��V�.���8���
PK}�r<c]1t�z���t��y� (G��yLǓ�Ǚ^�:a���,m���U4���Js}a�;LY���^�x�$u�+����(�70fSHPȊ��&S�����G�9��b��M��8���l��fm9=V�<C[��`$���Vʺ9���/dQ����hy���Ԩ�Ȕ�ѠW����<����K�2�`�+����}���?�Ս{�j�X����_ߒ&��:��?�װg�A�դښ��@E֜Y��,����Z˲P�,%��g���D޼/|�5����v���/�	���,�u�d`_y���Lן��<��W�Xp�����t^P\��wd��o���L��R���@�0A�.w|l���A0�u1�u��S����5W5��ڬ����`�����Tm�-�F�-)����#P��E*}��,c����,f}�*'#����lIokSZ��4�7E<�Pp��^7J����O9/�a���X�e�8_�)t��* �U�D��Yn�J�Ƃ��m���S
�`�w���4�Eg7Bۧ 	\}�3Ε�VP!��'{�J�ԃ��.����`�/���n��Pv#�3�l����<��]����%k���Am:�N��n�^��'����,G�br.�û��k`�7�#t>�`�G�-�.��{�L� ӕ�ƥ�0�x�^��/�(˟�0]��X����*�����>���K��a���߻��<�r�g�9��T'@�ƣh5��d �z.O'g�2����� �u:)IM��$A�u�fp���r �������ߒ��n�!�J4	���W����'?���w]'�Y�C>��M*('"���<X���jS�z�������ɏ~,�Z"��L�7�E�*�.�I�&��I`c�Q
9�]6˜�P�ɬ�%���K�/u!��g�]�8A�ġڊkC�}�\ȓ������*n[[��p1B����f���EjM�ڞUy��M�oԟ������� �h�Ms0Jo�|&ҽ7p����Ēkn  ���]g4Y�	+��Z��՞Fj�x�3�[�_aO�b���y��'E�bT�4�ձ�{,�
Yp��~��0���Ou�M'�@��?�ٷ�"|�;Ԯ� ���Ȥq����J"z�8���"�>�9xQ1j	�uxt�ߙ�ZɾL�<��0� �\|�_��t�s��s�*%{6匪a>c�Pɯ�)3O�� �<��O^�!�5�0�͘�I�&��^�Qc��e<��VG^���,l�e5f�O�ΑCO+n��
B�r��qS�d+�j���I�Kd�+[ QX&/������Vܔ��)i�[��`+�O$iD�sgO���{�BW��P��Q�C��b��P���
�d�	x�>����$�����ݓ��������0f'sYO����%���:��:����;�1��V�+�DFN-�^C4C����/�+��kF��k�|�T[����ભn��D6��M ���'�X��A�+��h��ﵹ�T������3����Q��Q8׶/�>�:U�R.}���%{�3�ݬ,:Hߦ�� �dr�{I��{Q[?c��MIu�NW�+�Im��j�ɋ�:)(ض$b����_���܎�Ц[�;
ڈ�~c:������G3�*��k�M5��A 2u�~릈�iX0�����
���UÿfWc�Xf�'�|���kH\���"R���g+�f䘛�:*��ʟ�{���Y������C{��Xߦ����P�Ҏ`m.�����nɬ~E{h ��� �C��cҴ���g�|]6���Ig<������߬�s(Gg��b>��Kd����K���������P��+h X�ɐ���,��:ޱx���3�u�E�9�H:8���|K��;� �'H�aϢ �p_�!T��@����$·b&-D]�\"�s��%�,�2*�P?����t�g�����ze��V{2Q�2��R{\�,3�P3�N	�]��G�!k��+o�3�F .�n>՝;w����L����RB���o�`�q��.�?�L��Z���v���_�:���̃�P��FM�?��	��`�PVV�V�!b��������5��g�������������!�ϼd���܏�5�/?wd�������?�h��s8.5�r�XԺHf��.!��|��F��4[y�䉌ԙD����]��O����N.�"[�B'I�`$��ciT��`��!�f�ߦ�}���"�QX!>k�,�~jLj�&�����:��X�
0�s3#�D2�.�Z��w�ɏ��rr�R��z_����r=�fS�������P�E2���kX���pи�f���S]؉>��j\�|C޿��d�T<x(��7n�ObC���!��z����}7�y~�����;�xn��@u�q�(�~�Vs��̻M�Rl�S�\n'��kC��� D K�	1�Ԁ����zlb���8\Pe+p-��z�9
'�'��N����Jw~���B�S?��HZ1wշ'��J*�l�u*����)�מ����^3
�ϒ:� �xPZ���ԁ�ט%4XA�f���=�S@Q�ؔ�@g\&fh�\�jH��N���K���[�,��e�;<t�1�6w�uN��d<��4jM12e��m��T7�i�1�s��6ԟ 2kVo���<��fT�%DmF��עK��uj��B�m��ƨy��)�i&Y�j�T|+�e|ز��=�~@��.ܽ����9)*����993�e鲡3A�x�K&�eIr	[�$�����I\Ld�|���c��V�j;���)�]x�Js�s�d&�3	�sR�þ��]IQ!Z
�����tN��j13kN�"��s'ow�0����}�7Y�Bf�����#�D��K�"���+�@b��6�c�*�)�Ѧ����,k��2��B��`>	3��=���-�=[��Z/}���q3��ڜ��Gk�"_v�P�ĺJ)}7:[�l�S�6�P�Ś��
�r�j+�Y̚N� �ь���y��=���}�|Dq.���;OQU��f�!_�6)e�룰�QA}�<�60L��t�j5{�߅a�W&�Q5zw�Q�5W�"�ṵjM��]�9�+8o��退�`����ז-��{��}���������-M��kN��S�Y�����O��}'a��b�Θ�@U�ah5�����y0��\�_��Y7�z�rlW�	BO��+��2�ׇѡ�`��V	w�?�\.	<m�$�)S�<�L�/t_�m�[�&��~螑����l�e��Xe=��G'/er�B��Dm����[�n�(D��'] �@V*��@P����I�8�_��
z+T�gs�(���7lBQ1���3	�d���@@�x��l��xoC��w�F��	Ľ����5�_�uo�k~x�3s��6x�|f(���?�����r�涴;m�y)��3��I�GwA��`��E����.�j������� �\��k��Kp.�GA�J��ɿ��&��},���v�t��^���w���(������)8���Vb�k2�?�^w}��ݟ��u��7G���s����E���èK~�.4,�W�G2�˟���OR,�NKPM��\�Ώ���T����H溨G���54{�F����FM�:��X��	�ɼ�=e��η�[oߗ�Ζ��BNGg28KG���|�;�%��򡜼xl�1�^D���)0C1�:6#u��|�ც�H���g�D��?��!�b,O~�|.G�����t7:қnI�U[�S�C�c��?jy|\��� t<UEv����rq6��s9?:�N���X�ӻ�孷� �C:��t�̧���w4�6*%A��IBt��/q���."�)Ym4+���� Pa�#V�F*ii!Aa�)>��ѱ��?��%0�'=�l��@E�n,���B��������HK��e�W9��NYI���<�:N�.������1{j��Ck�g�gT�������p=�`���,��7��L���s� �LFj�x�����錭
�%�2e�Ւ���_8��,Nt3�t#u���W����ܓ�D�v�"���_������5��z[��1i�%Z+ �9_�f� �9`'�^��^��wZ5�N`����i	j(<��t�ʂ�@^+�!ww��)k̚��6L����I!���,Pa D�6���#�US��SPz��f2��
:lu�C',3]H�פ�u�N�r�vW7�nS����!�q���@y6R���D����xC��:�9���L���e[�jΠ���q��)bW0�ֹPϙ�CF{����(t��0J�i�L�Ĕ�i_��#2�П#4�Wp-
,c�]�s�&���2Z
�ߠ4���m�Y�_0��P0�l��S@��bJ�Nu�/�YL�PD��B[Z�X���P ��K	����-�:p}�y62le�����Q�YG����Z�0k���F���g4E�S�ٟ�;�NM�zm�EH�l��^��J��#iӎBF=�] mA�vVT�u��ˮU}�<?9�5*�IeFm��{�\A`�@�
����y�b�F̮2��1�K���,us� �P,����H�9'� OL	��`l%�hfid O%,�9ʪy������^��x����mXg�Ѯݕ� Y�)��r2+%���!�ڤ�郍]�I���a&�猀0�q���j��C���~o�Uv��U��9��.�:@��#eK��u(�F2�`M{X�}ѵ+��zjqU
6��A(��~���\B�T@/����(G���pM����G���(1�5�~���S7���E�R�V�,��}f���N�L�E��9�ԞQ�Y}�D(h�QeV^z��օw)�ZٿJz�-i1<B��t�cM=|��>!�3�����	#�Z@{]�&��9�����������>�~my��2��*�ע�6J��O8O�u�[����;
�-�SG�fi곭E���fG�$��YȜ�p���_�@d����/[�P\u�?_�X��Z$�kե���� ;��Ba��?��/�N�K�іBw�� ]�\��T��XW��^~������ �c
}XAi��r[ӿ��&�����3��٩����Ï~B
��z�krgw_vo��8�ɋ�#9O�̮,@섓Y�d���@�3u�څl66��*����Tgv$�jM�w���) ���tp,G�Db�7ը%hN^���*6�(=�EZȆ�=�t�7t��1�������B�^9���-NN��E ��z>db����s��{6�E� (�b��G���ն��Xeu`L0�k[eU�8)�-���t��?�w���{������C�t�*i�hgB@��Y7b^��lv�"dWIΐ����E��a���t�sʨ;h�5]hT��={%���28?��Կu�m�Cw��r�#̠tZJ�"��|f���}��	�K�t P���b���3�7���W'Grv10uR}?�/�h���޶�vt�-R;z�癁���5X��������?�|2���K�n
mT��fa=D����%3���6l�A��n2��k��t�X��c�(�c�Q��̄f(�}pwVs�����e� HU@�G:���+!��P���T4
�Ʌ�mC�W������X��9U�|��^��@��B0�qT�x����ׂv8{:���e�Ӓ�,�Q����c�7JI[jz
� TњV(�FB��b�-m��A���4�CDH������6��^eK[;��AZ24c
���LJf=��#7UW��:'���5m�A���6%t�Po��+�<&�չM�wG���h�V�f�k�ʪ�<�J,��AsMf.���?,s�).��Z`t4p������g
��R���]��]�\��1`X�S3	.
k7��+�i5�h+}0�߂�t��i���X�(U�$�\�l�FNe�N��IdhYoy�؝�G�-H��v�"��*�׹9q�� 0;8�9��q�_t> A�Y�A�!��� uTƫG��H��aVN:Ǚc�0�f`ղ�Bz�.[���c���&���e�V�W�xӞ����:�gK�yoi��	��0�*j\��_�7��g��3G-nCnݼ)���KYߡ`��zk�JP���A�//Wt���
ʎ�d�MX����A�G��B+�/��Nl�ԔF�]eK�B֩�fsi6,�ɗqO�)�kj0�/����4V����l�hu�>ڦǺ�M�.4�<E���;��@����,WU����f��bU�C!�TH>h_�y��iݰco� ������b���߻��c�X��+��a���~��-��O��O=��m�C��d��B�g���M�o�p��A>@b�
%}E�2�$��O���̏��j؎ed��J���3� ��E@@QDF*_a8��-����
R�2�@�v�]�y�������EC����ɑ j���ΌS$�o��?���ɳ��H����՟��ᙺ���������+�ݯ}[�z�����P7]���C�棨)D�=Le\�cCj���v_F��P6�hڐ�B]I���j1�#u�u�oݾ#�g�r88a�6*ʪ�("�p�al��:} ���TD���LFCY��}AT�ߓ^�k�8���F�6�M"�qZ3Vg,5P�4 �����N*���5i�&`=��y�
`�����;2{̒��¡��=M4���H�dՓ���	�X�dF�]V���x �tb3�;@���W�՜^3��s�JYW6Pw�u݀�~���RF�9�`��$�j4��:����w�ٔ�FO�|M��[��������u��ː�_�����o���񿱵�l�����@ >����M���[Π����4�H�N�[��W8�u=*U�Y�E��3��?�PZ:��޸!�����\;S;��	�@�P5A�'�$T~3��j�	,X 
P�} %\���)�21�h�X'ޏ�o@g4JmA'""���V�xVaX�0Ω
Q����'�maXj�8�	�Ux2j�,c�2TL1/�ҽ�!Ѯ��nCj��t�+>�I9ʤ�ПG�,���6�]����-�;�sGƝL��T}#�up��ެɒ�8�w��UU��Ku�� � HI��f4fc2�4��^���1Ioz�d6���$����d�$�8�@�$�D��5z��ʪ�3�~#����OD��F/��M ٙu�f܈��������b���Z���o��a�{��nQQ���j�eT���=+`��U���#]�{
j��)D'�O�
Qq��`������Ȯ��ް�<���P촀��͂�-�/[�&�ȶ��IC�a�"�X�Fs�
�c�e ��r���2�<KD�-X@3攨�R�Of�������D�2��[g��b����3^D�Vepʨ4�>��n��N�D�ƨ�i[~"m��h�Ժ#�
!�߹) c/h�.���j2����KM�LQ�����Y����E#��J�ԁY�aFRCCQr�g��E�6�Ͳ7�Lqk(���x��k�ٰ���_|&k�ن�?�R������ecb<K�5��-��m6��H�VV+��9��%�� ����!�X:D�4��r��*@���? ^/^��	PEm=����ww���a�#��hN�!���K�^o�����:�T���J��[��3���H��K&�m��3��ON�M���Kk@�E�Haq�����N쿵�S�ҥq��w�l\\ϲ�	d�����2���&�[ϽpW&����H�AS_wVV=_S��c�eO}�2��}2�=��'���>�ӽtb/���^���öi$bOA�ɨF��$MT}�1k�Qւ�@��,m[��ƈ��hkWU�+���M���i���O]mW`��?x�5 ��.tFeA���A�Quuj^��� �Ȭ�5��Rs(Hb�A:�wz�և,�a@�!!�:W����z"�������<:9�w>�i חЭ�xv,�/O�a9�G�ȃ���a9�e�+�YB�-J��w5��s����LO( �+y�/���c@�岵5��}y{v.sutG[�lw�։>T�4�;Vp����I^�|�z���W��N 2�L�( Rߐ�5[���1��R��P��ju��Ņ�o�:/���3���[�FK
4�|v��x����|b_�2}�pQt�2L<�"�^�`Cpz)�zo0V�4q3f��\&JhQXK��u�A}B! �a�'�YWj}��+G0�`%ڼ#��2�T�����
V�w�|�U�
I��Rz
��' �c8��/U67l=]��d&ݲ�2,����i�^����������Ku��l�#�5�p� 3��������/�̵���{�����������o˃���wޖǇ���
�f��
P	?Y]*�,���tk���h(�ܾ-/ݺ-6��Bfz��H7����|�;��$xnQwB(�v�m�����Qӕ��y���h��"�xZ���1R������biY��W>O��Ǭ�?�УW���p����{[KXZ�����5Nt���0o��~�BB�p*��\�˕.J�ڮK�u�k��~{��+�:C_+�Á=c���B4/zN��W@��Z 'H�g|��f��O�tp�����b})=����􀍵Ffc��h�ӥ�kp ��<m���BV�dM�
*�q���ϊ���G�K(C�iL#:��Z��&<e�M��qL���4h2�@�g�U���r�!Y��Y���<Q;:�k�E��G���y��O�+�޷�oE�9ΘC��j_p*ea�#ʐ���=#d}~-�h٢�TLR�
��6^U�r휉��T,�V7�]�P;�u�QԴ`|�_���)����x��s�,�'@;o���>
i�|�MW1��:��@!Qg�F/�zl?����h'63K�[|�~<([�'����MH�Y�Oq�*�vmm�>��})�e�d��g�=��rS��\(J���<h��cf��Nn��4莥�RA�3[ �:�Pz�o���kK��1���ZJ��jQ��5E쬾1�S��۫���L�Ǐ�����_>�=�X�''2]�)6a�*�җ6r9k�Ҕ3$j�D�^�V<��4�� �7ف��|��_�U��7�J?�H�K����g�c��UkP����>V9 f��6��	���e���y�Q[rxx�_�r��M�C���¾���^X�"�/�#�:�*�N�5��olMq[��JgN�N�<�6)�)�*�m��l�sm�!������ߏ�(���d�}�[��Jȃw,�9` �_胆h�z�'U����<��F�+����st�j�8Y0W1�?	��;?����%��`���3���N� ��x��P~t��5R �s}��r-�g'r�@pqv)��Z��sC��\�P^�ҿ���>���/  /K5��p���k{��W�H-/�r��HV�3�V#5�Y6�����芜td ~ ��r+l���3�&`{W�̬kҿb" 3D����X�x��ڮmo[�=�5g�"�P�0����&׏L�GK�:M��z�eu�7&O�`6��bF��;��HQ2~9�GJZeƬ�S4O�yM�.�X7��]JVt��0�E��0x�
U�r�"i}1di8�1�������y�q����2��]F1lj1 ��7�����������������.&��5Xtv(*5�ൕt�Q38��ɑn2:_ �G�����$��Zߩ�s�ԍ��Yaՠ^��|2g�J[0�h[�����7 �����۷n�믿���)���:�jڌP�A��
L��z��M��ޑ'zO�-�Z��m�[�>��Q��T�2��nŐ��N+j沪�c��n�y�h�O�����3��7�z�=hSzM���t�1F�թ�E��ܳ�yʎ%:�����Vu�#���ﰑ{�v"Ù�����KG�nss�`sYmD�;Rpؗ�gk���m�� c���&�u�	�3��ё���3��G�:d-o�jMZ�Y��Xh�2R&ŏ���z�Vi9�K��ibH���T�YGwHc��;x&�W�0�l���')�%1��[$7�=�oը��O3�W��F\�s�B�X����^Χ�&����b^���J�_������Ͷ�mL����^���[��Ip%,D�S�9�BR�#�T"]�3+gcs&5�` υ^�����C^�c(Lc�߲xp�
��%E��NŚAd�g?�ď�[��|�b�4�N�
�4����u��3DT�MY�y�'������?�1���bc�?{;YV�m�Ȭa}E<|�+�������<��0jb���n��&r�X���BF�P �PxG�+��-�<��[
n�=�u�t��ʭ�H��P��@O� `��RG�~�� ��b���W �>�
~��a�S��R@�Yf�Whiv�o��W0�A/���<���n\�;jC./N���ʽ�)�Ѷ�:Qϸ��d��IQ6�I���yj>������n�X .x�ׄk��=~8�����gNn:�4��Zبɚ��y�^�2j�~��:^} 3�.����ZP��ɺE��f�"�e�_�����ϓ����`��
��g�u��݆Lm�~R/��2��b�ĲbB��yr�������� |��>>T�w�{�U��]��u���s$ ����6��]yT.H�#����1Q�z��"D���R:%%���iRd��:��X�.����ʝ�kR�Oe{��^�j���^����a���9@��rRZ�r�'竅|xv��Dvu!��ӣ3���G����B'�JV3�����e����4�#7�N_��>�	;_#�1Sô��nWzj(��g���r��:+�=d�G?4�~��FTⲂ�ʝ��K��C98~,�gg2�8S�r@�zW�5���yp4�ڊ���T r�I��=�b�2�UN������R�?��<ha��dɘUyNY��#sI8ъ-zm~�C���)ROS�KW�Ό�^5�߆Lph퐖!j
��8<;���r�g`*f<�Ύ�T����ˍ�{rco_�u#z
VV���ٚ�2�'�b��F��A��F�UiuYB[�ˉ�tN_�v����ťl��ػFe�~fT�9{����OY+�������Ç��o����GD����rk ��/���E�����������T�d��@��ο���aO�=2���� ��,S�o��vǬo@+�e�}�|�S�E䃗$4'�o��d,��I�"�s�?&�-6B%AH��Ƙ�_N�OY]�c����Ҕ��y,u^V�.Z��h*��Rª4��:I��#Y?Z��6�1�+X^�Y���қ���.:�X���AZ^�h��peF!lA����\�s��Ѩ�f����sӌ)r%aq:�̴��]qV�������fm�b2 c0��³�>晫J��Y
ڪ���B	NO71���;KI�����p
�k���e�3V{ݕ-ݓN.�r���ܿ�DӒ�e�'�xW)�k홁�τ���~$ǌ1��l�~ɾ&��t�:�WgX9j�\�9�5֕�7G�{�7�.=b��y���r�4V���,��QJZ�6n�U�g��YZ�cj+�)��;PT�5��b6$�G����?SS�N��'�V?���I���A���7n��X�<J�^d(�M�3���N�=(�}�˾}C9[����֕g���L Z���@S4փzo{$�v��;�0K���E�cfp���y�g��Z3Z2�����U����g)�U���^�1$X�������E%�j���	6�ݺ{W�#y�>�[P��C�k�u���O0X�=~���~�x-�b�é��]k��6Z*�G�(j���#_�O���}��.ͣ�Xd{nY����Qv�v��P�z�=�Pu�źu>��Hh@�S72,LC@���䒔�.��]��h8��F�P�A���j��R�R1��` AK�İо���}��.��!iL$;Ӟ���M@h��&�I�i���c3����-Zϳ�q%��ވ�AT��Yɘ�[��~��>�kQȀK��%۬�(Q	#����2�S��]�_����t!�f@�j>\`����4Zyv XԱU�N�bylRC��Om��X�\ȯ�}M~���ʵ�=]�KN`�_g���w��Ώ�h1�f+�>ђ��fs�<~ C��C]|}P��!��;�(8�I8�`�Y"�?(mӁ��B�@5���Xh��`hԕ�NI�~G�X�y)�J�Q_'02�������������;2^�ɷ:p�\���[*�ɽs)4#��rX���I\+Z`�+�D�hVqmu�yj?ӾiuU��W>��̓ƴ��]��4�M�I���M��Dok8���~�ZL`c�������@�u��6�J>k=�?g��6(�P�d�?|�X���ՁW����" u�q�(P<��ɩ~��L��^W����3���lC���)�E'x�����{��8?�f c�+P.A�}��	#������T��P�\�������:�~���s�='�0^�;���M��|��oʃ?�*��̉μnK�I?����CR�/��/��%���O���lyR��MZ#6�A���ւΊhu1R�sy�&�aM���*ޞ^m�h�ed��\�	4�] c�(��CVNA���F��]���%�O\�^xy�S!���*���� <�<�تo5�ѱ
��]��љ,/��<�	�(��B�7�g�(��u��fA_X6���/Ή�hݑ���	���b#���A��&X!z�w�m=f��x0e�|)ԯKZ&��C_��P�c�qH���&�~�q;���yo��}�����֔�:����&�
��Y�P@��LW�L�^q�މ?���KZ�҃?�,B�5t%͸�N��Ϗ0h;[y��}?Q��i{�v���.�^3��lY����%`�@jQ�6ڹ����z`o��QY��z�T�W� 5�*�QQ�Xɬ��k�IlIA�e��Hl���X�Ƭ��b[��؈ޗ
�*�K�>^��ѭ�s\	:�g�e����~Q�G6/ЄA���V��F�1@Ci�#x)��g~�K�W��x�Y���H�������q]}>֫���f6�Xl%�Ш۵Â����#�3�e��J_�'֧b3�T,?`?Վ���Cf>#ŘĔny�!s@�vϐ'S<���Y8R9L�!�[ U�]x��9����^�o^%Ƒ)ɼ@�m^틷liYy�?gI1�� �Ŕ�W�J��ٗ�Yu���mW��ĺdw�D4H�3��y�����u��և�q�ò���@�3������-5P`�P�fv9�b�e����I��+K}��f���|O���~��奼���%F��DE��{�X�v�@�M&ge��NB�Mv�9I=��=�D�����p} ���G2��	1YW�����׆K�v\��Mo����Ejg)5]�F$�3�A=S4��"�G�L��.�@K�g���&�^yn����>P/��E�щY([_^�~,�����o~���^����3D���iW#���u)楼u��3��P-�J�:9�:�'�,>�/���%�g�*L6n����E��1�[96JLv(L^���|6�*�X�\nwYg����_+P\˹�n�Q��T�aޣs�D}�w������З���)'����)��/���D��r	��&��`6俑ɂ��=т7X���g_�Խے`��Mc�&Rl��D)[ĵ�g��>[����n��_[����: ;�
��j�E�-Jn���j��h hpv�g}�#�<OTZcKE�:N�9�/��h���~i�R�E�W�9%1u��lpp~JѤ%��֖�*ꆩkO���wߑ�ɥL��ϰ��:�&��k���Kj�N ��X߼~�ζeĻ299��ᘴDɾ��_�/��E���|O~��Pfg{GvQ�=���1�^��Y�����o�N���_����쳷�^�3_ʠӗ	Z���T�f�������t~ġ=���B��:6�)J��!���+2\���ulUR$�k���S���"h��p��*�7�&�V���u�-4΅��V���`�V�f�:1�]Щ�҃�{O?�d&*�>�Ń�^�R��k2��6J���Χji����H�>ߌ5:Ua�4��[�_�Y�,����E[��]�k�ɶ�כU&�D����A���f�FTկ��8���, ��:�+\%./�Ъu"ֺ%m�i�s!)�4�I8!,M�6��ZT*}9O�1
u:��yp�H�E)c���|��Òk&�A��Z�F�k���[>R�F�=<�R	i����
�#�Y6��Z&!�F�YN�@z�j��<﹙�'P;�m@��g{[
���v(�B��*f~��C�Yf�J�b�z�@���8c��F��:�H�J�����W�FD��rG�*�e ��u���hOH�W�~����u�T�������c� w�|R�GHJ�m���W���p��7��E&Ӊ��ؗ�[�H6��bgK�<���2�G�rxzɞ��k����C·�Q`������6���$A/]�%�I��F%d]k9���QE��nC���Mϲ&1�1�y���dn��&p��ǐ�J�1Q��l��|-&\c���AVl�c�X�٦�!��ڢD����ՃGrv~�w��C�{|,��Mܑ���"+~�W����v���eN���ە��s�9�{��u3hYt7��,�k`w�g{��=�o���;f!
{�we�}�:u���b��P��$��:�.��Ci�p8��J~iv��ݷ���*Ţ�#��s{�Zj�	�%BI�ck�5��qP?�B������V��5ap�˅G�Ƒ��Ƞ$���1'�G��[(+��H�C���@�u]�+�7 ѩ:Ҡ�f�*H�W;�c�X<z���� ��b�_υz�E)�p���o�G���[�:�?��O���\v�]�D�㻵�%��k��f����%��|�@q��0�b�`��0��NցJ�L!�t���b�uQ�xM//)#?��@�LT�nA���%8�S��߅���=�k�"�C	�bc�wO������,���;u����ȩZ����G.�����Yn5}j=m���- [�8�J���t6-rV�f�8�R���L��a��?E�@�Xycz8�|/j S��FƖɩ��i��o����AK1�Ĝt��v��s����/w\�F�ʕL�d�Rg�ҝ��e���)���n&G�	?�'o�{����1��-�Ѐ~&��)��Q�c�#cH���')/�����X�x^L嵗_������D�h�`�~��^��k��k�Go�D~��~]��?�����(_�������G?�1i�l�� �4�Mi=����@����R�g?��CBVӋ�E?Ģ?"��"-�v4
L����,��`��Rn���c�Y&�*�wkȝ(_�{�@]$�Q� Ie5��K���j�\�(Ħ`�ڎK7ւϣ���b�I�Z0���7v3�G�l����.r���~���L����ƶ�6�X��ɥ��Y�+@Ld���j��f�m@4��Z_��p�S����XQ��i�>a�7/OM�-2��7K4<q�k�hڑ�|vο:C#M��k��j+��C���v�qF�Kw>s�Gheb�hi�ʣՅ�	I��Wb�n�g �1O
p���� k M,-ҎAo^�ܘ�^Q-"�I7���
���{�YʐG>QȪZ��ɚ�<���ͧ�P0��I�5���h^�ynuLi,��Ⴠ.l��i��H|�����:j��X7'���Gi�1Y��ҕDi�~�(sz���Ӽ�-�XRȒ��xF�@�Ǜ_��-`l/�?
�������F�PކC<���"�4�Կ��� ���qu C�r��j�͛��
N�����s����w��z�H�>��� kѼ�K}�T��)x}YZ/d������m���c��sۓ-����o_|���tsGz����#]�k��d�ٜ���-X��FJd����e+	f���=��%�~-XҤ��[���<�ql OA�h
�h�Tf�=$�ݿ����̾�k��źALl���3�2ʁ�8��O�fB��-����]�ޜoT+����s�)��G�w��xB����sSY�J�l�e��kܱ>a_���t^����=�;��uȱZ��ɤs��'gG����W'3�O
��r|�~���	�����Y��g02s�6�j��]kqe|���jQ��^�iȲt�]rG�����V]��gd����3����b� ��R�>��ߛw����Op�Uk ]%�̨ �1I�*�o::?��.�م|���r��p\;�9����S}L�*����0_�;�֛%c�R�.{n���P���C���)o��r���8d�{o0�_��o�o|�7�T'׏�'O.�e��&��I�؃l-j���w�l~����F�k����ܐ������CBj&�ɩ�?�綅���t9�X�K]����*`{wy.��7r��e�S���h�PNA�A��ʹ���<=��so�I����Ww������R`<��~e�|?�襚���������u�+ԯ���@c:��9=�H~Q���Y3HKC��B���@�5��Q�i���;كS��������L��c���2� MP���vD��F �02V+\Bc�,���A�xأ�Z�\F��XT��42EXg�}��:<x"7�;�?��R������2�M���僳���S9??�W������o��'�����<{�;���|����~/ݡ��^��7���7e������Pw�u��Y�d>UP3%%��ZYqP\8�:�LU�E��|��޶�I��c�)>�a�
w�Qg�Z.�ì��H}p�+SL����������嶣f@��'��Ѕ���53����kk�Q�X�:[��/�K�U�sYo(^��r������kr��X�D�L+J��n�YR*= Y�0Gr!������՝d.��1��@p��j��<S����H�c��=��
N:m��U1�bF��;?���^����e�r_��c�+h�#�-a͚1�ȟ�)d��1�Q�\ƃO���h|
\�~;��+K�Ĩ�]�x����%(Tϐ4I�S6�O���6�?l����g���d���]yp9��P�Y Z  #0^;e�J����5��FbuQ\���"̺�.�n��G_'�����U̐��4O��h��8g+ϞT�ޒ���"5543�c�D롙e)��E���I���2����$�/�r{�������R]��A��ʉ>��1&���b��4��X�=>���z #uЩ@�_[�<������#Ǘ���<]1�m04�I��s�o����S09�:�M���3�$��ء.K�����+Gk��m|%}��0z8�H+=@b�@�x������sb~d3D~E�$%��Z�-��l�}�Ÿ`�B��2���8�&I=>��@}�~Nu�}��M�-��Ii2���t�U������9��u��������}*�B_F�H������x����=�P��R�ߋD	�����SB�L����^��)�}��Jd�t^�uܹ����Bnݹ��pL�Ɍs�{%C�*L�i��U:�+�Z��;.���},k۝8�	�Uu��ꀈ?��|�*ӹ}2I���f3���_�@*�o;3���$Gb�ָ��)����.f2]��o�H������w��l����9�j�����Â�r]�b}-�m4�;7n�r����; o����SY�L�dg0�3K7�/_��W��;���7�o02�۹^{�ic�	B��kQ�J[O�;de����u��G����&�q�
"e���*��� pGg�2��b�ٖ��sm����~ 
P�Z],�-]��_��FM��]8s0,�mU5� jK�"r�9r#]�}.����ˋ�py�4�Dk��Z4�gx6�T�`�I�l����
��o�rW)xV�;w A���y�E��S���� �]�G$�/&��<������z�8�_z�D�[Y�X(�f�ش
n^����]�ht/����V��(���0�dˊ����L�����!]H9[���}��c5�7����{S�t!���|�����K~�;�#����Q���'����%6Q-�����`Q��;/��`�v��	�"���r.�!���q:[R%5$Al.P��:�A�%��f�,h�iӫ�?CP�h�K$�+]�QY*�"[�QR�-S��Ts�,�W�@��2��8z�̚���N�U�z��1T+�`�'���1� ;<]+�1ߛ{ �)5YK�#[:��О����ѡ:���exc����@4tQ�4cf{�����y=�CC�kS����omW�̾����u}e0��=F�ޘ�z����=-����+Ȥΰ҆D�*�Y�;	f���6�!%2�{qH�p�9o]Vk��?#��v>��y��j6B���y�.VldM �lL�-}�%I������x�A�S
�Cu�=�9Eg�u����Բ!���yt�Do6�`
��{�`����H�򄕃ƕ�tE�{���K�j-�S�E$[��ﵹ�4>�I1#`k�a\�Up�Yː�s@���8'�ڐƗQW��Y�����\�4N�P��5�7�q{{f�O���}�.�b,R�d�_;�\K������� ����>���=Y��� �4����k�>᭝krmo[���!s���+/<���3��$�[�V��a��4 E}��:�l�+�֙c.�1gtK�p�6�`� ahJ�64B�����1è�,�,���E �!�k��m�,O��D	��X���<yT����W�7 ��ڪ�"3���Bo`|ͿyV�L�o���jHx#%i�׃nq�k��r��y���7�/G�w�w���Ug{E�����&U*+<>:R0kC(�"��F�b��P�F�W�ȱ���h��2�K5�ZP���ϘIDP���[��
�
�)[������ d��Z��s�Y�Fe��5A��E{�jP�D��1�B{_��Ś�?�iߡ�c�X�ț��wT�|`e ���V�U�M�K���=��{?���9<9�b{d*�n��`.P���mf��W�x̣"�_�q��B	� �J:�а�ȫ/�"_��/�{?}O��ߕ3ݼ��۲u�|OA)���n0h}���AӒ@�ƕ��ה�/�����d�0�x7��+��
6��#�e��O��D�+Sg=�&�\�E)}u؃q$����D�}���9ϧl6��6���֥2 �Ϭ蚑�nF�DF*l
�<�k�(��	Ѫ������NT�j��{��&�������Ųrm@�TDS��մ6��Dxݒy=JF@(�@�&�j�J�c�3����lu"tS� N�(`1���42d<0��V��̢�%e���j���:��ѵ6#�
!��FH�.�UT�NrǉPCJfۚ�t^.�&���	Q��k�,(� irq�9� ��≜�ߟ��Aߍ�QF��X�����n���s��35�E�J��1֖>�)Z����L��*�/;�"���h�5�Ɔ�M5>>�H�ϩ����2T�k�X�X=E�ȳ���P��7ռ�H�q�盥(U��E�����3�2�B!Z=C�1,�����7u����v��oX��s�Sc����Z��I7g�"(4�S��(��Q����UMf���)`��y��hx�ql8��W�_�CX6�J��Ib�:ӳ��Z��A���uї�W��� �W����g{rn�?��K��͵���M�jJ#j�����gY%�`{� �����6F�/�9�����)��pn�*�����ku�$��m�^��V�B3^��^;�e�$qm��2���U +�:�	DT5���x����ۜi���9�6>c�)sEd4����f�ܜ�����Lt�o����m��[{o?��]}T�GY�e�Ѵ��8L)�`�Uʙ�����5Bn!�^6�ϧ��zQ��+��� x�S�C���1F>��V�@}"0��\S��[7���kl�uqzF:�X�-Uޝ
�ڌ0x ��E�2SI�z:K�
��)og�3а�R�Չ�6�����g�ػʼ���Ff�L H�#�H��S	�6�)ђi�lOK�4 �Ƅ'����샙Sa�-�����L�?�k���*j�Z�%���I������=�h]YOFá佟�� �\N@�D� 0dF;I��V��;�y|��N�����J`���VTk���tʚ�Ug�DGO��:�y'��l!O.�����\���@�~�E�F�����b�6�ѵ�Mh.�/���B�3��7�r�⣡��?SJ�E>�4��k���h>7֏��u���ΡO����ã���@̒S`��C/>]��2�Ld	Z�^��}9W�z�3Tp��;��f�A��*)F���R_�F�t��\rul/.�2=��'O�ݻw��/�����K�����,��ߓ�>��| 7o�S�c�Nإ��d&�^/�p�c��=��bbS�
�^+2�î����>pX-8�yMb�: �h�s*J4��2C����0�P	Zf�  �+���	
�bWs�q-����V?Uu�re����U�P���J�x?9?���O�xZ�kH&���N���M�@6�+$~�L5<�r��8����x��z]֠�*SI,��
K �h�j��J#��F�b�[��ʤ����ݠ���qd���׈��z;�YE�^�,��Ś�hcĈ_��q�^Ra5�������6�3f<Z�9s+��V����������!�
��زB���5[`�!P��"���,��s��.2���i����ӹ�ݡ�MY�e�s�\w����T�Ģ$P�Q��12D�*lXjt�ք>�����	J@P�>S��Ҋ�Ce�հ}�b�G���ƅ
3��5c��%Y�!�M��p��ཎbkN�Z�L���	-���6mSf��u2(���Ϣc5�3�OQZ�Z����\�ƥ̃�8q�ǱCj�c�i�:jq 1 �¥��ZS���Y��b��j57�F:i�Z�:�i;>ߋ`jsM�	���s9��3BSF���]�p#�ꟿvua�,]�u�����E�7ՑL����wY�r1����P\G�`�NNte��g���#�i�dL��o��r"�3��em� �S
5�����3�XO�L��$�cʚ�Ʊ	�W���R����)�`���1Y+��X ���N�Q~Ltx �����#��30o$�&�&�NqQY�L��'�����P��F8d# ��@3�V+���vD���hO�v@�����w�R�/ˀ�K�=Y��=�?B��g�͖�y(w��	���\Y��P}h(c�/����kM�o߼!�n\g�秧T�o�=,׹&r+%2� Fo���(0C���`U과�������T�Z�U���l���K%2(%s��֢"�7𲴾�k�V�v�Ddʄ�H���|0��)~c�y�pa��X�����j��u� �g`M�
}�i�-��e�&��)F	%��J����ub|͇��&�TL����M���]y����Ol�B�K�����Nu�^��
��Чm���B m!<x`��TV��������X7s�lGc���/gz/+�O�:�<��gO��遬����d���~Tp��Y�-Ҵ�r���ҍ��V�S6%U����������\r���n�m`�Ң�x:�4��M�>�оP�?����G�L`����`Q\7}�X����Բ��tP��[c�=�<��cE��/O(�.��DD/�`}͟�hHS�@s.#�{�Cyp�Cy���|�W�}������U^߾)�3=�[�Mu�o��n�LEƥ�KQ�Q?lX���Ag�5��c0��ۢb
�<"���~�Á:�CPf�U�ܩX,�J����>����b�I���|5xS=Df2J�[cwVH2�����CK�Uե�����H=���g��[�
_'Ӊe���>�D�r��x� ��G�M�(����xY}�e��!���^a��W�#�f��C���MR���Rf'I��E�P�\z ���~:�K{~��2��h�z!����ŔY*�DͪD1ko@}�u#Ў�j�j@�Ʋ!Q�24Nyr��O�%'��֎=s[���~�We������4Ĉ�E�'+\	���
�I���{����Γ���������U0�1�ɡ��z�ɊsW?�OVkU�r�vFgu��=�c=G��7J�q*����}SΈ΢�C�"���ik��ا?��	�`3M�X��*z��^�m2q$D�C=LX#&����3���y��������v)�2w�D�gWRlK�ʇT��
����9ńP���6��k)�
FR�6Wf��+{O����Έ�ut��0�n�,<�4A���}��s �6��v� ��S�3ZI�wp@��)={Kic{�FI��g%S��ى�5�=�<8N���)�N��u3F"[�)S�
 @��}��]������ugϴ4�3ΰM��zϤ��|�&z��4�����˥YZ�:�0��ʠI��r�b+�{�3Ƥ�^og`�l]�65Qj%Ҏ_�;��Ոq�)ժSû�g��X��G��1���-Q�5^��	:qn�f+����W��n{��m@{�㨙�?�Ǖ����G�:����0s�7s����}�l"���1u�N��&�`O2!4ؾ:�|������w��؜����D	�螬g��ؒ���d��� �G�Ņ�ǌ��VOF;��#x���m G��� ��$�2�]��oʇ:5�o��9}��Ys�d��QFl��a����Aj�BӖ�j��63P���S͢�����r��br���YcN�Zͺx��|&�~ U;#��Ջ[�y�D)JQ4YMf�
��l�-��ZRyoū$��=c�}�{������7����)K����ş�{{#�7��7]�����&�%�J0��������T�uC�����N��B��>�E��C�H���C98|L?-�n�xS^}�Uט���B}4�k͂��)���!T���q�=�&�d�ʋlPd��(" �v��ne�7`A�D)�G�8F����؀�ƹN7RG�ss����~)M}V��wu��%G�@B��٢��P���ewwG�u1��C��j(��}I�_�!~�@���7����K����.�ͺ;���j!�4L.�srk4�/���
��t����afl�|��/(X|(���_�׿�ey��}������ߕl{�:��=���p:�����
�u"AZW����:��y����	]VrYY�(�I�&�`��i�\�	׃��p��&�����,!��(�����%�?D�QП�:6��D���ue�1�^�l�X'�����	_���Ձ��U76g��1�$QŤQtK�H��h�����ܔn�S��UϬ�%P[3��+�n�,�5.Yo�F <}S���z����s	uv�p:唔�����9znQ5d��k�a�|�"�x֩y#-++���6��W<)��À>$70����k��*�NO�߿E�=�f�Yl�Fu^z`8����rxr�J��;���u������Ao䪰P�]��d�kd�kE(�T�c�����|�g�;w� �@mXsb.�ْ��O5,�j������d���gT���Q��H���Ӕ��i�[A�t>���Rڅ�]���$�:Ԋ��\ԾL�$�³�n	�K������16��dz,,�VPg�A�9ӵ����6����L�֮�&>s���FIzo�鐡�U�jjRp39,Y�z��ѕ��y�I���]y�1�:�9l���&��Pi�\g}�����b��})�{f���F�Ƙ�r�q�eKbD�u�3Yǜ[F�L���k��U���?��ꆮ�h[+�쳟�=��?�"_�i�y}4ɚ��?��N�,YP��?��V�4�i�]!�fi�Q|XA�5ff����Wi|�����j�K�/{=�HN2��U�`M%�D�:��3�w{�ߕ��Q�k!:r��m�f��<�g>�cP�^õ彎��9��J8�I��T��H`X�W��3�人܏"*�7�o��+�,�D��ۧ�؊+o=O���3Vx�ʱ
N�國�5e�2{+���5�=��c![2W��ٷ�Mz�6 �X��~�k�Ŵ`@/p����N���7�ŚX��fFF��Y�9�v�R���J�ZC��G�_{mm���m�N�!D�_�^���rRr!���g�z���m��~jW���U-��*���w�5˝[w(�t�}�+_���399<������B��\�k�{�B%��J������׋�y���e6]�����H2_A���o��z�N����P=>=�kׯɗ��%��]H��i�db��w��2�~��0/�2+���ZOЁo�LE�j�dNYX��k������D]
��l�Χr*�j����N5/	ᦣt�V�]H?���O��=�0��e���\y/Z����~���B>6�
Eg9|�P���=:����{
�t���JW�S &��;�E胂��*�����ȝ���� (O���T>>��(��P�ɟ��{��?yS( -�zld	�H��F�����bϨ
�#8=;���C�Sc��,��b&��-�`�ݘ��X��:�m���+:�Bk��1�c�{�`s�"��s�� �b�)K��V��V��h.$�I��HZ  �؝���MsJw8�I��6ӕ&��N3�2��X`�,`Y:�g��������e*ԅ�q(����Ed��NYRIu��4�m9(�C�i��� a����ÃmX0�a}�5�-�c!:��	�e�g�upu"J���)cD��Y�B����=�[��'̲z�t���ɵ�[VK9Q�g�Ѐ-3����=·ڎd޸')��VK�c���������� �7 12i��"P�p�� +];�2mV���-5��dȀ�<*�鵇ڶ+Q-���ab�?#�̍��\7'��K��Iݮ@R��`�8k5\��A6���e[�!��YnYTf~�Q;	:"���a,��iۄ�7!�Q����~���=D�3��:
ٴu��	��H���F�s�����46�Ϋ���̶�7���;I��'G��5�^s�fς߾?u��n�R�d�}����v	��3�Ofr	��^yF��ZPL���@�����z�*�k�1�֏@�4��l�]�t(�#ЀҳlrU�]h����n{-�T�k)Cjt��^jـ �t-CXY����r*�r2�v�ٲ*Pɗ�jbR7*f�W�>��e�H5Tv9Uk2�x�yզ|V���E����-��]�?;�f�-�H��2��͇=�Њ	��tU��tN,{o�@�go�!�}��"5�m;��H�Ao�ӏ�D��G
&��J����+�-(s:�bm���Z�R��X6ϒc�=:g|�#Fk�C����c(M�\��Fܳ�D32?j�P6�r���d6�>���A���`�$=w}G��ܥ���.��8���@ZqpJ|��4PX'$���	���
qi�B���b�nӾ\�#D��`%5R��0ޏ�t�}5�_�OE��2�ݚ�x�S���g�4�5���'�����=��}�};�� ����ũ\߽!��G��-��?�+����-ѿ�5��6n�U��l1���t딀��㭑L�S�j@��b����ٔ � �w�NN�	袇ʯ����r���b}����~T����xj��n�#*�Yy����i�l���ل�!�|p�I%��c���8åOJwbE6�}��ȼ&YUO�z_I�M�	�  SZ@j����U�.�����uڦ��-�3-֦"�����*�s��`�ַ��|���������$��M��l�����} (����4*�:D]�¿���e���o����<:;��`HZ�yT�v9����W���-�<���D�jh��tal*�h�)�B�C�YDd����ji
��d9����p߹9�����g9��}�7<f�K�D������L�ƍ�@fS��9����(8�]�s�1/��,�gs63�h,S������n
�����Y�`�L�h}�RD�J� �8�S^W_�s3e���4������u6�B���?�G�i�+X{��� ��&%�9��9���V��&`��
��nO��#��a�p���<�⡾���b��H�=\������ ?�2�x�j]����,��ԭ!���	"H�QRAtz|b�� -j�f@UN�հ�c�"h�oೡjy��#�ޥ��[��i��1̬n��^z.P7V���F�:ts�AgF��	�+֖U���syR�SU�!3i��;�
�m��l�~S�~�i��fy_+avv�ޡ/x�YL���<�3)A��h�T0'�2��eǜ��A��Yg��؊��"�lG��a/A�òÚ��\]�3��tϕ���ʽ�w��h��L���}61�S����)�Ns�wg�NvkL������6V�q����Ѫ#��^#�uե�Y�w���u�tH[� و��A1�F�u�C�  ��IDAT*ǅѵJ��[��(�)2ԓ)E�0ǹ�2�ޢ�`��/�-���Aط/do<��f��(|��EdĻ�b��
�ؕQ���&!4I�]�}�B;)k��~��<�N�hHf+��@b�����荢�7Z3���0����3���ؚ+�#R�{mhpyiTV��D������V�_��i	�xR�LTն1��O��!$��gх��,�]^h $��2�l��0V)`�����?��>=�t����,�g�E%�1k��cYx��2�f�E,�V1 g����>��fn��yx�h3��h{�T����\C���������yd�`m�^rt~Nۈ ���^�q_��ƺ��/	��̵+gM9���H�P�6sC+��5W���V<�Ez~ZC.0f�״ �iQ_K*�������01�"����`>�ҀO��&����.�*X���H�CQ���ut�q��YG�_���c�|�=�wv�d���(�@^�M�l���Ey�{?���S
�`�·}A�,�@
��������:�A_N���?ߑ���� ��g'dg��'���#���<~����/}�uy����]�<�/���R<H��m�~6Ee���J��LS��I/�!�M ��k�T+flP`g,��'��kl��Pj���i�^I� ���u2��N8,�;ȀIl6�:��7b��.~d�����bB�9h��iB�Ǜ?���?y"��oɷ��5ֳ�:�g�ױv"Zsf Jl�����K�B}���?��?�7�|Sv�#fG�Q_.2��sYM�������s�MQD���aB �zEE֥?�XF(ZV����x������92R:ru����iA Y'(����M�q���%��C��/߾%�(R��Tf'����v�ZX�1�H�N�(V������8 	H	�Rg<�LāY�%j�AҦ������ml8g�k�����k��5fP��;��^�t�#�v��f��؈@I�(�c74\j �V+4�� ڄ  ��Rf�^{���(qP�%Y[�k8��Ak2��PPC4�������(�PQ�"��0�Pc�
��:���;t0�s U'��2e��L	S����#�����%��b��'W{8I��H��Ṗ�r%�.��D��^�j��ܮ�"�^�e>=�S�P9� �˙tG��(�Ƽ�a��u�h^
vY���-���@C�l֙W�cM�)d��U�חY`���q�8�R�z�L::��Q˦6\w������	�3����M� 4M��]ae5�M�d��7�A��k����	f�0�,y�}���̢e�F0�!�����<�WYAk"o��$`cB��ɑ���x=aʤ��β��=2F6V�0{U(�,�L�t/�,Y��������@�O��X') ����T�+mE"�RJπ�T&�u�:b�O� �}'���m^�����8jbl�вg���g1��n��w�DgLT��6����Ԏ���Z32R�0��*�D�3����u�5v�M�WB�d��p�b�v��k���7�g�^�sw�&)~R2��=)��B4�|.6�ŀaY0�\�	��,�;Ԃg����I�b�ZD�?�jF��
0����-Za� x�y��~3��ɚ`�g��^�bPEL*�,�׶�;���!�/16c�)y9���
�`��Z9�u��l��,�\N�g��ew��R�L�_�g���M��.՘�0Ě���r�Af�Ihx���AH�F|K�䃯��=QY�g�y�J�>�
 K
��ܲ�^U��`�W�= MH��5�p�y�� �ZЄ�B��})1�j#����j¨�s0~��-2�|vqƄ�y�Щ����n��Sy�ͷ����L�]��aW��֎�����C���J�[ͭEӃGd[A%�S��^���?י��H.������B^����a$&x�C�5�@?��R�L�F��6+���P�10F\�S�Lъ���v� �A�ş��0Wd:�ʺ0��B�㺇�js��2e�0��(���"UO�Ed�g�?�|����T8�`�F���1J�o�����\L'r{|����ޑ^xA��o��98=���D7�K�8pJ�	�pfw4�����r�6�����s7o��e��I��b�2�X�`<�3VlVî:�+:w�4t��B&�� ym�B8�Ȋ �=p�w��Ɇ)d�BC#v�@"��`bfi2A�?h��o���C]`����Z�,�ݽ.;���}n�/Mw����j4��Y*x���b�H12��+Rк
�a������ʀ݃P�-˔�����K�g�()�����Vp�n�C��&[�B  �^Y�2����>݌TY�ǣ)
��G��ZT�*������j�r[�xR��قs(p�FF9���>k��|<`A}:�ʻ�8�U~�:e�ځ�*j�b,9�>z�dVr�ھܺvM���kjd�����nm��<��;��q�Ю��[��3`@����7����=����mX�uCs�[���dg��s�9�:#Y+t���l����af`=7�4[* ��Y;|��0NE��1l� NHs����U-�����F{�����.!4�y{�����0cJ�g(�P,�ޣT�)�!�PQ�T��ٻ��h+EdMo� ��N��\$%չf�Y^���@V�&�Z��`���5��G�}�9"�BU�<o��͍�z^=����q ���)���`m�J"7��J�7P0�����@��e�c�(|�$�tU �NVR��m~0�|���Bz�Λ-Yu*�����v �$��LYL�5�z_w)���lBtJ�d��(��S<���7@��Z��}f?�Y�Xeo>�DoKY���u�c�M�L
^��Z���r����K�]�a{ �l����k��od2��`lø����f36�k���F����V~���p��>Yl�<u �����ų��Ϛ,t��Q�^ЧL��Ls����O;��s��^�f�9�$�	�ٸU�T���y2�n���DMB�L�QƠ�8���X�3���my�-��{�B4e��d!�>�m�Fcݛ�o9��i�`�9��F�km������׮������G����P���������D�4����5ߝ�D�zx}I}�D-�Up?έz\R뜢T2:I��^P��{"�]����=���p{�i�����?��h)�ߋO��\e~��x�`)��y�I/�e��^���30����7�'��X��oȍ��2V9��?ܖ��o���Ӯ�����zK�cD�e\RAW�ˊ��E)��DF;#y��W�嗟W_��8� c(�qاpM2H�_��9�3(�:0�[��'b�~�WL3�4�:[cp����>wo��'r~vN�,6�T�dҫr��6�y]G��Y��8ZAia*B(�M�:!�/�� ;���=�.�����zFpk���Y�
R���#-|x|,�>lm����{�+��y�����w�f-���eN~W�T�#���B�=����k��w�!�,���;��1R�ٹx�s8�����.�JÎ\W#�|o,��C��؇�R��¢�1��*Ԋ �����Bh�0[�1OY�Pu�	N]7�ȵ�k
(P��tv�~����Ð�3��F���b�� �YR��7誁,�̎��Vg�?����, �ê�1`8fs99?���#9�]�:i4 'F#�P8���y	�Pn8=J��)��% ǾDn���53�ѡT�R%K�T��y���:�ɷ��=X��.���6-���R]�ϧu��ڰ�hE��.�]�TѾ|��R)ыFqkgG��@.�/�O���g�^�k
��o��96���]9=��w�G��}�����L ���|���L~��X�Q��� =�W��YdT@U� N���`c�s�������������� ����<<` A�=�7o�R��������������@9�Fa�}�ko𭟇�m���A��[��eװ��5���d��Z�
4ڞ^/�Au~�VS�ɔ�bR�eժUr/�&Ժ
�H0'���b��؛���ava�*x���''�p���X�f
�����^隀IP H��m�9������&" uV�bt!G���D��%�D��TY�}D����J�8��N�Ϫrw��X�Ԁs8o \򅉍�� [:��/.� !Հc
Uu2'1Sp��Q����$o����Ym9�)�'j�]Hy0�l��[�QO���Wg�)2��զ�*�O��Q{�r��#�H`��I��s#��F	��nd6����T83�)��j�IIFLet��|ļ��S��+������j����	��P��)H����:���")�����ye^_��O�i2~�u?׫��)64�rFև��L�^�D�bb�|�Os�<w�~��(zUX��gT�Ul��Y�|#��mU�~~n�6���zMA��m�R8�JC�SM]%G�k�I7u�cG
|�#�|�^���q>���5��` �|�5�H�k*C����|*G�}��3
r=1�:�I�F���fޜQE�)�9���93 ��mt�*��sE�\R� �+6/ق(��fʨ��2�vg^˜��kՀ�>�d�L��&���`3��d��|J���<�cϱ�$��j���g��^yS��D����3�a���o����2�\}��|�k���N_������2ؽ�������ڕ�w��\�\��b����'����<8 �몟2+�{2�衽��n_����Ig�QkK����`�T���4�KV��й����(yjʸzHeSTFw~u�������8��bPAEɈ�3}�z��Έ�_;Kh4�5��AJ��������H$rTB_/���	��@��gϐ�̣V���@Zj+�4^��X�b6���ё��E@������m˩�3u�wFc+��	��G�~m�+4^G�� 4;�T]4�u��֯��|�/�F4��dJ��Z�FJ��3QG���B�7�D�=yH@���o~�
(�ȏ�|Y��_(x
Td�#}���ə:��}zN�6/���J�!M�p����9�
�!V s���^K��_��_��|�&����ys����{4�+���/��׏�<{/ݕ�߿G'ȋ�K�1�a9թ�sQb̦y���OP-r�������2[t��-]��N��m9;;T����:�՛��� ���h]�E9���T��Er
:x��(��U6�U�ut|./z��Sƅk&�#A������B)��Xue�շ>M}mzgrXPk��S�+�C���<* G?̃Gr99���  y�����lm��7����/���Z���d�@}g������R���<�y��o��,��O���G���)�X��U��=���!:6���_�%������9�k_���39><�B����loo���}����N_}�2�+�������]Nu3�z]�N
Ыvj{����F��}}K��)z��@��l�>�p\
Q�S�`�����(��OY?:��gGzc���J���ڲ>c�*�:�α$=.�睿GǱ`༴�S���-<[�S��n��� ���|�{��~�O��Z1�TB���Z�2���	E�T���&P���r����>ꌘg�,M�pX^wH��X�ZB�_��0�ޢ����OB�X'�;���7��&�v�XgЭƫyhAꀻW?/���s�ʭ�T���hy>�l2���w��=��$Ә%��S�[���As]G}��\UV��$�A�UI@ʹ�#M�(�Bt9���G{��4��U�:9�)K�&n�C���ɉ����9J��V[V��t�ǔM���#�B���ZR�r;���\���6���#��0+��g4�s`kX�TуC���MK�fgN$��SI�g�6\Uf?G�4����ب�l%#8S�"�z9}I���[֪Ӝ*Z�����^0�]�)�^Βy�u����h\@v0�g���*�e}�}�r����%u���B����cytv,'�K]^V#V:;���Z6�|A��P왣%��2�단C`&�k�����,w���O<�cꡞpH��C
�� �C��`~%4GD=���#�YA����5��f�AE�^eu�����ٲ.1�%A�U�LA���G�N�ΌB���T$����S���<3OJ���|�������)+j_��3R������\��k/���}y����?��ܿw_��<�S-&v���zY��L����g����Տ�\�`�M�r2�����%@t������ݒ�h�!2��D'�|(��JJɅ�hlڇͶV�{[܈�>�ȓ�����=����MVN2uDs�}g�x��D7np����Q�M�v�Y�:J�y�?G�)�ڍ��Qɶs"�w���.Xu���Cf�䉌U���Cɇ]������쒍�q�H�ԉ���xG��j���(��������3.������ٟ�O�ce=�����b�:��ݐ�[;R�f���~����T(ku��/�����+�(_��~������B�,�2O���L�j���׮W����R����{�|r_N���Z��� 8�޽~[^�}W��%���f�2����#�Q@�Lv�-�7�eg�%��=�)$z����ٌY���'
���5'��_�W_|�E������~O���D*��s��HPi�oi4]���lD�27v��oL�)k�r<w�jdB2��<�5b;�+�~N�ҵ�+W���n8�Ѕ���J5�D�^�y����Ya��0�w��ܽi�%Yr汽=����ަ1f�0F�2�e��f$d����A��$A�F�����Z]յ���%"���/2k�mڦ�h�ά���Eܸׯ���o���nr�\���:G֤� {����+w^�����{�|��o��s�\��������L'c�����2z獮�"u:pe��jY����[�������o}K���P�t�7�Ad��[����.���:�p�@�Ɯ��[,d:|fԘ����~�U�!=kw0������3�yY[�N2�kd���AI�����@�đ����`0JG�k>�m�ݶ\q�\U`��8�m�D�pS��1&�hTi�gˬ�0e����#�(NP��`�A�f���B�d A��(m)iQ�ȰnM�9qJ�cEPl��@& ��pр����Q�)7sZ�Q�	�h4KV\gp�e��H�ԕN�������en����D.�/��M$]ܱ���j"͝����n*�,�(��{��g��f�{U��IZ������h��DF<��`5�V��h+��V'�^����$��O��f{Ҿ?c�0Hl�����ĕ&��X� ��4��h��]�b��<�O���L��4��[{�4�N]���yt�ݎfY��@� �U{�ױG��R�I�m�Wn,���b-^_���H�G��W�[��v�u�d��-PQ�jt;i��:���M�3␜�~d�2](�S���O�y��+�p�E]��Xg�!���3�{���2⮛����۫���{Wo�+
,Е\�?sm�f$��$2Yr�}/�ky��<ҽm��p�� Ue Z�,e-�Au(����5[~!���J��Ǐ�����w-��
�R�����W`��-(���Y@1�H- �4I��Y�wE7�O��@��l�m�Q 8����t/tf���ަp�({��,Ms���2��4m�[��f�Fzi�T*m=�6��9�Kk��b .XȊ~*51��{lI������C������~E|3�g���9��h97M�7^Kq���	Bcd�d�@��V ���	`#Ԥ��2��[��Ο����-R���C?���$���9�m�^�T�q��t�}�;(g�V�������콆%����@`��"����u��uzۅ�i�!��m���.!F�^L
oŞ�ؑ�"����j.����� �e����ـ��:�$�Qe������;Q@�1��%�)M��ā��c�D�r��2����ߕ�O�ү2��s@���{ �~�-�SGx�^�/�ߓ�}��'���f��2cFr�N�j2�|�&���:Iv��<��6��0B��!C �gPFo�0�~_�
�
�.a�����|Q:;xD'5zÆ�YP��˱(�LA(Zp���seow 7o�T�գ�:P�5J8��޺I��j�&�c��Ʌ<�wW�g2;��E7����T
��^��,�Vw���>߬@v�
x��T}����l������bh�j��k�Xz5��GC[˞�^�/U�f��M�D�<��\�l3�q��[*��M��)����V���ͩ��:�(��s�F*;�������/+���H�I.GG�����ߖ�,eY�؋�w-2�dWL/MY.��% ��� ��jk�5�*������/�����������P�"2XOs5��z���v3�gyz*O�k6_�I@l�$��.�1�Q@f��@����d}��ۣOZ�� Jb=s�=��9�]�%�A)"�j#sS�k)�AJ DE8i���l��c�[e�fE�vC܉u�X���z?:�z���v�����9�Wĭ-�3S���R�:�'�?ܯ�Չ��[}X� �ֶ�DF:�ʩQ`��EP�[�����Z�� dyִ	W��u qO �~�{C_1h���F�u�̢����%߈�S@�*�z�V�Hk��L��L.���_��k������.:5��e_��xcuoPva6H�׹����{[����p=�����lX�	��5lX�g�j�}D�m�0f��}�zE��/|D]����(s�<"ت���0im��ƌ����Ƭ@T1P�_l[�����yW3Ql/D��`s����>�b�jt�V�e���O��<x�L�o|>{i�é�B����/P�R9J�mmJ��i}��[��W|�/P<�?���f�K����y����[Yk,��*2kM��պ��cc�n ��[-Ya��+�3	\͖��y;+�P4��Tذ5X]P������o�UV!�	��9B��p�)��b��W�WOvԧ�"S����=<�bp��~��,�ms��*W4�4�mFP$�['�W��?�$�Ʋb�=�E�����x�ϒ"�������H�5D�J+��9I��}2Q�@�h��G��`�����*�5�%j���v���`�"��a�r����?�g�1(C������Cy��7L�����D�h�6���r&ظ�O=:����ý�q=>�ev��׸���<�Kb�����VsxO�4\�h����´\����F�3���v�ÛB&^���E`-�`0�"��������D2D\�s�\���`��,��6j9U:, �_��3�UqQ��3��p���� �Uu��mt�iݨUxp��j�� �yGF����9y���nd�u�F�)�D ��F��l�#��8����}wn�.������?����'}��}pO����R�_<�q����`M����Q���r4��J��txx,���^�GߓWo+�:�:�\��P-�
b
��|�7ez4������\Ab/g
u��*M�����6GJ��KAm�~A���B�����
���8��Ҍ9�/�W^�[�������t,�ɹ:�sR3?�{��3}����}
��*����ˍK��(~B`T6�O�+�F�*���(3�Eǜ5/�K��hщn~ym��Fҷ���VԺ���a(���D��V���F�u�c��kt��W.����+�~oܸ��Ç卷�&%�֭�2�_*��Ȯ>�b��7�ܑ�G,?���x9�iR����s�+��`}+T�(!�sfv)]Ƿ_a������[r���l��eP��`��z	��eIO�z ��ܒ�/O�!�	5�Mҡ$��-�D�����O��jmE����l�l�	�$&�U1Q�ڰZ�[X�����§���i��
�%l��=�pk�U'�?�§�7l���V�fO5��o�F�kH��������؊!t�jfY��5VF����x�*���B�2�h2&�A�ՇC��@�/��,�dvO�X/D�b��ڲZpd���xA栏��6��z�թg��UUE�	���J<�Py��--(s:6a���̜�+��)��i����t��a��n��`}�\���,��V��Mh)�6��(��g�͍a#�`Jbmﴛ�m�#�v�c���֓s�3Z��s������LT��.r+�dV!����t�@hgL�2�������m����~ː�t�ٟU\[���@zbrvƚ�d��L�D5i0��ȒH[��]�,�Ƭ5�!1X��j�l�UKq�X�f�b��5';i�H��d�S,%�u�Yi�F�N�	D�)�����8ڧ���j^q����~�G�>L4�y�`I����,�Ч̝�gJ�-�� ��d�7����	�dE�v����@!f%I�����Afz������UA���@�b�I�1�SJh���&����t�>⍽]��kkj�I����ԒҲW�q ��j�/������D1p��H�Ce���E[&��j�������pHt	����\yQg��� �T���i���M�lgY;m?x��V���W��	���(����1�h7<���|���d��Ϊ�Rvr���L����;#1���k5��G�g/V�ߣ�]�!0�
���?����]G����.h0P� >��Z 0%~��gu��<�Nf�d���9I|���\�3׋/f3���1}F�I��"A668���p��(|"&W��h�>�B-6��p(#��������u
"S�C��K6�<;;��>���O|y��.��r��
Q�0ܑ�Q�:k.xD��b�m@L-�H�\W� �P3XNԈ�B��H���˿���^F�����_��~�s���{2Wή��Q*4��{���
G�*{>y�H>���^d���=�Wn�Nq83預�~(������
~��_�;�Od�¤���c� �����	��N�h�	�z��U��v)B{
�`b��t�����9::����zά�C����9�q��(Po
Tiڐv0P�z��[
���&�Mm˧���]���`/+,Z���ʃ�w����F��5����6�6x1��|�#�fZ�.��b�iEcT��4u*�_�]n�vᦕž���� ���4;HH���@�z1�@�������D�<���?�g?V w���R<�/���m��z��(�o��$U��O�S��op�zK(�..���	�>�{���4�U�u���#0q2���΋B7��nٜؓ �G[��90��r���6咆�����j]��dm�̦jϐ�[�E��]�5jr�d���d��,�Zn�4�)֜���s��D�H\O���u"ԡ(O�2�w"��"5�$�����,�������3�jan���֞��@���^Wb��x}��C"=)�=�k�8��&Yk��E
į}�u��)��6><�Y����9ǩ;ͦ�j= ��F��y��F��G<j@�ɣ�y���$���D�_�%fԹ%^����&��T���LŨ?�κ��:s�z*]�����.�h�;�C�{G�.�>9�rm��Rar��5�x�}~�l�-�5��#r�(WVn�d��G�kҡA��j8 =EɖWn���[� ��A.?��5�+i;�M���+۞W\W�+�#Y��$�`.��su<O�V����x����豘biֶ�B���Py����F@� 9�.@���B�is���2k��{+8Aa;U���g���^��l�uibS��R�?�uZ�'�y)���1%��b���%l1y�;3{.Hp�6.�叠�o+�6;�� �AWe�B�ԑX6?ES��>�����
�|v�-�u�o��!���i���ܹu$G)�t���Gm/Z�4��K��j������깈�cu�\�!o�"�U��`�FC�5�����.�JrhuT6o��X�hﴒ�ڨ��݋���@!�ر�P�`��$Sc���+��K.�rB��/�r���E1 ���,ѶŞ�xF�D�,{hZ����(�EǔIY#��A�Q��J�Լ���I�z͠7N��f��&	-�6ƾN���C�!�8�F��DT3n�`+(v�"��n
I\,8r��5�3��l�樓�;��`չ�?8�����4J����2�n��t�|�[6>� ��mǶ�ۚ="�Ϛ-4���M?+-���-��f�C���2��T�ͨ��ٛ�I�
Щ�I ��)�E��O�ʴ2�p�7���Z�O4����1g����W�O��_�7oݑWwd��{���|��'2^-dp�/�D�j.Ӵ�'��:�֐���P�Bs��Sun��z�z��{t@�{P�7�VzS=|,w^yE��7���{�dя~_ 	a�AS��[̛�:,�8׫�����k�	�������=��s�ѱ)������@���YGh^?����������'��z����+�@�NcК1W��Y�e��~�K-�e��6�-E�$�t:\7��|��Q�Ė!��6���>���^� �#m�����9A��I3?���;�ƴ� It:<�S��zY��j���A&L�x`\�V�	[������@�|�5��a�"���ĒP�������G:_w��/�ܰQ�����b���ϙ��Mel�?�ǿV��`]�J�3������Sy��!�yu`��B_�NG�	��
��L��pG���w�D}�>S(��@�f<3��i8����Zp�`1� �	�����s�	r�;��^f�����������;�2��W�NU�9�,��}c���y�,%-J?s���v��l��l"��J�˄G���z(RvR���휭�����l��%?�Hoݗ�G3)z��>k���>Z �k�GG:FSN-�P23�J�ޗ*O�Jk'�{RL+�{L�Ƀ@=J^��N�M�4[�E`R��T�3��8�[��Q�&���U	Ё�
�n2@Y� &�P9�)X�&C} stpM9D8�U�-��+��̠6��s<�t^X}H�����=E�!��0*QC�>-,��=6�X�ʠ����kbu/���l�6%��KZ{�g!ڊֿ�?��� iܫ�\Z�F�xW��Z�"
h�mK�M�4�ŭsXH�|6�^f�e��Y"=�3k�66�����}ͯ;l��,MI��:m���V/��kOݶ�Yڜ;^D��fL4^\ִ�+��f�lG��s�����A�:��"%�h�n�uz	�8V�f�	W���^�i���ogq?�Us��m��*]��r����(w������{껼��m�}�@�zԩ_���ZyH���$k��0M���/��J@�B���F�[�Սu������l^��t
2� 1���ź��^��r����&���ԙm���W&��`H�C���1���_�J����h�/9��M�l���*����@��zPʦ*y�Dq(�{�iS��ӹF%��l������'6b9H:@�簒�u�ʈv�r�F*0~��$l��x�����ƛ�����֋�x/�AFd����s1IV3x��� :,Q��*�$*�����h��_ǔ�ʊ�!d'0�%Z-�Wg�bЪ6�ܨ�Y�Ӛ�;
`�S���Jr�;*�7nr"(�>�,���S�;�����e'�q���b�i����78�c4�������~����%m!�d!o�ߐ�l_.˥��5#
p�N�/���|t�P�A`�*�d�Qȋ��]��Q@�\N����B�b"��y]��T^����vwe�`��2��ɍ�l	ŁL��Q ��`�?�K5?T�!*����k��WP���������C�~�Ϲ��~�Y������<y�@.�OX�y^Ա�k����%��@`�`p� .
ɑ��4xkYc8*�??S�6���V��*m9wE]s8:�#� �*�ö}}ܐ��}\��Ÿ�Bx�n��3�?�v��=���g�-��`�=���\Z}0zB��t���{���e�`(3}>��D^ݑ_��k���K��lL�� 	2�u��>��A*㍂Euv���b-�%�;nv��.i�h����z��kZ���t<#HA��t��wi���K x<��>�9�̞��{D �< �l6�g�:��񄴥�xN�jX���NLL��!R���g
��~�PvGFaD+��)R�n��2���~m�c&1R�����a܂�k~s6�]M�R�g�^׮ڝ �礤�) �
fw�e�X�DAJ9�I�(hܧgR�k*b�+@>����Q��"[���KFÑ�-�:�<�\����*W��[�o�2�qS�({��؃��ZE��>*�Z�&
O�)00:��oj�E80���:e]�:c �:<��1�!�Ě���s(���8��&�Q�WV� �G,�C�l� [Z�`� �eU"v���������D��~@"zm�Z��� �u{@i��2�6�|&���fc\@-5u��r(?�^�\7J���hW�4C�Y�ف��ijD��:����w�["��|�+O:�4�7���1�����5��%i��g�G�7����O��/� ��r�����G�|��}0��4�o� ��%)�/����ڽ�Q����=�G{�m�������seɪ��E:5�Bm��Z`3�e"��& D�qjtJPED�>%����N=	�����u�aI�j�%��\�Γ�H�4􏾱�/�3�g'2��2�%VO��Z`,d��������g�am8{s2{A��K����	�o|_&&t�=��m��9�!1��e�*k[*���$��4j��r˦{Qp�,C�z���QF����`��-�HJY�˓6+�+~֕�m���/;V����6�X�kk|��Z׬�/�ҟg&bĦ�V����p��p�~4pԅ��`~i�0�E��~Xﱔ����%H����O�m��rm<��!��M�=5F
h v¦��61O$nȀ	)c�^D�Z[#c(/Ɔ�0��r��Dc_G���l8�G���یe�cv�z��F#�ld����0`V�8An��+-ũj�N���믽�d,�冋Rw`ٿqĨn���û��ן| �.�d����\��x��0�[[�NL�T�M1�tv)�M"G�"G�<�\ UWL'��饼s�#	OP�Wr��TY��`�cm����i� �H'.���㛲���/��f�x�A�>=���s�s�}�峁(��ޫ�`��>�!�^�(X���+�02R�w[A�\g5�z�������3�L.��B?W��l�l6��?t1d
J�y�kM:���E�Qi
��B ۈ�6$eQ�����3�QP&R�0�1GA�J�V��`�}��UN��\���-����E���̃��Z�[���v˘6�|�:k���>��C� �+&&F8-��;i�Q�|/DG�i�Bdsq���BƓsQ��PpV�+�7�'�'l�������t�{��sf�/�An2�T��*�q[�sE��뱦���l>���6��Tdc(X�1x?��f�J��Y7����]d�x�!�s6g�`e�!���fh$n|K���h�rg$���\�N	N�=.&�A��i�E�ٶ�l	�E�#����g��y֓%_��H�r���	�gȊ�����L��6�Ta�u_]�8~$2��s/��݇2��dWnI���V����:��Y��k:/d�����GYqQ7}�Rñv�^��뮱�D�xe������!iķbxS=�ҨQ�S�H�uxvۋ�n�ـz��Q����'�鋢/c𠋫���w��t����$�u���|Ep*Y�{:󖕩d�Qk�N�@���xM3���an�A�q��;U�Ҳ*����\#@���-C*�6I3�lnV��Y&�3 ��5G_�Ǣҏ4unMB�)P�vꢩi��B��I�`�g�ב�.J�>1A.�Iũ�-Eэ�#Ɍ 3Lbt<i	��V�l�]'���g{1n�l���������b;*��m�l��\�:@F�	���M%��8�̈́�
�=#c�&��1�#�o~]��@��_2�Xf����5��Q+����`���N�͜�^���$��]��%,��b�6�n���ei:n��@�_"f���!��'Oe5y"���=y�8ŀf
�`�]V�-������ؾ���|t�M[�1�r��?�@u��v�1po+z��Tl%>y����s�<�7�դ,* Y#ё�"���AP�F����k۫y�[;���E0�h�XZ�R��X�`'���@w�+�ʵ�uM}w��S\#���auu]����Mc#�ߓ��H�w��c�65� �9: ��z����.W��R�=*jT�f��j%,��̋�}R�)��`Hύ���٫P�B�&w�{kp��4�?ְ�qG���Je�~袒5�<�rs��;��Ɏ�o?X�l[�Y8��=@͙I�~5Gl�)\!���UC�*�'O��Gʙ�$�k,8����XؾL�៫�{��T�ꌽ���;"�i)3u��M,=R�&.��MJ'r�跂�K����_ʻ��Jw^�H�.PeR4���t6��b<����l"Of�<2��Q�3C��U���p��D�������(h����a#^�rs�P.��uW��ET���Yň��j�����wM��j�7.V2��cړ5��m����{C��k
g���N]��D��G��y���x�k�m���N)��:�a+~peMF���ڎj��D#��bJ�;5r��f�Ļ�]|�'2ߺ�kF���d��o���8(�>�t��lL��� ?Q���h�H.�D7+]�KFwAu�Ίnn��T7�.�E���l�b�W�<:y*���`����d97�˴/�2*|��z���2��T�&9E/N��́��bb���7{� ��:�7��e���zgЗ���<�2�R���r*��\���Y���Ը:d��`��-�-+Rk/O��߳��MX�3ip�	����
���AO�o�lu�$�ɘq�U�U��t�T[�,]{�����^+2�x.����S]o��)�{mO��߻�ۓ����G�C�t6�G�:
l߻'�F�fG�P,ݰ>��NnS'��IV�����о���Ro�KR����a��� ��ۣ򤅪�(�$�@^E�i��t᥂�u�!3��g��(Lܑ��nH5+�kK���9�@U����$QU4a�.D^���g�&
/��3p�dG��vo@�	�ld�f �s�+��m跱��A
�� 2b��{�Zm��h��M��#&����v�=�nA�n��;H�����V��ӏHc��K��I3�ży��Ǜ���^c��i�{aF@(�����|�H��S�S�m��^�AJ����y}m�}�ьQ���@�����m���@	[E�x��O�x-��ѹ�^���k��M��s���U�ʔ#���* E�1Lcڨg���V'����ﵯ?0��,�g�k�!�����n�s��*�(�N�V;2�ȀW���:�ϟ]5���V��
���A�])	�B�i���|zi��h��`���Y��1L�yb�u�㰗�e
��@��ʄ��/D����]�6�o�j�+�!$�//��⒢5�3�W�g�{hD�^B�����σ�+! IY(o�c
��Ru
a��(��{{��tQc_A5B��'2�����̞��sngRh��3E`��B|��7����V������)�At1��Q��g<���k�fB�_�_�E�g a��)��n�� (v���ڀ,�Zo"��y��P��X6�g 1Ly�QM��\?�?��8�LG���9Ea"��}��Eٔx��&6��@�m�+��R�
t����Sf�Juf���SY(x�����l,O،3��8�+�BS�&�tB�	w�F��f�Q/�9lП��=�9�D>z�@����	>qc�v��6��6_.$9�&l���M��yf�@��{8φ���.T��ڲd��=�=�' O6S�����c3L�����I����w=�C������F�:T��=�Y�����> �h%�&�gF�1Q��j`�bwq�k,rk�=|%���9S"���k����M�t�a[������;x\�PW��}��Ä0�������\Wo�
˅���ݛe}�6�����=Ca��.� +#���؄�x���������3Jk�=M���D��H��H�?U�5��j0y
ݨ��O��6Ѿڙ�ގ������ܙ( �L��p�)Ɔe�eD��?`�*����������}�vH��+��x��B7����K�F=
`��O�`�0K�ґP�k�*)+����K��ٱ��S�¨6jV��=uj����F=��5�]�
���e/��������A�[�b�Z-a�RJ��rp�/��Df��R�LM�VP���Dz}}ֻ";
�%��Ạú�ؗ�������3o^�f�����\DY�8F�e	�3k�����9���\�ъ�����b�S�%^�`��L�
�I�[vX B;]��� 3јze핐�P/f�y��j�{ ����d��Z����Yы6d=��6�Cs\�ƷT��!�,P�z\?5G?�%�2mz_%��;�}Fy1��8_]�^�A}B�%X�~�4����&��& d�2���ˋ�ř��-�B��d�� �r��_F�H�ښH���me��>H��z��p��i�KlYH��� Z�����y�j۠ڳ��sj��r�V����U��e��>���Si�"k�j�	�ԨUKs�!�l,�EUl_U�����`��ϥ��m�b���-W�"dꕛ�e��'�e�A�����y� "���`���ԁ"ҙ�� ��s����Zg�/F�q&Jc�b!�e��\d���@i�7��a	����I+���a{�CP�e�DAk��^���(��� a�)~¸`�,�������G�����E����X�X�q��d�,fS��c`����3�ƎJ\1�sTa[�8*�@��G��r1a�6�,�6���pD_�L2_rɵ�;ަ��=G���`���ϴ��252}5.��?qz�+��d�w'��.�Z ,���Nw�~a���X��eoP��W�2���f�;{�-G��ӳ3*�FCY�e�*@�
'�����hop物#��J���c$�wd+Pts�O,���}�G������@�7r����\Jud����������MM�iD92}�Ʉ����{�=U�Gh:����QOȕ��J��9�V���%��ٗ+3��Jj?�#%G�a+�p�9����w_�Cu0t/.�r68c�Z�X����Ef���@�t@虺Ĳ,�󼭏�K4'.�ıv%��4}��^h�Vz����#��Sekst"p�)���.��HV���%%/�u��笡v��}�t*�l݄VǜN}��]\Ndo�@�HJ��vp��H^7����,u0�'K�1���r"*��
�!DY����W~ {ٱnzV�>��^D(�H|m�J���y:����;^�z|!�nV����5�mD�괩��y!c��1�>#d�AC���7u2չ���G�p0��4{YA�pS�F[�}���eղ����p��c�����.�f��z6ȟEQZ�'#��y��<t^�;�&L+��a���⡮�ξ��P7�C�=�'��@tW����gG�T���$����ryq&�I�kl���R�6eVʮ��ȁdE���ޔ�WՖ}c�l&,8s���dɭ�@Y��p�9(�X��(h°_yi4ySy�Ӹa�� �C�d7�A0����:\�K��5��Yq����9O�D?c���x�sՔb�V`-�0��A.yW7���2��_�gw�V�
˧��N��W���<�6
�a3��Xa����=����ϲ.��f�=��4".���}Ä�t�u~U���0P��&_}���3�\tc4�z�pf����6N$o�n@�)�Ͼ�������8s����G1s������̲fI��t!���.�L��[��@VU�܈���������꾱��� ]�����$�H-��j���6�]g�f�y9�o��L4,�[�ä�2�&1{�-iv�����:�䷕Ml_�{��F�3F�3�,�EQp���z�fl� ��mPC6m7{�93�5k�X��|��]W�����Z#m׀������k��2�ݕ�9k2��&��NIM�=��
�:ίt�.�H�G���6Sa�'�'#u���ڙI����"��5�YO�z��^Q��C����\}�����	���=A_������a���2[��F�K�ϖrr �I��ѫ����q��'4 ��$���Ϟ���~�������^�s���9b3�^?I��/̯\C��K�u�?�{1��2��5"�Ȟ[�:�J��@�����.#�w?�/�\^�\WЙ:.��X��`2��o�����ː�?
�T�� l�t9������^ҕ�Ʒ���ȷ���^%R8C:#5�=��YTg+�O��O���%���u�.h�\б�c���U�x��j	��_���sYnL
�AU����񡜬�2�,I�]bL���<�Sξb�Z�l���� �F�y���TЋd ������N����+a�A�?�3j�g�cG*1��2b�����z+�V��bQR�M����W;]Sd�O�&FN|jq�*l�D�ˉ{b�
_V�|��hO�倦�̥�7	'P�D����Gr1]pB�i��7j�r�"�,��/礒�{#�a!���R#Ը�T=�x�LfYP =�9�u9չ�H!�łH���|e0J�r#����$���8_ˎ��n�̎e�3�c��D-tŵ� ��d��������`g`�vx�~��Ξ,K�B@�H��M
k�����66�f�v����4�QJ�'uN���� �ɷ�<0�H�ua4��6$��#�F=�J�P�h��ڗ\�ɹ礞�J�J�N٣s�NE_�x��:�2@�`^��!���#��A��%T��d�t-b^�L�Q����ؠ�hl�V�rm�>�{��'�JAF޺��6c��J�S5TL�.K-�yjn�`�����]N�)@��u�X�j��[:&���l���+�r�3�*��||�y%�u��;ky��2ֱ�����u���,����=��gz�s�/��������ә�cu���4�Q`V:��Q����i@���(�����8*�"�[��s����jG�%f��*���P� %���h��]��w ���>�[�suAxϺf���y��1t�� ��6��8:�ϱDۺ{{��F��������}����`HY��iހ��<���\�>��d��<k ��)}�,p��p��1��q�Yw�<�H�b����r=�om2RRy��o��i������{H�^��(R�g_��z� ����]f����] ���>�Mp�\��R�l�ʳm�5>N|+�g-ۗ:��T�L}�l|�� D�M��o�x.��v�r��m�@@n|J��9��M���da~ 
�-9_Y_�R�,��������ǈ�9M(��<k����j�fP���Z%�B����ڙ��V5i̶؍ƠfT�,�Ƅ� l��t���`Ÿ�I���/z|U�m���[���_�|�ki����_�z���&�I�2����/�:��msY�|ʗzp/���9~�#��x�\8�I}�@��vw?���n��?��������wߑ��\f��\�5� ��*�N$��xV!DS�Z?+��c
����(^j�;j	�����÷~W�K��LP���b��L�kD�;g74����ߑ�^��ЗB�݁� �<���OH9���~-�߽+�Ҧ`��0�QA]R��QWƅ�ڞn⽞,���$R�`d���X7s�e!���*���D�~0ɽ��鐠�bogH'��q��̊�q&�gEJ�g��m�9'vD�7oo=���O[��jJF,V��{oZ�b�ڦ�,-8���M]T��3��^���C��ϻ������@E�5,�2z��y[ϮͣT�񜞟��l�����ܡɞ]���ߐۯ�a��u�(`��LZT��|)ONN�-��G1<Z\L�r�8�o�η��W���_���\���)(���9-6&���#�W���(�o��)�Rݫ2����'@��bn�5hpO+O���*(�`��&�QJ���Jz���}�`|�׏���޼yC�KV�s��8 �8����zQ��I]y���w`]@�t{���M�����Y�Ɍ�g�
���u0ө��ZH����\`��l�x^�H_1,�*�/�3��L�Y���]����#��D6�  ��T'D����$��v�� 
B.�h��c����	�h#�+�Zt8��
z(��(+�%KuH�z�gz]jA+�����v���tkOvn��L�
D'�����e�h&��=Y�Q��9[Ou�q�b$�B��(�j7�iX�]�J�ԑY$2��\�|"�PAҫ2��eq2����+`�.;lq�>��Gj7u>�M/����.�
({R^�Q�'��@�z2>ș�@�i��v�L���B����t(�.t|�m2zE����@��rhN��w�j�1*Rhh� ��e/�5�=]O-K���v�-bt
�)频5AU�h�~����W#��_GG��٘�ׂg\���ߍJ���	�y[�$�'��֪�E�7g���2����KuF1�*.�\�R���l��|������Z׽�i����Cl�Z��[y]�4`֏�|�k��(��5�������2g�UɬX�Bv��^�)[#%�iP�d�	&mc�������.��4�c�)�cϜ�
��`S��s���#}�-y��P:�F��g���Ӛ�PP4v�wlQ���Pmcw��Ї���\=�B\�������&k��P�W���3P͓Bz�%�9l��7��<���V>�Uwc�Ň�i͈W��_�X�����1O�qmM� ��U/[���=���I�g���i�{��e���
��RK���v���u�߇/�9�0��i��"ħ��h��"���,u��^.{�D޹��\���_������r,ߌ���NCd&e&C�/-ȍ%$�|�;��v��	]d�~��|(O//euMD�Y��_�C�����\�9p"Ԁ-g39=;���3�����>��'O���)�5�8����e
 �zb��V��b#+�L5ct*Q"��N&�o˙�J����R��I䥩�¦������2@EO�A��`� ��^��z�)�e�r{8f_�XG
�/�4���t"/K�]@��j��(YB��i�J��2��ؓ�@6R�<ø%m6�$[C��?����f&���T5J��K��#�ܦP\T�L�b���{t���ّ�'O���wdww_�ݿG�����3��2�kG��ӧOIE4�p02�;�֏�������'e���T�&�R7Md e�V�
,'G7u^��Z���+k�ࠜ6*8����f^��Z`BCȆ�)p����rN0U�o	�X�6�ݏ>��w�&J��fI����=Y+P8;=S���f����y�
Z����X��\Do�˨�#�pƹ�����sJ�����)�f�fb���Z�������׎�Za�H�rXN.uL�z�}\��̦�x�u�����x���R�OΤ��_?P���_�k�d�G0h��Y���=}_��J��̍�����C��X˖]���uGϭk�����X�^`;��3uP�A�O&�P��読��)!Z�4E����
�;��4P���p�����C�:7�bW�N�F4l���]l���D��^�a��}��r��W�Z���KqcO��w�T&�����Od��My�z!�d%ᰠ �(�X]�xM �rI
��k5�b��=d�k��+���w<Z�������;V�c�C�{n̒�?�Q��� ���^K�^f+S�5S�����捺{kC��L%Ӌ����w]���Ui�l�g��qj����H��=��F����lZ��i`Y �ޝ���?�b��8��s�J �&��u'sR�bӗm$?[���O����'ׁ��x�l�\��3
J�뺹��,����il�
~��ߛ:���g�/�>G{��#�C�L�����3͢�Pe��%�^)�;��i�#�̘�6�bf��fν��W��p���cc	^��Ki����]=�<gx�ڗ��t\'j��0�6�A��T��Ή(+�
��C�hG�>��p�3���jh-'2��P\/X�95��W���ڎvX�D�J�`1g�*�ˢ��D��Z���������j���i�⢐�X�8۵��i�6��g�D��F!��~�D��Xw�u?����k�������.��9���\�kz�*��{�Y«�����V^~�/o�����p������R6��8�cG�~�לE�ud��×V�4R���_e�����Rk.\�0�1>�,-��>p���� �׿��<R��
Z�A�i'����;oC�YOn�:�fG�U���ш�B 03��ꤪ���1�零�Z)�;��!�K��@��tE��TyO$(�uQ}�Ѣ�ԁ$޻��i�lA%�b`]M4����z�1�"�qFԸuL�ցk����68Ac�vW��/3"E�u��y��T*�OԛQ5������~��i��&�yd1���W�|x��7U~���6[l�7akpc@#x{ +?s�A��̥�1o�>y�w(=0a7�SG�o�����r����M���A��/�˙ =�����������"*�w�/�����ʬ.e�@rU�xE!���R/�����L�ӱ����G���d���-6C�-QZ�H��(�+(��aV���Vn(~�Z�9�j>��dJ����o]o�./N-��<B�-d,�̩CbA�NR8�Ii`t�k�#]�a�x��j�\{�V��-6�A,ӞfV�^�s	)���1��L�:x���wO�K_�B5ȼ��"("�E���D_V�g,s=OV��OJ;����_J�eͬg`q����Α��Ԡ���:���P{���BQG���a���\Jq8��Z���@j8�:�z
Z�D���X�����z���g��R���3ɦ�\��zC(��酪�����J��ٌ�����#�W8�4�GOB �@V���e)�󅎅���<�lt��y��Z c?�q��f�u>���N�5?��_�O�T@��gt���t,AQ�Z�(��B�Xb��+Ucb $�1:��fQu3f�|}gT
�A�"=>Y����9�6)ve�u��8R������S�fȥ*��[���֔�=�h��f�aI��cC(���q��C��R㹌^��Aͣx�SC��!�c�;�&�
�-!,�ി���mk��F:}�$�����w��f�zy?G�Z�������:� G�Xb"%�d~_������<�\���q��=��IS����[+ߩTyO ���!�ņ�	{���ci�c����ob�b�����<f=#�	��^�*F�Pj��~ry�D��{:Y�y��ͣ����
;�!3��P 7������{:(��2萡T�>@d�l�D�R�&(s�ZP�D{	wn�j����L�_I�;`	Ѯ�c�ɩ���9C>�y�b��q��6��ĝ�5]o'�UM�W�\�o=��v�F頟�T�z���"k�1�P�E����w�v���e��v�m��L����yo����w9�~J����wh9��u���B�}����<mm��3JiL�^Lq3���2��2����Ixʍ/��P�3�����JԈ�
�����uꜨ���1�o�P#R��~�8�pĭbHJh�hdI�~ 2C���QG}U�S�¹�{�����jh53��:�C�ɲ@`�{G�V�Z��"�WB��@�[�@G�����ʭ;���gmE�Ag�q>�K��[V�����qN:�]7�2_�� �>���颍���c�:$3�eFRo�kb�� �i�B"�[J*FO����T���%�`�$��ٜI� \�-��� k�}÷G}��@=!nJ��O��Wq1��W�^j��e�B�F#	[e/r�������9c��M�7,��c3J����\4�=
��R�wߓ;7^��᎜_<�]����/�{�ͭp��?���x�X&
��\>|$�G���%��1�u7�I�&o做Үz6!�x��H����5�A�ٌ���_�Z�un�J_��񑂈��z]����6x�:7�u���LЭ �4�2��f��W��^�f/���lI��?p��:t땾�M�i9��
����$
 "���t�B8�rj[���-5� HF*��>���+2�"M!����@��\��C��J樂��Ӹ�@z�,�(x��ᙞg�k��Ynmf�J�l�"<B�u#=�)+�H��<8YK~��ZN�+�7$�9Rp�2'
��Tzz�ٚt��i�p	��_E�A3+��I8ʲ�I���5�*h�����ְ'���j�
lu�ww�$;F���Lt����L����}�O0 !�l�vj�f�ʥ�-e=�y��L��d���Hm1Z��3�Ηrp���Փ�c� ��3�گ�|��D�O������zGP�Ef�o��@7�-.;�p"�[���{B�|Q��ϰ��H"�(��u�YA-�l�ϡ�z*3+܋
*X���{d�0��|�N�J�E�9���)��U#y��#q������c�w0����YϠ���΁qT�N���;�5O_a¥p�a]̲#�L,��|}#��$MM��N͞�\�{"m����x1X�ה�uu���Vp k���D��w��h{��Q/+2��1k^b$��Y̓2�\}��4�p� ]���4s%s b5u �[x ,z��˂�d��u��]CvО�}F%1�0�E(�!˯�s	�01���q��zQ
�R���{� ���h;�������0��?�$j�t������/-�T]N�sk�0>J�Qĵ���j�{��U���� e���K�������\�$�z߿��'��&�u:�':�^�u��c.J_�c��;�.T��v)M����Q�z˻�]���Un��3L#0�z.$UY��&H�`�@����6��f�7`�}������4S��&�����m�a���NPh��ے��_p�+�<�����B~�Ǘ��~V3���eM�r[DO�!��bR3��R�����4��Q�2�|�����ϡ��K�����Q���ȕ�D.d|r";:��pfc�y�@fp��Suf��W��S��j*����IwoH
��]�r�����{R����q�%�l�����f��� ,�7+5R�L�2ڿ	zc����@���h��=2&��W�M��8�o7�^�Q���7�^�e*������Y�1�j!N�~y����ra����Tn�r�5��O���tw�F	B�ʌi8X�XU�i2�8ݨ%MP�l�D��8�*, �o�^Bp%�ɣ2��!����#��T�A����Ed�����H��'R.u�:4-.�Ą���`%��"�K�"��R�l<*:Fo�M�r~v"����R�v�u�=������~�Mݰ:��y�G�=WMt!��\�us�n*���Ǐ���13����~*��ɤ�� �����X��4Bi�h|~� ��������]Y���&aO�5j++�?8�����o������x]~����Wo*��m���r�\����?��yx�T�.p� �zh �)&D���ң���K�G�nB��u|�Q�:X� D�5 h�ևs��T7�cfjp��tcaa�lB���k��S�YB���k�`Y�45��o�%�=��g������&�?8yx�L2�l��Y��1g7�J�"�b�S�!ʬ�\(v�2��K���WV]�������;ܗ�P?��U��Νb��d�slUIy���H�p 56ECd_AC�ٿu� z\Ϥ7*����}7޾!��N�J�zх~��������g"�:�����:*zϠ0U�c���:��Ĝ؎9>W�~��O�*X��Y���f������_?TVRKv -K����v�)�+�<�b.�xu�!(L �=eYG-�IVY`*�5r��� F�t>v�i����IE�U @��f��w%��q��m/�-&�e�@�E�S���T'�H3f�����KP��W\Km�=�W�Uo}Ϝ�bΧ�,w�Sw�C]r|�9-R�G�r�nb%��yb-�6�v���"���*1�/��8�'��{T6͊��@�*n�_�M#�lq<���+n�[l�w�c��q��G_T����[�CFͧ�����1�����=J|2W�
��������d4�����G{u{8�a�ԁ��Y�����t��ˣ�jQ�G���k���U��>ZW��c��$��3�9����ծ���%R�ULP� =kV�v�1�����I�L&��2
�A�!�)�(��5Q����Q�:R{R���_)O��/�ג?�Chs:�?�2�.�6���阀��#��idÉ�"�Ic@f;����/�ܯ�K�:����v|t^8�3q(��h����E੎����=�o>[�u��}vڬ�\���6ּ��g a�S�L�H�h���i��O�Y�p�������Gf�Wq|��Y�����Oؘ�a�2�e�h�P�
P|_f�~:k�x���ک�>^�z
d 33�uT����tn�[ߡ��;�/u�6jX�޸#?�����n�fo�{��{���'OQjT�x�^����o�!��L���?�SCŔ� 
L�N�¡���I�#cP�Oͣ�2ܗ�ވc��F��Y8@��� K�gA�{�|[^OG�zx"�.�٦c�^�N���p��+��]Y/��l��Jm�|�"���t����o�%G7o�;���:vK�Tf�2B�T���w�Q�V��y�Ϸ��c&s�j���%K�"���I����a\��>���z��<����f���&X�N#+���^D��Pb�v���!z�U�¨��o��
|6:��'�L�
'����dݭ�r������T��sֽܼy,�=��\��[����H�QW>|p_�R�M��'O��w?�_~�>�D�7���2�{̮#c���� ߐ7^{]�>~�ހ���:���|��h���_��_�����͛�o�%o��:ۖLgRD������w�+ݤ��L..&�
=F�/dK��a�Ջ5����"��fڳ:V�rpLs�T��)E��"�4��b,�׎��[R4!�d�S���ºj�k�m�]�2DQ�;��[D6�]���ދ�1���P�e� BG=P�
��"�:F2�>����,O.u�_\XW��KZ�ZV�g�s(��6��GY3�F)U�+�+����֍rE-^F��"�)�IA�o���)(@S��9�n�[�ds2�MQ��T�Qc� ��˧c�wr��w�Q�e�A_G��ɦ��$�n��A�h��e��:`����\?g!�dɖ*���ޥ�|UP ��a�S�ٓ�����8[������Y��1�|?8c�ND��̒	�| R�H���z�e��n���׉�5!�>.�-޺V��~lqt�H�E�.�ri�H�VG�p�����p���Ik�[-��D6&`�qs�Y��-(t�E�ֻ�cQa�e^��C7���2��vB`����Fa�ϑ�Զ�-� Q3�UV��"i����XR���R��$�����w!{4����Z\qc�54W��<��if5�d? ����Ef�ϩ�b+ج����
bJ�f1�@�ρ�`E��:q�$�3�bc�����������qؐ����QL1�"�I������@l7���.��O���&h�=Sf���t�s�����L�,K,q�k���q#'�\puRKl��i��G�S*�0KM�Df���dH�PD�\�:ulCDڨ�|�թԙ�]�����?�m_�en�g`y��/9sDHW��c�7�x���`0��ԞU��i�flW�[�HQ�'��lΛ�*@U��*�Y��e�*�q]$W��gN�3�_��-��������#E��m$�
�lR��n c�+��8�5��-B�V�BB���g
���ȿ���F�CbM���2]��}�k�?~���/>�@��t��(�
w�۷�mu��?�9j�2�|�+��3ߌs��kR�"���(eqg}�%��I��3u ��6�<��� ��WՁC/�Z�W^C��_��ə�3���f
O���b5�R���S9Q�1Q��lr)�N�2Kt�?�1�T���Y���K�@O�酼V�����s�Fg"���Jm�ö}ƶ�z�4��H��3k�������o��QB�f�����캊����h�&��?9��$��"PP�i�4!liɈ@wS���Z��\7*����R�9Oeo��N�J��ݿ��G:��[���:\k~M@�U��x:���(D�������僻1X���d��9��� ��M�M�������[W7���	4*����y��HeE�H��ۯ�)�������G?�����L������y��$������򞮙��SnL�޼#����_����G���]�b�&\��Z�
���-٪AHCF]����0vH�)�S�I_7��_�-��uY��������2B��Yte�� S^��Rd�^(M�
v��:Ǭ-
��qQ��)o��lCd��G�A�-�B,i4Cl�a��wQ�^1���.�� r2��BV��R�3�����j?�k�d�דjґ��Q�;(a�w%핤@S�Q4�L�l����\�{v��_��Av��^K-�'��twexc s�Av}g ���wX�����I��S�'�t��zσ�Y:��	��C{�<a���rƱ�#�;Y��ñ�=�*���
�!׎@�م5�F�ʱpa��P�\b�'�60��� %ՕA���vkv�ΰ�C�,��'D@�rP���1>���ʞ#D|����6I�
6I����`tuN�&ML~k�^�'���q(?���8bWZ)������G��VV0ı
~��_������ڂ�!���F��p$sBT	q0�0��2�4���3��\'��,��=���ZpTF�����Z�~C��k[ǞB5��mOa�`{P3n���f
�^�ֹ���I�(�6+�
g�{Ue��P��l
��i��n 0�40Ӵ9o�2��g��|Ant�Vq-��묨0^A!VB�|�6�kJ�xOd�J�	P"v�C�f�	-���	v	S�=(�f�5�H�@��?�<L�~�[��ڍ�(kN����c�����||hMQ�H]%֙3*�G
zӒy��i���V�ַ�o��:u���]�t����������~fp6�x '�ng���L���k3�9QUx��F�;��x[������CS���k|��[??�zI~f~����v��.>`�)&"�rشE).mM:�!O=�y�����S��:�/�	
;����nX+u��������8��́�����yOV�R�./�O?���!?}�e�SC�=�$N<��<�s�:Y#u��7�(DX���k�z��&plĎu�����U0��8�^��ť�;~*�>�	��:�l*���6���9)���ߗ�:���;z�%���͔�P�S��5��<+z�SR�v�_��PpC�t4��S����S頧�~&ˎ� �+T�,-ր����M��Yi@a4����u��G44[���0S���Y�.��ut-j���9�s�"g���4^G!W�+kLl?7�\�	�R*��pN�3��3d]�p_zG��w�Y��'�S
�:C^�z����c���K}��x�~��\^(8�#�ۥ>k��������R�JBɕ���R�a]�|:c�C�Gw��O���d����uW���������o�΍�����p�X~��Y�g�r9���R�W�έ��|������2@��E�Ќ}'���hWv���ٜװ��+o�qM�����ޮ�:WǗ�,���8c{�[l�ѹ��M|����y={p��~Gҝ�톱L�� xL �u>�2��UEg�u�'i���u���
�ˮtC]Kg�sF�r��/��^�z�x�V�l.���Zx�6T2<ޓ��Y�f��K*H^���.R䗝ZV]��ve>;a�a�G��Z�JO/��:�a�Y�5�����I+�DF{9|eלx���{���Lv�w��D�*�կ�_[}.[ ) �GS}fk�:�w��l��@K"$��-X�J�.������ɻ%����5�|��p�+����s��S��͒\ו�>�Y�\���	P�%�F�����ϼ��3�F1�DR"A¶��ז��4o���ɪ{�� @IA⢯)�y�>{m��lÌ'ě�g/A���C>�q�y��d27�V�J��~�\��K�7���D����+#����@A�RR��v�X�{mx�ҩ��E��ߴ�:���̼m�OF�4�4Js�1& G�#��\%-;֮9V�@,S]E{��):���G}���@k�c_�y�_���cdn��^{�/ʬ��E&��%�}e�6�^[��k?�K.j�o�,i�e7�cЦ�'*���(�����ȓ#�p��
$�s����v�<|����9�'$�)�����p_��{W����++� �Ydwe]��LPf苕5<+�$��{]�ʘ5��M�yf!��RJ�i������j2ם�	��V
h��{�2��0ȝ9D�Ii�Jܯ������d?k���v.-4��N=��ȇI� �Sev�Zk�n�6�^� W�s��>�b�^�b�ȯ7l��� �ˀa����yh�i8�|��45���3d�@zW�m�����7�>4[�[��l+�RT�ʱ�O,]�,�_�4Z��7���B� _�a�����1�?�N��o�4@!�45�!46Ac��F�C���Dz|c,�4�����7 ��|.�����?�X~p�r����qp$�nO担��.�ן��|r�XV5 �.��V����������z���x�N>J��&Ӣ��ۃ�P���F���`��t� �N�!>)�r�@��lj�G��v.�� ru.O���,׫�]\�M[���H�^���d#s�]rx(���<����T�{9{!W�3fn�n�w�ܕ���/ԉT�'�!%��sy�,�4Le����L�>���UR^��u��:"��i�p�IS�e�T�8��_r��� ��*�r��ړ�^�N�ef� ��.[ JA6�f��e���K�X�$�ޥI���J��F����٭^LXNE������	ųQ�<)V�U���sM���MY4�}X��X�^�QG}�Z��bt�@���^)X8�<��rFÍf�����ͅ<�=g/���z8Z�?S������W3B‴	��p�'G�5V@xp�m9��w������?6q�N�,�Cx{	�o��_�R~��?�D��뵼qx,դf�t	�Q���:я�@�)YYЎ��u����]���\bϒ�Ix�Թڋ�Kӟ�쪗��|Ό�%��z�(���M(���D��T ��b�}Wg`o ՛�R�ѱ�X�r^�dt��%m�H���T��:9�@��֚(��桢��%q��'I���YO��c쀤�.��w$L�$�7E�2�

2a4�-gW�2��폇R* ]�0f�l��ǚ`|s������{CYl�,2_�t�S�=��4��`(��oI�W˼3W U��*/�#�&H���M7����QV�(�Qj1�UЁ�]����jù�|��C�R!��u֌�C�} �ͥ#�7HS�{/������'d�LXG�s�4Q�,�X�
��?@$�-�ڝԒ}r�܄���zZ���,��#l����)�j�5���m��Yl��a��q[G�/1ChA[/5� ��n��
}�m����=�D�v�QcEQ�NtM2�����e��$>N%לe�)kɶ�����v���wKk���+����v��3�v2��y� {�t�ǂ���G�6�Ij�&(!_7e�_���HHg��[£�Mv�֞�,��נ��p��:�%�Y>;jk�]��P�/����4�Bdi���v@��ʿ"�J��й*��m_V��� �V��L���bϙ�WE�D�俰2fB�`�� /~��0x��lA���`�!�v��uCfe��/d�^�^�!�c7�$�/+O*@'��,��� :���|����'8@؇�;::�.*h���@A���{�\�DHˈo�Ƕ�ʂ/�ȗ�:����KXF�z��2$_�%�
��v�{�|�6 �Eޱ�O\��7�-���i2�c�b�q0�s��������,�}B����19�,�?�����ߑ�5�u0Q~�V�g�7�i�3j�������>�_>���m��ܢT����Zd;D9^s������?D��Ot6l�Br�	�P���R*��`)�}��
��j�f �����Vn��<�s2�],Wr�O%W [I.�:�pp���Ӌj�m�e�J�N�F�{���i� ����r��|͠��4�P�4e�Vra�(���A��%��/���,^\*���5����[��ؿ���k���C�5to�}�c)��$�}Y�c�C�+�S�6�R>��(��,����?�T�So����9o��?W��յ�P�YHR*���JK�|�7����JA �
�A(d�i��4�p4� � ��z$�K=�A�1 ����Q���l���0#�I�p��]s��NO�޺#��]�Kz���]:�}�<}��r(�up,�
���w�����?�o}�9�ߧ&{��� 98+u�^M.0��l�c��H��7۬j�L�Xʆ,�F� � �6՚��`	����k����\�S�ڝu����V��G�4=��9�Q�k!�ué*xZ��w�}N�b���a��.W���"b���suT�c��Rd
�L�k�=��ݰ�IG��ұ����V�u�z��d+����<�~.��BJ���r��h�2Lؐ6J+A@�\�>W�4V�y�@zw�e6��|:��;")�勹tQʺ]�5�;�'3	s=讂䗺� �+��H�hm�.�X��2js����{YV��a@I����uUgȴ��A=й�<G0��/�����5Ic+=EX�4�������%�%�j�{����x�f�]
�d6*��z.k�:�X.uM)���)d)1�_�Ks˔r�*�k��22�h^�0��?��_��Հ�z���u2�d'��=`}ſ̱��6�0����g��k9w�c����A��>�$p0Xf��s�v�S�gӎL�sfQ��ȭ���0�Bf�ndb��A��j~�FV��Y�'d�j��|�@/�f�Ś��@{&����׹g����%(k��Z��gZ�<�
�`[V�ܖ͛��H� :�� �����[�ߠ�DK�b
��|�������|���ޮv֒��!�����P'�Ov�����ꭔ�.0��I�A2pHR-�� 3J�ѷl��>svz��}���J�}��^�3��{ɨm��l^���jp�����G��'�'Ԑ�B)/ؼ�.�dv5���y��xqfDC������;�~���e�6,�@�Wm ��d��П��6�I\j����M@hV2���bH�e��1P"����������[F���14�a��ƪM��ub��m��ף���t��ľ�CdY73D]
R��yȐ-�I�&5���}+9ķ��}^0���l���.�tޭe�hc�=)�$1�O� lc���jj��Gr� .-���C�n���6K1m.Ht0�	k��0+TT�ZfK�ƣrZfD��jhg�Է[)7�1��+Z�O���"��T��I1g?^W��'WWr~9����k�|��5�Ú)i���$^��8y9����)�b�%l���c���0j�C��Bz/,3`�iV[_Yd�9�$hX�P�6���Sh"�+²x��{��)hC�� E�4����J��0l 2��mm����s�����G���^<�Ǘ2��u��QW.ʕ���P� I|�֘��M�<K�ٺ�����������̱�}��=�~Z�T
J�3�b��(�\g5��d1�ark�'���r ��{<����SR�d=!c�o�+�*�)���ݣ������s���ǒ���P�ݺ-?����G?���z=f"�ӳ�O���D�>{&O�=�G��7�u���3�F&�����gR��+��
�q} ?2����%�S�>��q3�E~� � �Yj����b�i(���]�똫�@��A_���z��R�kݫ
�ciGy�������fcz|({�C�SǦב,Oeru.�|,W�f.�?��ɹt祌���Ks���DbR�z�DA��!��@p��IWy�&�+��l�s�_����P�L�ld	��~W�p[=���t*�Dmź��J���R�$�DzyKZ{=s�0;՜Y�JǦ8W��F
��$�x$��.t�Қ���/b�ƣ�L�)�\L�R���[�C������%��W�%����B�b������%��%q�?c� B
:���%�s�ҫ]U�ժdpo�q[D`=L�i�A�22j�9�HtĲ��k������J#�}��w���� nO����kB|�6��O�@[�'�:��돗��u�Z��_I�K��'x�U�l32��A�Kj9;��%XJp|	Пj����h\�+�dv�{�s~��3�!bb-I�]��u�-K.D3Q����`��%��Y���'��T�-8�cܫRt$4��}�l�gSo!oܻ���-�/��Pg�۶^3�A�V��e�&O��I�[5Ab�<�&�1�̟��ڊ�m��'l}�f$�S�y�H�$�A�g|�U*�S�H�L��#i Z��ȎeM��'�D�j�U�-�}�\_;�	���y�`���u�-��~�4=ܩ�x�j5-S,d
�Vr��=�{ru>���RN��ȧ��D�<yJ��A���{I���z��ۡ_[����/d>.^L�;��c�K�>:dJ�{C�2[̤���ڂ��'Q��4�D�w� [����W_P�n��v�|0�5-��?Q�f�����]xu������|��e�&�Ӂ��%�M��*�iS'*��B�͑*Κ���O�-V�'�t�x��2pf��1LBט��۞E�"��^
�SZܶ��7֨_�ܟlt��vSsё|έ����K�B��������2d�ѵ� ����0L��/ ̡��pS�M�-'4n��gu���j�BUd�2KA3��Ibezp�� 4�xa+��C��o^�Y!��q70�>G��M�<�*�e�M7*+{á�k+D���g���!���O>���H�3�y���@f�XAp�X����ŀ����Ny�r��Ɇ
����mύ_[��7ߒ�|�=XK�|z!�
\�q_��2��˙Q��t@�me���e��������Pn�����j{�x:��
t����̈́�.BÚ�{����FC�340�������='�W��{o�����kw8��O_�g�Oe��3[��~�o̷z��}9��gO�f�"��m�m�r����Ǐ�ѣG�_�Z�H�}.S5Γ��{þe=�� ��p7��Qc]1�}�����-��,�Ğ��:s�ӐPǪ	��� ľ��ˀ� [<�y�F3��fp��J�@k��z�
c|[B��V�t�te3P{4�	4�ץ	�U�k�Jȃ��e�j3.�2]M�V8�Vd��D�/^�R�|6�6�EG]}/G��9"谿?���M9�0�k�/%���|.������4��RG0��|9���w	�V!�k�sOn���B�^�BW�Yd��I�R* ]�&
�+�+�$�x�{ 9ѲX�P�U� ��֣��Ό}u�vL��۵�j[��ֹ��"��:ީK�l���ie���##��dӑ�u)�rE[� L:��F3��u��"3Xq�6�ͫb%ü�>�dm�s����,�EfM�Sp�"|ph�/ӄ�WP�����G��y��=���[���h�5��WB�CTV��o��Ia?G �s��'�?vX�__�w���[���j����=��hlP��X�$�ٱ׻���溝$�Xr�J#�� 9ȜB�` �(l쮉��Zϡ���3�f?^-[���� �Z��5DL�afS ���Y�Y[&t���rr�\R=F��@����\Z�F�ն���й�UW��6��Df>�Xа�6G*F#S7u#qtl9��S�>�G��+f-��x6z�&�w{Е�)�5&�&Em 4dMF�U��Xz�;�,2/g��(�n�G�Z����K�@�Wx�Q���̪8�����F;�����4̇��,/���ڋ���6�Q:f�?��յ�����x��(�}��cڒ�ON��>���=������,x�"x|�p_�����k<��X�����9o밴8m쭄�ͳmY�?���'���=�}�X���a9�����R���	�f�z���k��ߵ�x	�L(�+?��#P7M��LX̹��(y��k�r/i�}�ב�y���Ohn;F!c�����N��dQ��^�
�p4H4�
B�:�=] =u�::;pΐ�a�_e�$�p�;D�7^C#�O�(�a��iY�u��|"t,7��S���jD��K��T^���%VMj�(e<��N��!y�Xٵ�a����2��-�-@�k�Ed������ě�m�j��ۤ�"�0^p���L�����ǟ����
��������
���1o0��\AG�"�:�d�D#?�4����F^����y]x��� t��}���I@G�$�qf.�d�.~x����D��sJ��� �r\3��y0�	K�$���@�}�2��#��J���%D�Y?�_�߸+�g�ؘN����5V[�fBE��Ƅr	�@$�F�,ƐS��d�̀ �����d]9h� F�'8��/�Z�����=T`v�7fo�	[��������F>��e�s�V`��Ɉ�t�Tж�����������L������A��?���{󞼩��`��H��CA�N��}!
���3��~���z���3y��!#v����*���zq~"/T�хY�헂E4�B����|{��?!9�~�`쉏�Ս���^���㿵٭�A�k��1�[�|d0{�s��I�a|��#0���=���}�6�`\/�vWrD&AJ'�_���~���Q�<^���X���s��$�>2�X�O�k'���+�ө~]��zO)����v�%{�K�ց̟����S�x&KaYe� oQ��tg$�}+��o�U:�
n����T�K��钕������ Sh�E�\E`�$ߘ��ԍ=-]N7
L�_����3Ԓ��۹�(��Mf�Uʉ�:�K���6�76k'��������a�h?0�J���U�Le��\��BoQl����"ӍH 3E���Tւ�r]dU�����v����n�EAyw�j'9x���ep�u������P����[""�����M���y��4��۾���@��/���2���K<)��Q�["$��THYK�%��t�;�L�̬��ds&K�ߦ10�Y����CdE)�>*V�X�t�W��'�(S��
�~ʦ\�����8��n���V�u������Ǔr�-���{�K��N֧��)]w:XV�ڎ�c(��~��r*���IO�S�����s��{`mhj؛� j�#X2М���B���� �'ɵv��}�����_�#�x⺲
0#-�4޿��,�|�Z�d�gv�ӷϦ�WM�,��=�܎�u�����M�^i�r:pj�ѸVf�_+�0��b���7ƀB]����W��e[��r_߇`�4 z u,����'��|(��@�W�S��y`���y��V����� ��قㄬb��i"�C����~A�Փ����������������oJ���>K��@i=��c���f?Í��5@���
�LF�>�A��~b��U��&���R'������/���[�y���/��~�7~|�A��|���x��erP����W	R
�ק��2O�q��jus1Wx�T��z	:K)�8u�o\e��9�Mv��|�Ѕ,]01x�Ղ͡}�ϵG��I�n���:��1zS�1$L��%j.�a�~]��l5�r�+��L�I��P:�(Z��g ��������?�g��;�H��2Kj�yDϘ'0B���n�r�V��=���x�jc:�b"��B�`[��+�#�n�nڒ�t%��A�0�u(}_%��ZZ���
��G�r���X���#�^��ܽu[����!�������� �g}����J��� �U)�����";6"����\�+����lͲ@�BI�R{�����J!V{�b�;P05�QHÉ� i������D�Ϧ3[��e2Md��h�|�iu��z��ܻ}G�
2>�����-��]A#��[�s������o���C���S=��
v�?�\��'���y���W 7�;w��t���^\ʱqZ�j�zrzy.���7�B��Ʒ�%W'���:o߻�{{�챴�՗�U�s�ِ�%��,��Z�^�|:޽�%��,mX��%�`�1B��ğS�� pC��G�ua���w�끎]k�R/@k�܈���p��K+S����@&��nW-\�>ͮࡂ̅�.���'�{��]�t��2z�Pz���we�ZH>-��ޓ���t�% W��3�!��$�b� �I;z3�ч8��R��b�K��)�r��T�zS���Z��:T�U���?Py��r�� �|���a	Je�|�E.e�뽓P���<=d�'�gÔbΠwgO�`mut�[$�)�sY��}��z}
�zFT���������wv"�^Yu�r�z��zi'�]�=@;�2sTЖy�WU����Y7�J���˙�{�:h !2��I�:)[��x+AR8K�mD�GD�O���=���G��?'����`�'��u�;h*Y���"�Rw>h�ǎ�F�V�˱�L�uE�Yo�J<��s�ױ�_�"/?���gk����ʳ!赮I�2-s���Y�C�d��u�*�,-k���o�k�g ��6�|#p?�m �:YmQ��ŸR1I��l��'��r� �qd$���ڢ����FN$|�\7�+2`ػ��*vK�����5�▪�AAÈ<s{����2����Y�{�`}��8��M���M�_j�BB�(I���b��=��lf����Rt�b�a3A��W���m�c=�N��2�(3T�`+�l	�x�"�:�V�q��V]Te�u��;���s�2��ͫ���W�*:�|�d��yUo��}�h��dd��@}��Ǐ�?���$�K?|K��/;<8$ �?�#|=$�]��c�_�	N0&�'k�k޹��|��oe������/���~�r����-]{<����7_���t�2��z�k�,����W���T��k�R/���_���xs�dݺ/1��ىks��7������%�k����M�l�+��%����BE�]�[�e�|yC-I�꾢)+w�<M���z�^rOb�7��{��em�B���&�����X�<j�񩼡�q��f�^�+��	Kv�e�*���*��
�;��M��#�1=��f�9��Uf�(mA-��<9����'�>6���l�^Q穭�QO��w|G�z���O�Siz,y(��	���l��DԑX\�g:0#R��C �~��L��l�U��$�E͒�2ZD��t��7))��C0ST�
V�̡�r5�u��o6}�L食	b��ց�%�9=qN���.1����L�^�R��C�V���Z5�HA@XZ��GY���v��&?������#�~L��H�.z`�o�}E�C��9[�p��5,_N�ip�D>�����A\�����Tu}1 �G�C���CG�.����#ۢ�n��"i"�6�+ "���w���rpx�l�������� ��7ߔ��g4>O>�G���~�+��>;}N��v��_ s �,e��j���B�0����l��>�DF|�ЏN�v�Ց�C�f	�Md������l蜞<~.ϗ3)�C�jE���>v���K$AԒ�����OH�6�wd&t�.���/t��@�P����H�֞<�d�+e��(������g8r�I��A����6ےB�d�;����F{�&�[�^����^�Z>�Iv��e�)�k���Nu����Y)(\��=�1#�œ+	gkB(�NL��2&���r��U;� �B�93��
r��pȶ���m���1��a��@R5c��B�K�H�o<T`�gV9_,u.��>]�K�n�Ô0Ï5��v_���!���<95ǿ��y��)�H[F��H�R��� Y�	�cooE�KF����u��9��k��
}��E��s�������L
;t�1Zh=C�3.P�ҽ2���ݿG0���lM�m�Y��m�yK¦6W����W�3�#�u7!�m�W�ϙ�5�b_��1��ɤ���Po��Ce�A�4IY	*�d4��݃7���P��*m�SB4������m]�B+m�n��f;�)���ֲ&$ok@����nw�:�ַy���5�����U�[@Z�FŐ�?0�E0��>�ŕ�B�	������w�������=�����T
$��qw�[���Z3,0k�B\f���7'��S9�2��Uh�v����-�s�]�f�㠑i�
��zt�B.��d�I�n�Bχ<5�Ǥ������l�-�g%����!�;����#v��q�n#�KDc�mb��H�([���͗y�_2�1�m�����+��\�5zC�܇��/�<���1޾�6}����,�#��YZ1��2�u��m'�(����F%�1�Y0��@ϙ�̖S���G˓~Œ�w��-#��/����K������aK�s-Cn ¤沉%�f�_aG��wnw� ����e��ȼ,=�D^��HH4��Q*���k�˂��K�q��9r�S�v:6�u�Xm]T� n�������~��2J��g��m��-�
�=E#�R��Hw& �M�~����������N#23�Z�	�����j���<�6�n ��o�l%�QۗI��YQ�Y<6Y��D�5+WOTjL
>�v��X0���NX�?����ϩ��t�B����P���C5�^j��`K��.���U�� ����i��x���Q��W$z��tf�
��0��U-^�as���G62�i���g�>��r"W�Z��-�2=y,�"#�l,��S���h���tA9�F���M�S��B��U^"
�ĸ�tN�ĸ�N�@����;p�;H�����޾���.0B�ZVtN��`G�����m4^�lb֌G��#�~�@?�h<"�P��{j4ѓP1�e=]��*@���D>}@
��Ϟ=�����{���g����'4�`
�ٷ`���|� i��} ��=�>�ӧ����^��o����R޾s��r%�=�yz����)����\���Ѵ-�˩�������U�h����f�b�)��l�����j��m�.[�0��[�}t .<#T���f0��`6۴-��+�c�� 	�"�zSoH ��������Jy^]��e��H�;C9O�%�>ؗq/�a�������i�`�,3FG��p��mM"!�:>=�C
��&=A���Z��Z׼�+$6 ���l[���|f�m�����<5� ȥ#�j������g�g}�
�k����is1W�I{S{��F��BAiW��5�6ݲ+�'�2n�JV�BZ{ڂ~Ց��H�s��I�k	.�}x.�w:2U2����A?kqN�:gv��R$����6Q�~Ւ�́�0���ZEBA�d�t�#���6(cF��}nGQd��"�8��Sf
+]��Ē���Gg;�Z"QZ��y[�S�HC���w<<D�u_8����~��TQ��,���i�s�4�Οﷶ�v�E<���ǫY���/��f��<�jq���� 1SZ7�?!MY�]`�!ݦXf�����a_M���ݞR{9�Hl?0)�P8�67����$��[;��s�%ɥ�?�e��z�,P}">dh��ӱO�H�{Ƅ��x���Զ�V ����2��Q?v��P�f���J�,�D���5�R�^��z��H�{���Ę�9 ۆ��R܍��j�d�
�Xgf���V+|K����/,��v2fе�ۉ̑�n[�CZ�k�ߗ0~c�TsΛA��Y�H,�(>����4���4���r[��rjZ�vؗL�u0�\�Ĭ���v���������|���r�w(o�{K����1n߾-C�6�+O��t;���k�T'��9�X��d�ȁ�6�f��߾}���@~���(���i&����8�?���db�z�[�����e_zh�0^vϸ˛,�:���-���W]R_wο.qU����	��/}�MҪy�MJ��F���0�cx����������-s���!��D2 ���aҘ���m�͎�xQ[���2i�|V��Wi�}[z��13����61:���GsD�؟⽂<�d�"�>�Q(3xٓ��~�#&xIjm&�ǤUCTՌa�MY����o葓X�ȺW��c�puj�\�#�, wA�b�[�4���eO\C(1&2 8�-Ed�h �ױD�o�up�6�3����9[�����j9��:����c?Y��޴h����I���yZ�
ѝĢ9.� �ڑ=���k`V��t5��b"�4�b�2����r���zhYAG�_wdO�� ��j�Qb�i����+�����W!e#�Ha�� ���ۓ;�U�Z��^�(T��/��N�K��B�����4��Zv�pͶĲ�Ȗ_���W�`��y ��������}lLGI4D�Xo������7�r���L�}��_��o�X-^�z��?�D���F*��9��t2��~��ܽ{W�2�J��O��j��[GG
&7����L��#�-8t�VG���=A��Y��W��WT P��j!��L���cFf_ #����e�&G��/N j�&�R�|6�C�#��p��"#��f�8�Q�v|�/�d.i��t���̲�TYI)d��j���J��v�z�z Y�ݤ��-���GR>:g9��xK6��2̤���1���f�`)��DAs�&����(��$C�#���
��p4�Ym�>X��F��W)Oג��JY�˥Y��@��Ю���"��3n]����ո��X�+d��������ɜ��x��f�r�YQ�l8���TA�\�΅�e��]#]�'�z�K!��yJf8�NC����T�R��W�ޔ�y�jV/��X-%+-3�>'��M���9:@$r
$��O��7Y�l���oA�mJ �B'[�- �
������ށ<�q$��&�4~��~��=�쥾ɜ��a[�V���NF�I����s-�qX��Yo���O
�H'
ـ���Y�w�; 2�\s�^Y��u:��)5�J|��0��=F���X�ɤ$x��!�,�@���g�0����}f�
#Hc�>����eg��W����X M6�~�sl�Դ#���i�_:N��\�u�P=�
�,S(M��2�U�6�e����{ߐ�ў\�&���T6j_zݮ�e]9L{�`�<{��M�?��j�α�gh\�>2�Ǿ�` a��J�ز;�`m�$8��F���ϳ��<�8�3��ť,�|@� �u�>�؎�sy'O޳����0x�6Yö<2^[��v�7rf��b�H�C���-��U��>��!^e��_Ә�L������ə��׿�G�?��������WP8�	�J�OT�#
l��6���I��+��4�ʄ6������|�}�stK����w=;s���~���������~:f�e�Q�>f؛*��k	��PGS�J���h�Ղ|�n.lAᗁ����2�ݐl�d| ��G�m�.TP�k���/��%��k�k�^w���]�� $�M�1�Y�KpJ��"w�UV_N�;�����Jr�;tܗbu�d����s�V��g�RI�0���Xl�C����+(1�Õ�G��=(@�%�,����d*�Ę������f�F����y��۽���4s�X�gL�,��Ps¾(�ZsN2nLF���q�=3�0cu�ct,(T��i���#m�����[&%�ʻ:oɲ�2��;ߒ���O?`v���Y�7o�!��?,��z�v)�P�H�M�RV�F��,��Cs�%����m@=�F�	[�a���Z=�ݥU�f��yE�G�s��aܩd��2� �k�\Z^.G�Y���^�ly iu�2><��o���vGz�=�*l%`�ġ�&}�Ytxi���0*�!��3����m�ٮ�Xj� �I���%�LB� �(��HڷZru�at�奔�z�H��L��R��I�D���\:�{�WX/V����K�O?�[~J9��9��g���L�NO����!���@�����G��&i3��j��޽�,uN;�)���^�G?˂��-�!�po$g����]�VX��^	n�@y�{�r߫}��j}4��ř�xo+�"�pu��(��kɋ����+h�M<Y�R�JD�a%�q�zV0/�(kG)-z� ���42Ϻ^� �u��y/)��HП�E/'s�m� y"��IA�6k��o�j�Z2�\���m���^G:U"�������u~��@E��.'�Nw��ǲy��RR�R�V�	�2oj���s���R\���
�	�Bfv)rQ�ft��Qp��R��t��,��;C�%��-%��2P������r��9wID��\H�t.r�Kge�zI1ujv�6�1�-�]x����,�B�p����u,��+�A5#��B�y�bl�~]�g��f�dO�싲Ĵ�[S��e���0����G���}��{?kzgK'RhhZꖳ,��-��9���&�D� ����u���g�~;��g���gK`<sY�\`~��,�r�W[�#�$�s@b(��W�$Q�n��W���I>8��Ψ��N#m�����%�Q������V!�e;�pgւ���>cԲ�g#��u1�����XB�	�g�i�)����>NL���WгS�p-�~_�~~�T��'�`w�V��=����C�c�\�T��2�j�z�0H[�0�-n�(eeGb}���d�`- ��W�W^��u���^wٱl5l�z���˙\̦2�s2H�Rm�ڑ��Ap[�����w2�\ӧu�$��SXx5����rƃ���[쉭�ot`YYR�Ȕ�Abf菉�yl�v�+�([E\�~��-1������|��'��(���[ߔ7n�ak"}��(/�)�1D`#e  S����`��{V����aR�V�fR��~��O��7ޒ����������u���S��d8��^��C��L��Gx���1��`O_u��,�/w������{�$��H�?�7~����,��V��W����/*��j��-���7?���u�z@�:]���ؔ ����͌���h�6�9vRL�*f�J?�V8�*3Z�Z�k���w��c�]t���0�^V�qP�B�yIR�ҁ+���ߴ�����x�E�o��K�d�QwG�-���y�g��߃沶Zq6c'V>#�.##�oRſ�&X��k6�������F����L`i�ڵ׋dU�d_9ϸ����#��{R�7�����W|�@��>����),{uv)��\�{��ޝ7��3 ;+�_6�r�Z���`�\AW���%�����-�ܵ���^[V8
����ZAL<�_�d?Q�� ��դ�yuOA�@࣬/���N;�D�k�ġ?%7p�!�	��;T�sѮ�#�����Ql1���|m�xuJ���qd�8��u�a�Lg��svk:�u����ac����KX|}�=mL����}�g�"cy�`�{�}��_��_\^���y�G�2��|i�:W�WWV�{�y��`8�1�ȭ�[��V�"���wd���!l阾��z`ύ�1���\�~������+����C�o�[ے}��B��\z� `nј�C�{���_Ӑ��ћc *�W�{�(�.d���I��a,S��xIJ�M���Ȭ�b��
��N_n��,��*�3Sն�5�7t<�QngNdE��N�#��F�E����J�C�hՋD�������kh�X��WǾT���%�_P�׷��\92��#z�#}�Ś̂}�4��T���L�#
ռ�MV���R�5����E�V�����ggl%�Ezx��*�R��#�=��*0&D�H�f&7���u䪞ˢڀ�E:�toW}�MY*� (NMTD�A�ԫ��X��R$U������e��
��x����7��\�̕�E�
�;K�%:H�P���4��vL� ����������q��-��kſ����x�;Ϙ��[5%d� R�-��0S3�[�{��pf;	l?Z/�A'�B�_y3��� �K�֢��ׁ��P��ܹ�9+xN�fШm(���*��{��?ˇ�����Y��%�	Y���@�k3a��⭴cm$��52`���r��YeL�=`A�m`��_���.�EF2R&��eb?W��RV(uL���ʃ���h~.3fБV�$g+ؘ\������<�_��?�oI��X�*P鰍٣�	Y��חR�aશ{��=Cί.���J&��� b�v�6A����a����o P���^�������F}�j����<.bpU9��R
���q>#x��,e�J�k_�^�A.���c>Vb;����D�c�|�܄�8l+��
UP+�'��/�����֝{
���D&�M�(0��(����%����Ay1��	�J�B����Rύ��[K��S{�,	M�L|��FC����k�`��=����7���ш�%�Me�cee�C�v�U�f�<�=nn���c��1�Ѽ5`B��e���^�(bMx��>ź�����A�?��8�٦�-��:���n2[��x���l/����(j���^Zm��b�
k29V�q�!"+ؘh�b�w���rG�V��p�P���g�$�e�-��͝1ނ��s�8�'�\�bYZa �����if���Q-���	��z[��4c��$�@��0�i��V�n�=�.����`e���u��!��a�\b�:֓�4  NP�yn��铃7+��]���:�g���QS�J�j��V�gF} )���H�<T�r8K�ʈM 4)���a�)	�߸u[޹���K����H�8o(j�u<�b�H���ʘ!4s4�c=AsL����X�v>�.Ƣ�#=`Hc���Lr0�����p�3�ͫX��� %i��<z(��0�j��=5`}�-�2{�L��߮�4�T�v R�M97�$4%��:�c��A�x�&�B�����B!���v�u�	��^�l�ɥ����\������o�qG拕�t_�sy����������Մb���>���bA`{��Fy���'?��Y�|j%�:?0�0��G�)C��H'�P��%ݓg�����g�#��(�L�_R �5����3'�`��Q��U�)σ3�r���"�h9�z 8`��y�\A�{f �@��K��M&�\��K�7��	K���:�Ⱦ։U>�ܻ��ﮮ��|�^�D�ZcY�X�޽}�F{r��{�;�eur�NMGA(t�@����̲
g�+�H���B���}��ݗ��k�'%�y;�.��'ruy%i��@ȃ`�l&�J��\G\�d�o�@�lW}�l��
]��WGAfa�5_��cq$�����L򋹄e!ݬM,��\?g�{/+�=��<ݨ]�P��	���N���d&ݵir�u���d���G$�A�2D�Kp)�t�f`�X*���� 2xx6�C���7Evq�3�P�,/�/;��;���=eb�j�	�qm ��ݪc�Q'c�`�R�\���7���H;m���9�ͣ6�g��>��CP� ���71�7�N�$c�����l%�L��3��ؖ���Ƴ�;1��P2����o߸�j����E���J]@�Y�������_K�Y�=����/#i����
7�!��ݟ�óA�ҁ���C���|}�
�CX��7�g��j�ژW���mD���D��}tb뼾A���J�{U�ӱ�?�Z�Hd$~�����Vm���6�L�X_mP��|˘Ƒ�C���+=/�����L^��(QŚ��@����U�o!Pl}�(�O&̤�6KA��*���g�s�������L@��u0��25���e�E?)ؖ\�mtڙ�!V�625<������Ml�p6�5�=���EY߯�C�3�s>�lB����D�B�-������p����BGK��}m�i�$��v�ʻ_��F[�ޮ��8>��#��z�[ޒ��#f�کIR`,U�T)-|����M����b��8��VՒ+�7Z
��}=��l�N�or>Q�7���ǲP��������?�����Y)��w�vkv�㾨C��q�+X����ٰ�?aɢE�k�K5���t�˻��l%V�_��nvK���ɇSTY�`�p����!1�Pֵg.*�lFx�&�ARR�\���B�N�%y�4ᚬ�qɔ������Nt�zM��^ٽ ��Em��M�;s�͸������?ɣ�g�>ȳřL���H�VIF �����KI��q�#a�Ce���k��k�,�L�c��T���!Y[9x_Q!�8��};����zR�F[���X��u���b!�E#;q������	e��Y�"2$�4ח:K��N#m:6B�Θ�7\S3��. !MaF,V�D}T�V��C����[�B��3�fc8�X�  k�V��j��ŧ�̱C#��1�����O���B٫�5�UE���H�ʙd�9V��J��F���$�ɋ\F�c�.�d�k�k��2���=�ء�RZ�$v�}=�����=�b�7�� ��*�kj;��]��#�Q&����D���0�,`�o�5(�=~�hߏn���ɝ8|�fs9W0��䅂�3ʿ�A��8 ���eooO>��XG� >=�$@�A�X�w6@�	:�c p8}����@���?��w��g�0���(�C��kEM�R �~��2fHo|������N���\f
r���^��d��L_s��!�iڊ�_�:2ف�� ����=���j�bp4��&�Ү� b��m�`ʇ�X�>��؎�F8)md���U��gĭ{�Ş�z��O�eJ��F7
��VN������ Jy�`���|�L�~�Ǯ��>o�|FGp���R���l�P�_�D�L�ӣ�8Q����"�#�+x���ҫQ{�@n!�\-���x� /���d.S��j���w��[p@ �RYek��Ã=��Um��in�=����z�5�L�`	P��H�2��������P���,��t]U����?���0o���F����^*3=�����Z]�Q���&dL� ғ�T�{(�@�A��k�^5%�@���	�����^[$;ځ
_Șl#��sg5�W��>��EC�l7��*H�0�SJ�WG��,!���I7��ݬ���6�J�ٌڈ7`�'�⹕�m$�e��Z9R-�����S-¶���d�]���<\S¦���c`ו�
�e�l<&[@u���2M:��Y[n�U�dT��8y�|�c�l��O$���P0{��=[�߂h�X4̧����|�6g�y��^j�Y�n-*L��@|�5�Oe�c$H�1p���c��;�b=�Mz���g��NS����V)mD�ON:3��E�s���e6)�Gy>9�׳��A�IM1a{��Y�3(�������N�X�,e&�!$A�R�Ǚ�`8��dC��ũ��?|s[�^�'���Փ�AU�E�D6�2{wr}�����Q)��*�_E��	����e=��C�29��їx��1������9޿��4`�ںVB�n� �F�Tx�X0rI&�J�1锺!�C+�;�#{z���KjWڽ��+�9�;�����������ȣ��ut�gc��J���=�a���a� ��e=߬�BO����p�]^��hOn�FdqCI�Θ��n�k��B��aO�XE�6����h��x?]\X"�~��o�[ͭΠ��5����p
��v� �����2�HDFS�렸$}+c;������pn���0}�?1�(D�Q/�:w}ı���;l�_�Qz>��Cx"W�B�aM"4ޖ��[ �,k��J���Qo���H�L��E�<Wq�a��́[�I4:7I^�/U���D�/"k�;3))�Sg�1lc9d/�_o<?���D�O}qqΰ�4����$��L]��2��1��=տ���k�w:{N���g&#�ז���6�i�h`qF��}|!i�˟�x.����7�ޠ$��F&a!u�������[o�3�������	��F2P�9�\����M9{��� Kу%�����7�U`��\ @���[�yӵ��wޖ��B�q�.I+�s��vG�AaMj�cϥG�j���D�M+lA%z5�<���@������ S��cm�=z��b�}��l�ܔj8<4"#@��	�0cת��SC}��/U��S��=z򔽢Goܕ���M�Lg,;���ӱ���)�h3��JNp>;}!���� ��6��C�a��J�l�M* 8y�B�߸#�^WΧ��?�_��9�\�+y����-P�|"�;{��e��4O���4��7[��-֩R7T�V�LF�[��9`4����0��C٤�|עR`�ֵx��Dz�F�]#xF�`U�Շ��8��U��.��{
t`c! ��1����Å���t��`��{��^*�[��>�lņ�;��ޑu5��幎��^S��A�s���b<�1��g�e�gv8S�`my>��l)�"g��0�f!01P����b��虌�nm��RJ�,6��h,��X�s�Rl�y�g�֐���J����ҁ(�������UJG2Bf���Zf��l���/(�be� t`ӞgJb��S�!���U	U�c��D�n��� !�<K�xw�5J!t��m�q��	�c����u�i�l1Ы���v��D�3q-Zf�+��,��r@!Ry�6�]'R���������<ք���I\׮�j��lO���ׁ���~~z�G|V�i�HC��t�*��P��|��������ˠ��;�uh\�?����{n~�ݱ��H��U�쒕�Ie��B�n��� }$'I,X��]����W}l3I�\yv���V��T"��9%�����-�^�Z1镁�RxUG���EM�#X��O���6#���"�QO����\1�jTࢭ �a�V�~>Q;ו���w��e?�ZϞ�~r�B>���+7�a1B S$[J�$��������_PY�Z�c��_�[�~l�~�NMC/5nH�����*1�e��j
���� Z��LF�Gz����ShE�� �A|�~w,Gǲ7:�$���Y�㚓X�j�x�:��g�}ܻ�2�h�P���r��o��2q&�8�Z���W�o�����-�~�;���?��?�o��I9&�d~Q鲛!���3�ɪ܄�ŬF��ə<���ζ�y|�/Á.��	[#s��G�FK�U��E@��m�ѧ��,���'�BO�B��J˘�B�����01��Db�,��u ������L�j� w=_�c����k�stz3k�i�U*/7�5i������m�OM =8\S�z��}����驼X^ɬZ�)� 2ԙE�`����V�9���M�����A�n�+��lGݳm>��o��L��;����Cm~e{1bP��������;����-0����g�����v� ��o�Ѧ�_j��<��o���ȟ�����Y�B��{%=#�P��j�,���+��_ځ�U�
��e�o"J.��(�����S�W�upK��_8>멃ݖ=p?y�r��'���w
��d�P9�z}uz�m�G�F/�%V
�����2NP���8]���c��Aϻ����^�*FUjY˕:�����*��^̖g<��y�>����zY��ZT���X8(aH�5��m�hd-�=3ism�R�}���E���n�z��}���/#�@4̊<��V ����ԃ#���˫)�XB=WGk���\A�u��yu��)�1{:v��L>��o��GHв�@Q Mhuu�Áq}��K5֧�ۏ~/���o�tvEM�0��& �AN��}0����9]�UL
�d��`�0���|�6���a�(.'��lx��	:׭ʘB�e����mܕǛ+� 8uj�i��K7�A	ю+��AG�[}Y��v-G�����,c�,�Gr��7�i�D�-=�×�`4�Ξ���-�����J��D)�I��=��3�e��158W풙c�-�����R�M�u�6�˃q���D�dxw$�Q[ρ��gsҨo�@YM0�����J?�߾�s[uI��98[]�[�)ヌ:�53�[�
�m#�v;R)�?�u�u=�&m�K� �k2�fj�%%Ef/���2I��{�������"Y�:XZv���qA)����%%�EiFM��pC��6��Ih��V˪ X
-��up�k��#���X)[�O?�B�����m�!d&���e�2�g����!uArw�ͬ%�;���%��R��73n,��-Y{@�O��J�@�"����J�Y��,gd�L�ر��Iў��=���ucI*_t�����<�ZK���o=k�n�v$�a��.�i��o#PJ�+,`�	C�&i��C��{�/!�uj�����]wR[������v�����/�Y>�:�������7�h����8B�k�$FV�G�}��1�e�
�d����\�`!-��$�J�.@+	*0t�]��Ї^A�V��Pm��y�ԲP��g�Ajd�zM9���t�Z��s�v�H��F���*�$Jm�o� (x��\��ea5���g9t��/8P���K���}y�������,��'d���������2���ւ�Z) <Up6���Jh-C^ko86�1���J�&���s|Tu�ǿ�b�R+!���~_�fO.W9�Az�&����X������L�߂URw޺%�a��e}�1CxM�З�KF�tSgI��+��e��\�ɴ��2nz���:BT�/���D"(��n.�M8M��E,�I�⁄��ܿ6,-����_�鱡T�Q��1=�m����^[ߙ/A:��/;h�YkK��'E�+Fh!Z�@J eH���o2�Y�j�Y�R�$�Y�.<d	�5Us{���9�3y��<���� �?Dn�6ʦW[(/�Q��R=ך�q�$�l�YW�`;�F���e�TB�cH%4��E�f K�F�Íq,/�4 ~��Ƣ�����,\Q&����T�գ�8r[e��mϣ��m�X����![z�*��7���<���\��bd=eF������E`��k�(�}[��8���.'ώ�1�5a%�(y@=�@�� ��X�I|@�_L�"��	��˩T����*`�멣��L>�HpxoA�n9��.@L�>}N'5yd(��kAWQ����|֯�:GT�V�v5���C��1���l5���D�˘X˘��!����;J�<�#c�����7;Y�2��mo�k�6F�$�Xi^�y�l6/��	.�o4�۞_#
B�A�2x��@��V��Õ��Θɷ�S�g'�%��>9?�G/N�r>U@�f#�O4�C�V��w�y[�,�@Y9��Y���`{��8��J.�`_Φ2[/�����_?w�Fx8�T��<���p(�ސ� �$�z����0���`��N�5�n��V9��t��g�+e�ӥ,�f�(���e�
�!�{��D�꡴I�C)R�j��9)m?�DUǲ��o� /�l鞿=`�~3�{	�v����U�ex4���H��=\�ɤkH��\��S{�	G"QзI
�l���<
���&
7�R&`Ãf����w�A��+F��q��}�`��ft/���aKz����pA�/Łܱr�I����H׶ֳ6��J��:s �An	-̈́���! �`p��6� ���x��bd	��ekEa/F[Ċ�ȡR�/`�!-�.tn�7��EԞ=3��dȼ�ݳ'X ��=��%JY�5��D�=8�=���7���>��H�q��N5s�4���
2{FP����p,�k���'d�E�#��i^��Ot�:z8�q4�Ab��/yw
i�[3D�C�@v��ٰl�M��,	V�a׸��ݬ����Z'��S�����WD|݅�p&x���I��9�_]���)ɩ�Y��dM�ӌ�'lϖ��������^�	d�*o֡�����yf@j�g���@��{�Z����lӳ��`����]�R���Xʓ�3��K��z�m�s4<K{�o�rq�0����N�q��������M��7VT���ـRV��4B�:����h�K�d`�Q�ʺ��,�	�&waA������v+�v�k$��/A��W牱�o*�o�[��NO��dP(3-��eܮ����n&o �Fk<I<sWʳg��/�[}�������F��)P2�9Q�w��~ϵW���^1��3�%�b����:><�n02��eAP��k��B�{`5_�Gt���PΞ���Օ���Q���B	���/B�8���������4�����<]O��(2zqBM��\z6���}%ͩ�HxmG	��6�DQf�:X��~U^6f6Tc�r{)ā�p�,��b(��pj��� �VW=ү1P���J�
�J�<�6X���<���$^�K�ˍ.Ev��&Fx��ÈOp�����B�&'Rgm���^��/��E柛ĨH\W�"&u��Tb}m���Q�/�ay@�o�� k�px2��Hc��G	 �<�����E�m���mz�#!u���3��zDӃ�nޫH������� ��{�S�j.`�<����4߼V�mư�Em��Eiö�$�1�T �3�b ��ÑzT����T�(�V������7�k��}�e\XgХ��`�KJÊ�TuO��0�,i��:z�}3rKg�m �S� d2`C��@�]��J����O�f��Ǹ�E�{ÒR�ݳr���P�Z�A�Rw �9��5�S$� �ph^�V��k6����Y��0ʿg"q-�!�T��3#�,=�8Q#���mm�\��](�������E��5����3-6�[�D�iSRێ�(9�sPJlN('��-��N�	��?uo�lWz\����Ϲ󽘁��XU,I�H�RK�%Ybt�ю��S�a�o8�7�ڎh��Ў���v8�[jIm�%J$�,�5�@( ���<�ke~�������Sq��g���˕�r��{Nʧ��C(j�='Sf,�{�c�Ո��ϥ��@�dkMA��Q�m�i-�&jg@�A�{`]P�ѣ(�ː�>Ӄ����j�n�;���]����c'���t%a]bU$�D1X�:2԰P�9��!*1��5i�ِ��X���yҦ�)z	�ǺƧp~թɖ��Q�	ƅJ�5�V�T,2FMh[6!�[k����@\��F�w!���J�e�M����9h��S�����IQ�<p# ����OA��ꖣ��s�O��%�������teoA�Z0��:�R���{n�`ʺ��L����ٚ,��u�.��ڳ<R|��3���ױ�[n@+M�u^�����"�A�]?�b�;��M���hRw�ٚ�����#��2�j/E>TɃ3���qN,�).�UĠ Y�'b弱?#�"bD����L�z���sa ���iXb�h���'�IMi�d)a>+�7ߧ���(�Y�H;S���}����r`4��nl�$���1�!!�������B�(yB��<��^3}�l(����ݡE���''���ݮ�S�WNQ~�����r�=�(��+j�'��� ��R0��0K��I-�S��Mo�s=��h��*��[n�#�K��kӺl��^_B_�`f�f�<5�/'�u�3���
��{���$/��;��NU\����Ӱ��۸�DB�����FKAX[�߿/#�m��"�}�d�?���|L��tN�.��#>���!k�ufA������r�m��4IH���x�عs²̕:_h�e<C0ZϽݝm�k�v�$kѴ<�n�^__��:������ӗ˲$�N�ʩИ<*���{
.G]Ԡ㠿��/7GGz0-4s9�/ޛn�g��4V(���^��
��k�(���~2���/~f���`���Պ��S�2�+G��L� ��Ʀ�2��u\ �Ξoj�ǅ�+,u�ӹ6����"mD��I����[CO�ف�l\��VDt%��e�Nɢs��T�x{������`�%g��*93,�g0혱�F���RΈ�� 錙�K�0/L�(��`Ʀn�O�:^itRD(�hh���{�3r�] �����JQ�_��)�t:2���* ĺ��8�� o�`�{�a.�̈́s��[h뿡��u8S���wz��D�ƄN�0��\��
w4�9h��WV��i�i� 8��!4�:7�xA~6�z�A���C��8Mt�b\ٛ��$`�" k1�����x�*��x�=$�E-;�v���s*��Q�NkV ^o�eq��p<!em1Y2�DQ��2̅G績 @��q�,*k��m<+XT���w3+���@�E�j������K}�3I�o��%�6î>�Q�L��
-�2���x�'гgϳ�`ⵜ�����{�8��	 
��,��P�d%=��>D��*A�\"���>�?n<��(�� ��"!���
�Eўdc�m@V�-ìn
�hQ!8����?`�0�� ����f8�j���f �0$��4;�d�$��J��9���Y��s9��0ۄ�1�0d5IZhY����:
Z�zе� v��0��[O[��5'�=�
�i;���)�oktPK@�EH�cC�\����|堸��g���'DZ�2�-���
FJ��U�����uu)+W0J'���<���żԜ�[�����#h����A�����l��'3�8�(ҕ1�pfG-f���t�ֆ�׏g�8B���fb��Za�x��&�F��%�AJ=��E����� �k��B( �U������Q<�\�)�

�n5��]ֲ��6�$��Ҏx�&��y0���̛֗4�Ă`8K�ia��0$�|q
�=��������^L��z��@XZ�8�5��35�����S`��:�Zf��`L8݃�bl�� &� /ی$�~��Zl� 8$��2��� ��|���-�3�C5��q������F�6P��?� >��L0��A��E<�]��lcPK�tYnd���t����<@ݪA��.��u�o�f�e�5#��ǄV�^��چl)�@=����%��
(���_Lg�R ����9l�y����I��I*~����qg� T����`��h�5_�-�PL�Ɲ[��<Mʠs���(�������yv��?��67��@
�+�>O�+s��*ډ`yY���Sn�>���N��o�u��oJ\��>I����(\�r��E�v��;�p0�V�� y����҃�~�wo|L�P������3 .�ij�����H#pb����1貪%dt 3D��m�T!�z��H{MŦ�ʙ��_Q��C�/Y��{�ΐ�Z��\Q��Z���º���`F���1F���p6ɤѱ�9{�'�$��!�E�B�N�H��F��I�N�e�8�:�L�7�{�Y{^r-1��%)�b05�[��RO(S�Xw�9����@b�v6�F檡M�Q�$�>��L��]�^�N�����y�Ġ�TA:X�i�0H#�Vx�f47b5�=QU)������w��;��׆s�h=LvKbM7Æ~{m0����{�[�4��NOv�F�d1#>��܀p࡜؅4|0Q$�E���� 
��ʠ@(��GM7=Zl(@<Tc7��5;�S�9l�e����:�Y�0�cid�.�B'��X���[k=H`�3J8�ܐ2��,H�!r&^'� �\�VO#�t���L�����ǲ�_���҆ʡS��ht>PStꀬ ��ϖ�3;�P�Ŧ><bPcf0�Y5��^?R��~b61F�©�]k���Cf�ҳ�I(� �22h� 0��&�nn���R'C
� ��;k���Z�yP!�+E�O�pPE�b-,��sؿ/X���G�"}�	��30�u1A�������ݦtMA��bb�n��f�%���5	� ��H�&����Z��H��lu��~�Y̊A->f�Ps�L 44 V,l����$Y�v���Р��kflr�C�b�9�]�r�z�3d����ն:6&��akk�����Vn��!�`�)h�?��X1����xx�N�ڽ��iq&7��z�P�U����b�:�^Ѧ�݈�L)�85(����)&f�t�s�Aen�Bbࣂ%�f ՜BcQ�W�PD�:G�(�d~�tn�T��T (��x/X�S��de��j����M�����y�%y�ǚp*$`��<������kr���G��!�Ty3�g̢J��h�X���ҕ� @�\��ԙ)��B*�̿��I�k�̆`}���H�O<�KƯ�Z����6f��3UT����3��%?7f��_���[�}	z�S����e�顉��%�ΨW��<Vl$_3~U<��T$C\S+q;R���#�+�F��,��!��l6�/Eq�B<8�OZx]ka��� �N8�4�|�c�	�,��X1�fS���;M-�^wgZ T".�S�={E�� F�b�p{�3�"%����\!{� "�5�SW�N�� QH�}kSe�h0=���f���KԀ&�P���w�ɒ�ga�	���.E��IR�N��|�1�%Q�L���r<�$/}���ɀ��@�ϯ)��FR�fN<E
�������)��rsb�6�F�wj���E�Xp��y���b���S}:���d��@M!��t�ݶ������d��ni� V���q�}o=����I��X��Gc����ZV�dԠ�M�բٌ`/������ЮPgTE��cY�F�)E�uh�9d=Q�z5�k�P:��;Ƒϟ���b#H����@�.F��ꌠ&0�8 ��T��(|5[@z��b`�mE�S�O��Q����tsջ���w�=F����ҍ���s���ɉ��93���v��'a���L(8��O�ά/�'��&"Op���δ7e��Q�`����}R�z=�p���nl�8�l����ǌ#ƭ�n�MPK��Ѐq�������������򥷾)'łc�ٟ��<�qF�AC�MuY�ia�M8O�.�_��f���z-YH�|��"g
>8���v�/oܽ�@������j��0n7��K��3k�r^�}M�Ɓ�Q��T�@5�ʹ���.��0v��@ �����@(�Mǂ|~���O������W�d�N�C
(]�m�у�ޣ5p_.����{��*j	Q�U��O�sMA ~0�dE�q������du�xF�c�S�XF�d���ʸ�7�����h�j8���,�h;+�4�ZQB/�1� M��2����Q�����à�4�*&{k30R],�kq�Px�`�=���~�����*�5�b�Q��QΠ�
<��_���dogW��Ʒ����V��^X�T8�3T������؏*2b�!�-���`����$�j�Db�_�Jy�g����E:%u�������<7�0�Rg݃LG�2����&G�fA*�ad��n���Y���͜k��ݪ��A�ta�H�-1�M������e�ކ�&Z���K�����6jaY<�E/MXiB&	�as:�=����> �c����38� ���z4�������\gކG���o����u�e��r�Zd�!k�>�����=����4�xJt�f�����¨��3<��NP��6�؃��
�h����KX�N=�L�9	�ym�c���X%�N뭆�SՃ�D#C|OZ�NJ f��C?*�h�c��[f�p�O��&v0��!`Hb��(�S~Z��5��@����=spW8�-�,ފ��`N<�,K�]csV�Q4䧁�=V��j�N0��V,렂�g2S͖�U��vI�f�n��G��O㣬��5U�
WY�#�+[�0�XM&�����Y�4�,�
���'�_�>>�*��B��a��5t��ߡo'���VY�*)�u0���(S09}�9=+�)b�n�d3��Sޠ+��:n��(d�k��x*7�ʆ�Oo����̰���'ӱ�q����#�t[���#�z�Eb���P���db%i�х
�����)��[z�����HuE�OdMϦEaڤ��)��$wLd�a�;�n�����`����۬���d �&�E�3!PI�����aU�`�g���J����D��������)m���$�Ml��*@���e�4�IM��as�<")�n<����Xo�P�]����dE��G��)���dj�m�3_�(�YxN5r�<�S�e�s=�� X27��S�"�>c}GBЅY����3u���fݚ�V�� ��&��뿦��\AW�l���E���z�eT�N��f��NJ�a���} i�*�΀�mu�N��k�x�G��)��1C�����T{G���_�s�M9�]�һ����]��-b@*R�s������0]��eO7�"Ӄ1)�|si�:�pN�|����Ͼ�u9Y,)5_�.�n�/��	��g?*�E����!��XX9D. �eʌB�͍z6��h��FØ�Ee�2�S 8�m���κ�����odrf�'�z�#�ꅧ��r,�zJ�킎N!m�jH)GO\f�2҃���)��d>cVp��s�-�{xO�'T/Ek>�U�1;��-����&������޿��m*�w�Ȟ>�cd���Y� � ��~Bf�6��`��5!Btqm[Kon�n*8�ɹ�y�ge����t����[���y�X_����
~k�L��McY�ǼN�W-,�x�̝���*iLR�`:���y�l �E�h�UL(M���uk���
[
���]�D�R�3'sSM,d� �r�!�4:���dYg�4TU`XT)N?
���̊��Ƶl*��=B�d����H�@�c1��d�PJ�������_��\y�I�����rGA��d.3D�$Z�����-F�Ye�bv�i�1�{��3���P,K��V;{E���L�(8X�ömu��@�˩�6�h9�j�Đ5���z�ξ�ij�>Рp�f�6ƞ4q���4�Hũ���k܏sJ�X�/fN�8OK�en�"D�O /���C� �Y�>+2�sP��(�dg�2�L��?d� 8�5�"U�~+������`���!7�]�N��ڻ�� ��?+ה-_��d"����(�\�s��m��fJN9�怲XZ�ݚ�xI8MY�٘�U��Ňj��2鉶� d6$6>V�c�Z��4gR��"H��hpUE�8���o��ڑ*��F+D�Q�Y9:��a�t=q��$M\4f�2�!�U �4uSV͝����s�o �z���g�XƁ�d�b�&��U}���}�D��=ĺ[�a�J���b��a��2�I��q�C�!�U����>q����Ʀa�.��̲�bt;x��dWJ<p�m
�%��y�}���	\��R����[=
���@��D��Dmu`W����(,���Kw�S��_��p:|�V�f ;	��О�T�J��D��io�~��V[nݗ{�Grw�@���l�����dM��
������=9R@�L#5_�=���[��Р�iG��0!L�2�jV�;T�U�vʸ�ݥ����b,�
�_���n���<�y?��� �H	�̼02o�ˣ����UN-�6�>/�2���!P��q�0�K�R,{1;5�����m&X?�����Ij}�=�;�V��|YۊăO+;Q���!@�L��k�JB��T�e"+�0]�g��S@i�JND+3�d'��8�0 T���� T���H�`n<��"/3�{�Ĝӫ��P#r#����c9+Aa�g{9j׿/Rs
�ꅍ�%qJ/��V����X�W<Rh���6�)���+g��2�n��N����$�%�������5ONd1N��/��A����F �(��^$z�h�q���ІTxƞ^wFy��&뉂��m/��rj"��XZiۤ���ں�ٰs���)�������Y��m�A��?���MY��|~�΍�	>G7z5�'#�q����^�3kt�L���x��1�j�r�[�<A����ӱL�a�=:��d��|�!g~�M䝫We7�d/4���h@�T��{ׯɝiF��t[V���5�yE��&��ҩ�M�b����?�`�  ��IDAT��5ϲ�O��|c)�'������|���՗?*�[�6�������]��ݸ}C��	���tE^��<�}Vz:7O]�,�NM�Wߐ�q_�<3j�S�cP3����{�qΒ�<ԒU��#�3��\��v:t�-yؒvKAtBQhF���2�ψ?�����D����*�w��G͊zʨ�i�Ф�y��+]ɽ�`��ֱ���?������9��EQ���a����
��kߕO\���ٟ�ݽ]��_~Y����1P�Z��~bk&9�b2��}Z��j�bS�XD�������iBu��s�0!"����zၚ��6��(2�Ę���'@�&�����F��!��̲���)��j��k[$&�E���"���.�tTpguҴC�y���ˢ(k)�]����A��Q�X�da�^�Yn0O��?qMݞ LYM�		Q�x)Ӆ�K��Z^� � yi��x:=s����B��K%��J$�X=��T�]"�<��c�/�;�(5A��b�H��5����@ca=��l�0��OK�9����}��Iv8�|�3�WK���g3rC0�,STxcY���8J����lt�yYF���O���VY�E��h"�����VN���SQ�H�^rKgv�D�(FݴX�nX'w�7~Ӆ�E�L����z)3s5�Up]e�:��:ψ+�����r�?��p�.���Ѡ��m�f)�"F}�{�>֝ڏC��16��&Q�����|U揾j��|��<�)V�.!��*�[
��Z}�p���&��3�Ye��`-($x��pz�~�+�%��w�q �j���x"�=>�J3�[F-�Ɗ�P\�i��=֛i)�C��׫�=ֳc��ꌮí��(����N�Ⱦ���N���0��Y��Y^3M�i�ud
h�џ^]s^�J�JY�mS��`�J�M�HX�ٔu�O�٬T;�4�������
�%�-]3��̱��Zi��t�4��4���M�n�꩹ԡI�Z) ��-�/Zz��mV��#��y9��]����Aqˀ}�n�e8y�~�P�� �!��I���4Sʳ=�TA�X;
F@q�fFU��"х4�];�$l�nj�3=B�|7��l{�£��4z���ri�l�GC
^9ˮ�Y��lgjc3�i�X,rs����]h!��G�,�K���}��Z�0��x���w�7ޖ�˱+"�!;0����K��X
. z�Wkʊ@s�3��uY*�0E?�n�k���u��	z�i��A�t\"(�ߺ��\}�m�3��&������@�D�+6�9&�4����j$ ��5[<XR�NK�Z]�7
u���_d;�&i�-C��hӹ{�������rT�Y�g���,��TY���,��y�TL���[���(�^����C��Wlb�~[Pe�C�]^woܒ=����
8���t�n�s ��
��ةs���c$%�"�0�(| �*�^�k��N�o�W��OK��&�j4r<��Ϳ&����s�w�l�u�u��V÷��#��xW�uvS���ʓ/� u�&��l�?#������{8/�F�� Ka�1�<�}E4(ftĩa�����\��>D��{k<>'�1?c9��TLYK�}\У�*�ԏ��O�@uWѢj_aY7�bZC9#n�H�c�U!�h�@���k`0~��?F��=��Tŧ�R��`��3H-fp�A�G�ө������y�/���/��?�*#�P2{�ۯ����e��	�4�D���'ls/(JL��"@D5�"/�&w*+���9��rSI�c�~�Q�}0��?��mؕ��Nڲ�Y��TLP3A����8xM�
N�:�C����k���:��z�����!�b]�������C�����ӧAeO��s�Emau��Z,�NcF���ڬ�)��h:#�Q��[
'�Ϲ�>
ۦ�q��~ʭG����6���v_��v6"o���褪��e56uf�Sn<Y�i���Ώ�� ����0lOA�� E:'�E�����T��]�����P�Ґ� �ஞ�F#��@3�^7�,dvzՂ���+P �u�Fu]mcE�gQf�j�:o����L�z jE��YX39qo��v�������Ͽ���4h�yQ��� O�lfV~O��6�Sx$�2 �R�V@pe�,h�n�к'��ţ�W�I��Rh��fs�'w�����K��+L@��S�>�<��g�?��������q*��:}�ŕ絛����a��p���m�ͨ�����g�~�G����xm]Y�XFU+SP���0��?����+��
W�/�DR��?(����¹P?��휕�;�Sq~��~u:� !�}i�h����C*��e;���%52��l���;�@��
n9Ct|���*�Ҫ�֒��Mi��o�It�¿��+\���&~�����1W��
Ř��y+��>���1�|Eꨞa�ɜ�_��q1��Ys��������]p&8�4~g�t�-�h%�����E�TI�b)�Ϲӗ�D� ����u��c�&�a�7�ǇALB-�k��Ͻ*W6vIE�y�����;��o�{Kޟt�el}��%�\�(�|�y6v(���{���4s�y��t#8B�����#`��oQ>F
sk�{���/���V���ZYS���-%����e��w�C�uܺwG�ݿ-G�BN�������k���ӹ�驽� -uǡ�hXsb���
(&Pt(B������2�E��$�3�{�#�I��L�������K�h֪�HǼ��k�59����FeR˩
�ŗY��K&�&ramKz�B.�=��S�,d� �'�/;3���]=I���0 a����Ԩi���5���'jiƾe��,�VG����5�]�g�bb�]DM<��N[4��@X�2���'�՟��ϟgv����%�ln���b(��ܜ�iұ���L��k&��=C�@�R��\<�Vr�@�X�7iG_��V�9ȗ���ݿ^�ӆEϺb3+��~���V'k��b�����$�9���r��L��tH��j
�3���+���f$z�,�P���K�u�l���}Md6�����	1��I��"+��J�EN�B��7��o�����%��V4�ɪ���<sC�l�"3�Պ�/�H-sh����֜����z�Za=���
�܋h�{2��h6�����~��rW���۷��?�i����䥏�(��"�|�;<���]���q	2����Ei�j
�LE9�a]���+��^��2`����p��&��;�������Hg]����A ���'�!�,#ĉ��\+��c�������uO�@L�� J���~B�a�%R��ЌyW�5:���R����}l9=K8���H�M��jf4W�p�+�_���T�bQHTӘLF�b�w��m'�'1Jpⴛ�-(L������vEOLK)t�~gf5��P�ƫQ��k�QFI�,�gJ��޶t���V��d)��e&ét�P�'��A��%AFH�yF�j;�C�}M�����T��j(�ީ�t�/��i�d�h�uoG��ލ&�bR��ĵl�p���an��Qy)��G��u��lg�r�����՝Y ��?Me5�M��y
16�x2�!�R"��CG�v�}��H��X0���c$�	��^�p{�"���%����Q�x��-��E+0�|��:��p?OL�=q�&oV{D�\�C�=��Ȇ���%��h]�<Ø�ϫ���qz�аx���?�1�����	�r�O��������׌�OC�A�	�w���!��C-�[�Wˬ;�8��\Y�0���j�Xx���ET���՟#5>֋�����'O����"���g�*>l`?��K����;�&�g���.բ|�8�u4e~6���H�0Y3���a�n(5��@����+���ᾝͅ8�glQQ��=��?�V�j�N�!�-�����\6� .�ZI�rm ��:Wo�G�/����Q��6����]uf�}u��}C0~YC>���'>";�6���M�W=�qkW��g�~8��?���hw[�mXVC����"6 �G)��+;VL��=$�>oE�\�d�,��]x��I1gt���)���
Tf
Z����-/\|� Y.�d�� f�y| �����T�C�}�ŗd�ͬ�l����{Ro�"�C�40u$�ui!�5��TASG�T�AǺŶk-��Մm
2
��j*��S0o����� T��^�eR�-Z҆#!��)=���]+H[�wecc�^�,?�D-r��V��qE}��N��l(!6�� ��Yp/�l���ϞM4d pz=�����4ʮ:�7�zW�:��w���T
��xf}O��r�׷T#8ʦ\WA6j�%�������:�v`���Z^,F2�{l��}��H��y����1�2��@�d�(�����]�����"	p9����ۆ��}����Bl9Q��r-�N��Uˌ������3d8z��,uL'C�zb���ˢ}Lb�R+���-��fA��tCPVSEÐZ�Jl�E[P�1Z�>]1��L��Oi!+c]F��X�Q�ĭ )0qo��)Jy�ި>/��l�v�4Z�ҲK)���h$Ǻ&�sp�����P3�-��[��Ȼ7�����g�-l����_c���ZG�rnB3���n��ZǷ�k{���dp,���Da��:�uu��u��g�LI��G�	�g��@[�=��\!��-�2%��n�%a�6��@�yC�=�+Y��`V� ���{���l��<0��a-�9��������z�Հy��V��N0~0D6��HM� ���=Q&;�}�9� eI��Jp�r���@aȂ�����ex��\VQ�U��e�;�
�j_b�8�����cĻ�"��o�ǳv���e�Ј1g잙Q�/������Zka�l�8�eǙڋm��։�oKs�p���pF
�Ϻ�6�=W7&��,�p'� R��Ⱦdp�������{2��OY�G{~U,?�G��i
̕(�#�|�w��i�x��g�|_I�{�[���:���<D|�_^��V��◔����Nߏ5m��*��~i�E�TY��v�������3,F� hu.ڣ0悗٦�2�ă2����d��$+tu��{X�S�K5Xyx��S��<}X�0��`��Z�HY����Dd��/-�o\̌a��1��fORW7Q��LK�8)
��eK��=��x[fs`�j�Q�S��M��1�%&llQ�n���Qa̢��c�뇊j_}����5���e���Z_!��}�i5���=�RB��gGA�GiUa�U��/�V
1����gLI�tJ�ښS���)�>��^����j$�`|���: ��Hu�j�fk�X	�k� ��^/��jiNIi�U��4 �y-�m��۵Z��ŹLb$��)����FW6�m�{�|�ݷd������碏����/����o~��/<���;/w߿+7߿��S�(ouz�̕'$}��T��yG��T����.��L��|���P�J]-r��@9�/�6_uQc���A��ߚ����ᔇ0�lW�wd;( B]Z�'���(��?�"J;�L����n��ڒ'6Έ(�+h~Jz�P��l*�]��˝�.~����M���6(��:����ve{cS��R����Y}ju1td�*ȹ>8�����P3CĽ�`��6�$,n�,�(A  �>���R�t����-�ĥ'�|Җ�Q_�fM�=qYƋ�|���}��K��l��΍7���ߕ#�N��cst��]�[6�xp]��_`,��7�����[�n�!�թY����wK�wW�h��{aO�Μ�����~|W�8�-w�Ck"KI`�J8���6Nmn���-�r��q�@A�dqͺ�-dH�P�T�����2��)
CJj0#8"C�/���♀�g�I�+
fS���s��A�����Z�������pEX�������{w��k��ྥ��h�d�a�N �I�)F��Q>c�^KaA]q�I�������PF�D���Kbgs��30�0G<��	O3�4P�5˶}g���(Q]0�+M��`�A��%�G(�Z��aa�Rܗ�~"{2�Ψ.*�P݃�P��jx�zr8�ڣ����_�۷��?��ߑ������o��4���w��֕3�/X���9<<q��x 3z�zK�?�<�����ѡ\{�#���Hs�G�d��e'��h��3��L��3ę�7dng��3�#7R��^�}��t�`��h{}i0��fVc!^�\��-FPG ��;w0Ȟ�>���B���6��tv�/� BYDtꖹG����K��F�+�(7�0+�ܫ�����+�X�X[��=?c�!������WY=:��{���3i�$�:3u�}�S��-3�Ń7�0���h�\3�W@�G=`��,���nH�?���#9��/�#Yo�Sy:�1*s�[��a���Q碑H��!�	��(�� a�鶭G�~NhE��l�:ԝ3�k����������|UK��R�?�y'!�5�R����JB�Q��"�TC�������k��z����UE� �='q�3��+� �lftdc ��C"h�ߜZM4i�e�*�x �In�b�D��U�E+�Yݙ��\�y(\�Yx��F\Ɜ�l�$�; 	�ȫf��B#�X7X��2T��9�־��?O�(c�ȕ�9��7r��o�f+g��}Q���%<8X�g`�Li6����WlI�'!��B�+���g:[b-�2Sf��-qoHY.�����=c�^����.(�Z�ܐ�f�j�Q:���Ȋ�S����2��k��Uπ�
��Z�[.��ɠ~�%��������:|V����3���M�c�)�9�V�7d�������X�2n��Z�a>�32]Xv���"�� %���
؅�`Y��#I��~�����(,R=V�l
W �uM��RRt�
 .+��M�C�=�#q�m�PQ/����L~�����+�ݢ!kIS�tV����w������Ob=t��m�S���ƶ\�;'�����[�*���s��j��s�+!�"��4T3��es����V9��[['V�{ʡ��F�=�椊&���9yb}W�m�@Fl���H�X����ra�=8����/�wߑ�:�
�(񻽵%��H���f��L"�.�7�d��_�������&v�dm��4���ܒ�مl�oJ��)�FO�5�)8�q;V N�p2f���A&F�)[`>���&�ai�/	�
3����d�?����\V��lkCv���=s^�g���k�]��c�h�tk[&�p�ς�{�t;]9҅ˏE��ᐍ>)�:-�y"��	��IȦ�	���eS熎E#���zG�N����+�ɥ'�������o�u��^s�d�� �Α�h=R�>�4�M�hJf����e�j�Z
�]�B�,�>�q�N�I��S1���k��"R�_��Tf@�|ގ�@P�}摱z�e�.ƌX�`R�^�Ϗ���Sn����F*Tb=)pQp:�����K��f j��Ⱥ�&� �� 5i0H���u0̍���T�zf�L�Z}nX�t�0���EۣP�5Pg��M�r�݁F?.҂hY�=�̈�	J�Z�S����%���E�I��H*�0
��4��?�&�8O�ZDǥ��B�e:˷n\������W�|^���>/_�տ/��1��[w^#M����W�f�w�{N���{���E��_�����?�����yݛ�����]�@�s
u���q���:^�u���G:��z} &{�-����Ԇ������G���E-������pF&���~�I̼E��(��h���{�=ƙ)$~O^R|ʺ�/2*�0�����	w���e��#���ȚR�:̋]��{,"ݱq {mv�K��#|�xZ�@��Ml��47�v�N^�A�K6M�X۹9_Nl^ja}9չm-���t?�r�;�IrOρںl�5d6�3��?Ɛ��b4KD��W�(�Vwk�z:t�7���G'���'d�����2�+0|*��czx{嘹hϣ���"3��$��pj�}�r���(7Pf��l)��U��������+��)�4��-XH�
�B\���C�%�2Ķ��dqJh�?�8���I�1��sfI�X�	#���CSa�c��	�tC
�z�sI.��<�Q��7�=��iZ��ǿ�����P/�����2uԇۭu��L��гS���9�߹-O4��,d��&E��%�P骡J&�&�O�d���Ƕ���G5�)d�,���@f
�A�=�ɀ��<}}�Fޅ����6
�Ӻ����v5�p��c2����)Z�RS?�68�/��S`0��'�&�cY����dR�ն��N����[BH&�^��S�-/L�z K�=�)�`0e�P#E�g�SDa�#X��,�W�]ό�UX�d\�h<����L&2P?g}}� `������q
f!�=X*�_F8,ݞ�6-�D_���Բ�
��3�Cg�PZo~�kȰ��>��vg���O�*��Z���A��K����̼Q��wK�fg����i45k�7�L*�4f5l�x�+G��QB��fS��@�47�Vц$���م�����Gj�@��g7��:�$蓵�����7d��=fZzq]D�u��K]���p6"E������oʆ��a_���>i~��In�XT=u*mp�<��/��zO��������}C>��_�.��۷��z�'Á �Ъ뵪��#Z\Ο<��i�2�������󑣯�\�.�5urh���F ��Q���q�Y��y�h��������}�^H󚬫���qy��%���ɚG84�Z����6we��͈�ă����%��LG�4�����8Q`s��Yi���6���CԵ��z��&�wTE���u�:���0c��&�hF�W�ӛ�-	. �����W�g&:E�"mEQ���f���e,4�hpxo⵫s3�K��^����u3�d��I�uw���r�G��aϢ����tN��o�m�`B�+�b�і��wdǠD��?a�u\p9���t�%G'��2�{a�w�R�u�:^w�?�AVm'jU�C�n-��!��7�a5�5��Ǉ��h|H��P�̠a/��"�vj�Z3[�c�	Ś�t��a�ϖA��ߑ�����{ ��wW.����3����d�p6�;����y��E�r�"�$=��/�ߗ��yK���_�s�[��lu��.�v�{> ˽���@�Fd�Z��6M��B�M/���7�ɽ7o���Y����D�EX2`U��Vts�r[�|�陙��EbNZ�k�M�p�� Uߧ�;YZ&���m��vX��5��(����70X/	�hr_�G��C�Z�՗���\E�� 0�VW�g�� �kd%�[Q��� ��F!���6X�jpIp����H�XK"���B�w�HC�����#ِ63ܠ���j[O�c]ߵf�l%�SLlksC�������5j�~8���"/����F��Y��h�B�B����$����9��o�Q?������2 ����k���3Qz_۹S����*�xIe{見��?�*?�@>D{-3�\3��� T*�]dE=����u-?��j�!�xx^��3p�f�2�6>�I�WS%�f�z��%����N�{�:��Ƒ�ѩ�M`5�>�A�,Vؚ ������;�S���j-��9���X��j�I�L��p����{�������3R�9��%��^��A-=�6�?k����>�go����-�Sᜂ2�ƂX]��2�d�~,���C����#�he�Š<�5�^����c}���Kꃢ?�`
�5jd�P����R� �{�ևLuQي���z]�f^.���t���b�Ȳ��m6�כA�
��E����cH�l6Pf_�e���+�+��e6[X�G�9�3���p"�єl.��[[[� �F��b>���RF;�N^fy(�	mCĢ_��4�5�M��P�� �5[�yK�YJ	����sQ(Bm�4x}��
O!e;i���5u�ҙ��"cDau1n�riϗr��-?��+r��y�����]�Lf�:�E�QF;�;Ɲ��Ո'ރ�f�4'�^_���%�ׂx�*q�42��G@!E��58zQgvwe�ّ|01��)���!2<���t��~�h<�t3��N0гg��MY* Bz�����%:�~�ꤞ��8g��t��F�� }�,��I���'
B��K�B�E�XP,
��(Ԁ���Q�aВ�������uQ�����s�ۓ;�rak��?h2��R�40�eM�9o�tLYSL�A�e�CF�:�:�0��$�{S���/�(�e8}q<��g���x�IP�x�K���+�N�ƪ1O�=��S��,Ys���&� �	�����'E�"��hj"��̾�A��~���6^Kh��6oT��Mֵ�  ���j�����5���AP	e����f8G��pG�&�M9�C�9��ei��l@oKǪ�Ɗ�u^�kJ�*
S6���΀E�� 	R�2sh̡C?.��fe[���W�E��F�G�}�ŋe6_�;<���ޖ�wn���G.�����1iԩ�>(���Aa��ٰ~r�ߓy�v����_�+����?����O�S��?�#y����˞���#��Ay�_��5ewc]���s���������C�<W��ˤ��@�L���]O	�" 6�`�
2;����I�5E�U�] ����\�.)�L�X����s��F�8���،1���d��uL�	��Cs����~h��I<��zf'�:JL�����{[���c�v��*J�A���b�9�,]y�j\7G�3��/���_K< -`���+��H<-y�N^kTs�f�������8���HG��t���T���sS�?����#?����z�P;���;::�k7ޓ�~�5��$�[��no��O<#�/]�7�}S޹��Sa�=K�̀��d��xR>���t�t���Z����Ld=="@��
�xD�-�r�~��
��� _��4O=���acR��JE�]�Z�T��Z������h/1>\R�Db�ٮÂ(Ie��i�r(�T*o�vl���u��\^�$�}��.*d�k�kX*��C�{O?"���|ĠUi�b���i^
V��<��~ȼ�pᇥ�Gn��^+���\��N|*ry$��,d��_{ЋY���D
��W`����T��r����uq^�m��x�������^�Ю��%�eu��6�R��X_�#	Y?�t&F+O��P�:��g��L�]�[����9d�����
����L~Z�<d�#�u��=���
M�.C#� g`����I�© �G�/�Ye�V�i�����}}}M�'#f� �1���7�`U�ɍ����l��R�b�T�3�:�� P����3� ��o���`<R����O?%�n�l [4��.�<Ny�z��|U)�YNЩI==Ó��H�>k��Q[��[@i�i����d��"��'FzТw�8�1���"hA�R���+��/=����ޑ{�Ⱦz�-���>���j�h���WVtP��PO�Z���$+*l�
��v�5��S8go,��B�@�+O��]���u��b����á"���`$�����
�Z�ꞽpYƳ��߻'k��\z�<������3�!�[��x4�CuxQ/���i�:�R!���=�v��Z�;��u�7��/���d>a���D_�~2p>u)J`<t݌�N��9S@�K���������O��3g	0'2U���PP�jrY���@�R/���ڶ�vG��/��|�7�=W�~���gr��Y�x�7�o�!����OԱ����ߖ�|��K_�8��c�Od�g�w|��O>�!�C.�;''���`uYw�~�(6�#��2ؤh9�d�����#q��[56�>���E^����g�1��� D�t� (�Jd�f����oj:��F��0S������_�r&,��>3p^]t�B�55_�l�/�	�F˭gd��ZX�iL�O�WC�*nn a�x�%1*jF;��A,X�}e4^F���H��Y� �Vz1u]�ku�={V��z�����c���ލ���ߒ�ߔ�tP,g��F�X��]i�!3�����c?�t8���6�?ؿ'wo�/�v����k��/���x�=��ϣu���#�}���ULa��:��>��|���?��?�Ṧ��D�dQ�Fʃ��	 ��=%�.�v.uj���0b�[Mt>\���P�L����P�۪S���Kέ�+#�_� �1����":6���R�1[��M<��<�8'�Df HQ f�� ,X�I�[��oQR�	�ZS�lp���� �B�	��Q�F��?��J?��\�Z=ʬ�g!�س���i���pɎY��U�Yw�(� 0뮎K��ֳA�i���%9ɤ9M��?�yf��ܗ3���u�I�����#_��7�����Ψ�}���҅s�����M�6���q�״�ly�#/��/�,ϩM�� R�����E��ԁ�:$����T1.����UC��=?�>�qf�s��qQk	����y��F"�X	֪� ���������R�/�,%(dμXQä&ų{I�<!ø�:#6R��_:�7�N��e���W��zD��.:�E�F���`��G�w�J~b񠵅�\a�:�_,��eVK�y���f�-8��$y9���ҙx3s���r3�-'!�W�������@��Ē_$��HO������ݕi{.�������{�x2R��C5f(�cuGS=[�2=�>������5����8V�j�,����J�=g��� 2x������4�5Z��E���E��O� |֊��m��M������ڛm�M��s�s_� �ITY��2x~��__�� �tm��+Es6����-�C�x�T>W;2��\p���k�j��[����s�NF���{]#!��e�Q�� ��W�d<f������G�J�+�g��2�b�)2�V���[�$����bk���:Rj<ǋ�lw���O�0X��z+��FG�ڻ�������L�T)8���R��u�ęK�g_��g�ɍ���~�����͔/z:-*Q��Ę��Dܡ�8��[uE���"d`$�J,�w��<���y-�A6j�*��'�'}��^�"g���@r���_������ڔ� ȾN"�x���_ʝ{w���*��;�C��/���#��?�������z���Oј�u!�/���D���ё�u˞ \#3(&�K~�^��چ�=�w�P_^ے}uZ�cuJ��a�7t#��>����s�)�!� D��d�Ӊ�3:ѐ�����x�kY�	���a�f�9��D�j(� bШ1K����X�����\�ՏR�]��~E~�?��"����Kt�A�HG�n�uD��3m ��͇#i���#rgs[�fJ�9�hjb��8U;��גF���a8U�݆SوR5+��}�����c����"�3Ŋ����������hi���AX������n�>H���L�3s��s�u��ņ�xx%r�J+tA���έ�
k�)�M��wn�&�Y�`�L�M<�O�<:B��w&��T�w�X7V��Ϊ���N~tM��րK�ņ���c�����Ν� ?��OR���~(���r����(P�{[��)����YrpǶ{��+�+/�ݺuK�*�|���ʕ+�Ky��3ԃ����]fh�z`�t-u����O��g�F���o��\�Xfٓ�����.3zPd-����_}AM���ѽ���FC�f���m�E�d>�0�ReA��`�5��Z$So��]1w���QA�H��|m0S�,\��.Hdk!xMOa<��Jk�)����Lm4~b({t⇑k��L�L���`��3.���Lb��J ��k��?xv�@��z֛�M�$�՝c������p`�^1����ڥ���z?�k_��|���ɯ�֯���@����C�{{_n߼%�{g���K���O��d�L���۲�6�ez�, ���,~�!�ti� ����m��g?+;[��o}[nݸ#�:\�|�g^�gί3��N���ҳc6��U�V�Td��х;u;���ão1����W����v���U�'R���D=�d$c���:��SW������;�N�%񌤿����7�����ޱ�{�*�?���_Va�ex(�� .�y����*�C �!Y���tEs2���Ls��aF-�EBr{+��������7|�g�?�Z�E���n����P}��<�e=m���7��T��M���p��4�"��e���y�hmѯ`6+_���Hn���x:�1D�8;vY۷ȼg�e(H��1K�E����5���G�m��,Yz0�8�?8���/�s���4����X)���6�

�}�>v�㟹��A�I$aP�28�^s]����P^��-��;��d��a���.�
K%U����G��Թ�:Z�П1;F��b�3k9t������W�&)u�
�!�
����>\9?�9�Ԉ8G>�V�g�ZW���CA�'�w��?��v[T����)�o߾.�߾���i3�ٙ)XP ���y��+��'������;ߖ/���<@�v�}��FYx?B�YvQ�J>r)�[F\��z~9$0��]�͐���j���92"��4��o4f�ڶn�MudO#9֍XW���^[��m���)��!A
��K(D�䯿�U��W�J>��K�ۖ������d:��������fK����B��N�Ҩ�p�J!���h3(����nC�p<�U�9��z�ug�
:89�E������Tk���|n)��!���slҍ��l�Ƹ_���>�t(���=�V�?k�eck���Ȣ�����~���:�[�\����D�g��y.���4^��_��N%T�,�u̖;�9l�C���Ҟ�{/�d�2��+tѰy�<�{ڙk+yԎD_�aZDt)�,=�"�Z����S�����)�����~��h�37��!�=�1�{�z��u,3R:�>eYK����P����ҹ����Y{�{�����E�~;j�Y� Ln���O�Xtz����q�+ ��"xDؾ���2tU��P��������H_�䧞yF>��O��˗y��[;|� ��3�;p���|��Wس����~�����c�}8$��5]��U�yppȠ���n�ޓ���ɳ�=�57U���X��7vt�����뒶�rG�ø�?����)�⠀`���A��9}�٨�Z��ܫ@���P�!�X��H+���]ܑV'���/��Nu�D��|��.m���NP�ϛ���S�F9oX�h��W3f�D�)h%^�b�U^f�c�=�|��j5{Q��`?�y0�Q����Uju0*]Q��X��A0�o����rxma���^{��Ϫ4�H鮆���&|�q:���߻�(.!s3ұ@i
���-٨�e�ߗ;�ݗ�c�|�'����o޼%W�^e�c��.���.(�s-��Θ-�&���2X�׶Ҥ������W��:���wd����)�u�R9����5r�F|<\aWĖ�3�&�"���s>����YKV?�s nת��VQA[N=)�e���f�p(e_D\��;'���~͕�KuB(�k6w�%������=����?�I�C�����Պ%�q�K��&ȹ�JY)�\"�!�Q05���e�Ѭ�E0��E��~0�9�g|����G�B�`=��rfd��u��Ѩ�~�Aux�]�\���ѢMԉ�[5󑗦":ɗ�}���b�%���ߚ�%��T��pN�C�������ʽ����Z��6'�mB�'f 3S	o�.Ե����2)H��V�0�����Ţ:<�쩋���m��;+׏��}�)ͤ�����ku��,@PVA�<�����O�zE���]�kj<�� �1ӌ�6�,|�`�q���|*}���/G�+�N��W~�IER��2�~�F8���˦b����P�ϞF��4��答Ŝ��k�`>Y���s�>�������W���w}9N3Y�Eut��zv���G>&Μ�����_�oݿ)���3��f��s�D��Ԋ���t��;��!�����XQE�Z#��4~���R�� 	�&�b�,7Pt��͖�������Ȧ�d�J�8��y���ڭ��F�&0�Ql�^��ݗ��u:��fMnݼI �	t5Oe��#L=�H>MIS��킑邒������Ϭ�
��n���Ȩ!{��>�%�,Y�@E/���L�0�Z8$&ڒH�aR� �pJ0��}����V#��wސW?�	����,����k�ʗ�B^x�%A,�v������n)P^s�DbQx�#�%AV���1�-A�A�q��`�����naQ���z�=�U�Y�p��'t}�	H\�*�c9�<�g���2�)전=�j���r�Ӑ�5Z�]�3��{��@��ڲ������[�,x?�:]ȥN�`�����u�P@���@�9�5��Tb��Y?44%�4u���3�n�q�xSUd4���|V�f���DR��
�eUmp�ǃ�|���T*�롁���?�F�6����ŋ\/����>m���Rz�6��֦��p^���^��^��ᱼ�W#�ޡ|���dwgWu�� ��y_N�G���-�.\`����.��K����' �v�=�y�6�ŭ;�l�!�uQ��ۃ#9M��b2V_�q@���NМ-)� �c���|;�%M����:۾T�Q&������f��#9��l����2���',3���XZ��d�*����F��(�B�^�M-���x�ܺ�lK��f��<�>������G��r�`OC]6��.XP!��1��Y�G^���I�����1y�M-*{��r�7KI-��yBa�|�ߡs�չiM�*�'����Pֲ�l�z�-PN�ZfU�� 秮cP���������G�s4�o�)�x.����T���Fŵ��u���y��`�l2�(��^���9��ޱ8���t�����Z�e��{ԐR�2f��:�P��)_�?�t���m�]��=��p�@�J|�@X��?��8�w�0�,M|C �&�j���H�O�e��<��f��4����AŠ�7�� F��8��@�9q���!�r��q|zͯ�>����A�Ïx���<�U������{<,2��Q]��Vb~<n��<�gRG���P�@�Z��!���r�Ӆ�1�P�o�ų�i��c�f��`tg^Km�2�1�
�|�K��A�pz��`�jwQ��:�Ş��4[Mi##����RSSFh��~_�g�PA���J+��!s����IO��wwGn~��<88�nc]6׶d��S�S�z?�uG ��[/i��x�+o�	d	-�+�O�q��	�L�4q�d"l��:9�˽{w�9����|�rmC�lF��d��a=q=)�v�@��ݩ��
=f�͊3^(;�����`��S�/�2�E9�7՟A>�[�9Hl���i�3�Xߔ�<�����sr��7o�.߸��&F4A�D��*�hʞ���we�2�:�� ��JX]Y7(�5�L��#�b:mQO��I ����drt"M��688҉��f�V��pW�Vo��^7�#�AA}�z���&A_�����r]���r.�^�6�X���PǇ6(ʭ+�C#LD�p�k����F�������Ԙ����+���rߜ��Hd��CF/Jb�v�����X���H�sa��Y���N�H6���<-���Q�����K.O]�"'(�u���]��יn����:[-u�ăh	�L�D����aY��N#���X��l�`6�H�A2�ײET@�M�E�!�ݵ��1$\f"�5�Ra<x H>�H[N���ilѸ�����Q8���@���Y��$��5�\�c�T�c��/����ka�'�� ��A���T���� KHgܝd ~d�p��F��b����@�:y�k����IxhL��9P�c�¼(�a��""`�gqR�	���4φ�hR7P�luT�pB:�Z�ɉܟ������j7.�*кq|_���WՖ�e��m��ޞ<����dGA\�Ӗm]W�.]d��j_���a�:]C-5�]�i�r���'�Cvnuc�И�mn����eM�D�t-|�ŗ���K���8��e�t]OP[��S��_��ǕX�%��Z{_�t�� ��@ܷ�H�H��֌�s|����+�O>3��,Q�NP$ � @�]�]{V���qo|�ˬ�H��!�R�U�/�����Fܸ�V���W�C�{��vJ����"�9��$��"���hC����Td��l��fr�cY�}���kH{�9�Jv*"�G�"�4Al���QkG��5�z����M6�/y*h��(���$�E ������u�~+r�P&kl���X��_#r��|����b��Ҏ{&B�F(�5ޱLc���M��d�;f�"R�7��-~�������N��F���Fr���?b��,���IBw��l̇j,��6�ލ�Ri7	꠴���+G�V���`�ψ2M-ë�g͋�k�j��@w��ģ��G�}����������zy �w�x�_K��|��yJ�,�E*fp�,�R0G�ڙ�2.�^�v�Ӝ����?�}�}ɰ���A��Tpd!�����>����p�~�7��G����K�����{ i%P�K
���ƅ:�5x��E�Vj;g�XJ�L�4�5��	�	�岨R����+���A����3�q�ڊ�Z`K)��zp�"�/*��PU_�f���^>&;�hE�x��"vٵao��l���+#�����~��"������!�S��a0��/��VPOF`��*�Z��Am���Y|�X-.�H�(1}
��|�gT0��D�^���ȳ��Օ��C�8yZ���-{�7es�)�AK:�K�T���=�A��!L�v~���Kl�0և�g�d3;KVզ�Xc\f3�'%��n�e�>�n���w�m���ek�|�_R��$|^�� 	@ES �%�m���_�Q���<V;/P�za1/Lp�S�5uRp��>ʵ3��k��d#K�Md���hX>ұ��B��6��|kM>�������2�=�[�]����R��YFC�M6��-&��ɞ��Ή�N��e [�{feܡe*�@��  ����OI�@t���5=�v�5��qL��i=�rk����de�("��:3��  �ٝ�J8����e���#�7��?����� uC�xs&�@9ޝ�m��̼@Ru-�^l�}�?E��hL�MVW �ICA$}O�� {YTA�T`�M�)3�(t#��8����ޗ���:��$P�EުԬ�Df�O�vw�����+��*[[[t�i���6W������	�X$��v
�z
�+����x.8QpΓzU^z�U9z��4��dW��5d8yØ��]kz` �	6)���d��pŘ�P� 3����T,��\_>Y:�b�������|�;ߕ�_��6���:O��k`4���7�TQ�N��ʭ����h�b�Rn�a��_�;7�3�ר4����O>^�(^Z�LA5�; ��O+��"�UH*^������O �	�)C}+���lJ�.ڇ@e�h����� ���V�9��aЎH���|A���(M1���܌�V�D� \S�Ӯq������Uuܚ �gO(��:����My{����̜����_�Ϟ�����\?*�uY�e���vw������Msfq��&n@�������7Yv��)�m�wm�S�|Hvnݒ]��Z��Ҍl�X$�P��F����Y�#���b��rS�H��\��b���yӔ{�M�W�_��59��"=�HO�$��0E����lr�Y�u�BL�y��Yapm^kzj�q��̯+�ýLij{
)3w�}��r�z�!��L�ջ�A�!g5�7�� �FY��h���8�@�AvX����_��Ï�nYz���p��+����f!�SO��V�tT3���ݮLo��LAz��P�22J=� 5\u|��:�~o2`vxy}�����50�R8C�F�4R<mk���
�GZ�e�R=�GyT>���I:ݑ.j��t���=�iQ��w��c���͝ws��j1���A�4	�N�v�����CA�?.��y=m����u�=��A[F��V��C�~��	Zrab %�<�����Zf
N$Z�L�YP/��Ew�/��v�C��%a�0����v²�R� ~a�ʝ;O#��T�����{*�F��������y�Lq8�5��g�C�4Cfd!��g�=�A�!:�9k���ۺ�� L���7ʁ��ju&���eg����A��]��<�Qo�f��A*�v�4pS�,�M���NP>���@���B�E���M�E����v� Dt1�WA���#P����4��.΀x�b�j�^��?
_.0��U� K���TR�'��p��2�(iE�v�#�Ο���m���U�`Kڍ6�������`� �"9���\�aÂ-��R���X��4��S�<:U�E| c��Y���;��֕+��[o_�����}�ߧש�s!.=}ʽrho�[�2}8��K݇~<,铌����_6R 1At3-����W�u�76@k��P��QP����Dڑ�<��|��E��":�g �?rYv�X2�\i/ɫ�ɋ��&jo����>?�!"�:��oDj�[���"K��� EN5��j�_ ;:%x.�F*Kp�A��Pg��'6�l��V0u��t:�rmgK����B���d��H�?���?Ea����a?c����d�1G�ҟ�ٟ�/�$/����"kFanuo�/�s^���� l����;\@k'�J�Q��n�1x�)R��l�P�Wpi�2K��5�M��T!;�r���ߏ�~��M*���>r\��s���weW7J��^Sǲ��=���`ٖ�:��󭭮ɿ����k�_����}��= #�iLH��$w�ԉ�����q�� <#+y��Q�mߩ��ƛ��`csc��"���a�X�T	���Mࡇ�g��.|t��=�;�����p^�"M���͍]���5y�sLN4��v��Cq0����v��ju��jrSA���+/�x[�ҙ����\C���|��e����z4�w�u�YA~ot��� �	�"��@�{Ń\�2Q�V��0�P%E[�#���%�6�%�a��YQ9\�>S8�h����!����@�La�0vȀ����]|��*Ԁ��>�����1��1�	lQ��)�C�ߏ�ʠ'5��j����ڒe�u�4VVd����[7佛7���.�Z��u�驶2˚�ݹӧ��;�ʆc��3�y�@��m�vwv���-�~�\���Q;�qh)�Zk+��5���9��t� x ��MsР��gZ�ĒjR��h�EO����S�ېckGY���^�/���*[�Xﾽ-�>�����U9�r\n�ve�|$�9�Wj�T(̼p��%/P#V΃��ϊ�U[88��r�w֢9�-�\���v���\���������+a����$D�͙s /kM����l`I����E1ROY�B��m���"^3�v0�NȆ��'2�S[���}����zVP�ey��M�=+
�'�8�W����~��S�/Ԝ�gu= �c4�D/<����W8�.<xQ>~�)���ʏ��N����]	�{���_w;�sZ��ʚt������m���n��")�?��Aq2�"��8�b�̡a��w�+.�^�E>P��BJ ��x��ջ�F�͋�{/���
��S���/���Ƌ	�,.iu���K"W\�f�p��I�3�3��,P���"�Z������rf}i��0�����W8�)�LjY}ݿ�9�v���"�j��l���� ��x�8�S��.*۪���8ǡ�۷��βm�5r
��G@�ڕ�za�N�Y����h?R�(W�b���g�xN��;6�0�eI`�X�.���z�J����} 1�[�W�,���=f}+�V��dJ�o̯��$^<Ɨ�^���c��Ӽ�B Bg̒�Z�S�NIw�KqhT�Qj�h�;RO�]�`���?OB����9{DKn��(�2ǂ�3�ǠF�� b�[[���kWe��'�
F��}�Q�	���B�Y� ���5_������f�6;�F}�O]xc$��6b�,
c����^`���]dӁle}ٍ����I�7��E�z�b-l�T�UH���A�T����:2:��W�l��,re{C�޾)
'�#E]����#)��I�GƑ��o�P
�W������
$�Qy^n(����/��-�� }��32�%��@'G)�FV ��O�\�FlJ���Mq(�a�5X��U��K?,_��?���:����'���S
nn�c��W_~�N���d
�H7��A���3l7Zr��Qf��}>E:��Q_�k&�#���f�T�q���,KXo�͇��i��-���՚TNEVb�w �w��\��u9�� ��Ɔ���T�
�ŔR�F�r���R�c������q�A���_c횂���=��ڣ����>#���޺-Nǵ��.�Ӭ�N4�yP��3�)x���7��m�n�d��8���Flf=�";�0���s��@��9��5����`�"��"UFj��`�>��Wޒ?����~㖜;��i\�q9�6byoS��nʮ�]5�=�H�LMf��p]G&�Ӊ}�2�+�����M��o�6i���b��`~XG9�H,jL���s��H&��-��Q5�q�u;�:菈����*�Ǫ��Y��.|=�t_6u��c�TaX��C]�UB��9f�As��	�y�aU>��WtmM��Ԛ�*Ufm�=b�?�B�o�ו�����h 5}{�C�u]벵�+�h&玞�sg�ʥ��}���`������v��3���gA�5������3�z������󠸪��m�	�����_�ħ��C����5��!{���-/���|���� ���L��DΞ8%�|�	�t�A)�
Fƙ�g#y}�=��k����r��󲾺$u8�1����r:a��$�yT���l� ^���u�x��@��0_4D^�/f�ގ[<�"����P�|eq��K�<�YF)}H��_:*��=R�m]x����o��D=��Q5T�԰����]K�;�'��g�������%�M%���R_���ou��ထߪ:k�M9�&�˰o΀y���h��,3�(�Z���eR�����jm��q�x�#��59v�<�����|��I�owh��w��W��G6W��q�M��ؖNp8��	{H�g��yQ�|��������"r��B�+��$U��k���c�&���4��-{�Cp�b ��"��Ԁ>��%%#�t ]ȕ*���~
��$�͡�������F<w��ߍ���k�ߙ�1�)17���c�X��{���g�"�X3[�f��h�v���_�U���>��!�%�����r�W��252�g
��sR���,z>�a~����yl�'���C��F�����i\g�A�;ҥ+55���P��km:�����Ϭ�>X.��,�{�鐵�����Ł� oＧ�	Yw�`�yU�H��΂&3g�	�#<�@mQ0e.f��1�CbQ>���0�u�X������o\��B�7����a3j�'Q�E͂"/�T�h��>�L �v��马!��Š�6�yټ�I0�}���uO6w6��ˏ�G�Ġ�D��m�f&Rd �k/Tw�ǉ��B�����o�`�E��ɾ|��ɠߓm7ѳO��؆�&�V���=U�vC��w�yE^���$����rVwg����~��-]5�N3�9�/6In��d�  F��f,�o�)XL���: pi�)~�,�lqg�ws#o�V@}�2]�� ���z� ,��o��N�}rt��\y�]��l
���
�.�b�d���y�D\�G?���Ci5���o~S�x����C��o�Œ�5��@Pfuy���ýb�����2cup*��=���#���$rى�R5���% ��L�N���
k�\V��4'��uQu���+���k�g���˨ח�@���
nf�h�pf�q��v��)����k���/ #f#{��W~��Q��o�3�ە�IA�j�5]����u!���ϗ�V8�ؔǎ�����F���F��$g{����*�����RitщXp�«T��ò��TŴ��9�3Z�Fz��������G�Ͽ�r��)k0:���LDP&�vS�w��zM�ܻ)�%]/t�
��!C�-�lldi�M� �T��r�`A�ڞ��:7	k���H׮�~�5�Lt=`;~����7nPbz���瞞e-M��G��y�Q����hgY�BAH^��a��=3[��X1���g&��*��3��/�n:
C�W�����˩#Ǹ?X��}����?�w�_c��
����=y�#���26~�쳤O�w��W��T
/]�$�׏��ꎘnd�q(̀����>cSݙ������>GP���xb"ChK��Q4��RB�$�"�L8�(����|���<�A��@UU`���G����Oʑ�U���������KO��3��ep0�>�dY�P�і���w���\x􂜼I�i��"6���BHM�k:q�Nm�6�Hh)"R:�:'��:,N��ٹ����ſ/�bG�g��I��Q��LYh�`���({4eT�8�7�/�m�?��F�n�[�?�Qd�Q���R-�����Rgk�'r�?�3�����D��}���
N,"ㅫR\�����r��QL�t��]L
:���b?5*&��t}�z�8�3?z�1���"�O�/�����7��s����m��h�}�=��#�C��f-}���~�Vtl�V#U�d�O��e1k��v:g��a�b��x��ޓ�3����w|�|�ӄY%^+6�P��ҟ@ݴ�U7�����=�%�3�w��~%^<��<���Ĝ�B$����,�h�޹tч����+��F��*7|��s��/Q�} ��=٨<d�"��Y��Tk���$�uF��3^���t.�D�5cO�u��0�w����"
��v�b)֪���cy�Ib�82��6!E�&	��*)�2gjz�.ךL�t�����k��L�����.t'��f����Q6V�M�Dxɹ�c,�9��ݎBP}�%�ע5 ����"���Z�C�rt�������ޟ�{g;�E@h��N���s�n��7����L��}U޿u��9��l�M�^�l-��G��-�Y`
��Z5a>4QPUl�nxJ�B�����!7o�NwWn�g�}���G�����Y�����@Oc�=E�ʠfq��2��9ލ��]Q����c���g�7�D��j#����(Ң ��B�<�Z����j��� S�9Jق���D}���:��t$#��!���H�6EF��/�1xF#c u��V���CŪK�U�g"���)���6�֘��m����KR���m��)��J[�в�|J1a�d�EaR=��8Z�?������ؼ%��T���Og� �،5�.q��߿}劜T�E��?C�`}�M��~� �m5"��?Pg���D_g��b8@�x���Xj��W���b"
BGs���7T@5��q�"�
B:�.:���yKfi�b�>zZ��q�O��B!L�sG:�(�E���Z�T>�[�,bf��$C
�L�ڪr���܆���������g3o��T7gkmU�軧�ne]7H��b[����V�%� ���������Y���B��;K0���Sxd��"��a��8L��4*���V�OD���L����K��/}�s������L���`W~����ҭ���d
�����ʼ�������ùyd��X���T��}]�b"�ݿ��`,�N�"��L.����.=,������7�]^�w��ه���e$��|����M]3c>#�'ӹt>��!�ǅLeP�*���'�F���Z��n��f<$��� �����
�H�~����z'��/�g���~����xH���X�ӷ��]�����d�`�tг��������<x������6Րz}���kP�ksk�j�tO2���caYA���Ȁ�W-���N	�FCƓ!�[aQO���d���ٱ�Kgσ�
���{y���䅟��v"`M�+0}�Oɣ?"_�������*Su�?��O�g>�I��ܖg~�cy��7do�'�G��}.�'���U������Ϳ{V��%9��}�
Ȣ�{B��(�-I�^��:�N%�"_��+��Wp^ߠ8�l1�"F��� Gт?:����`�i�ӑ!��e��`d}8�0�^�#��k�+͉��!\��^j�.3�2g9��B%ݘ�|��Og�q�D��п]��,'M��F_�׺2��3s>c3嘭> ,��L����6�֋.�[���d2�Ku#z�e����O�cr��#���7XË�6*j���dmeY�&=:|2�����ԏ?�|�������������_�������?&<?-�nV%��}��p �O�
l�u�EYp�"��yn�@�́-"�e��̻ۑ���1��\����k��\{�i���.����|���t�y4w'��
W��,�=dk���#O�f���bTH�� � �i�޾ʚ����^��` ܇U�H/�X�Qyv��I�k3}��زsv|[V�׼a^~� ,�a/��!(D�2�e�+���֛�32g�Ƙ�B��r���432 2xˉd�r��qnYD4�v=�P��v#V[Uk��`�^�k�Y�ߐ��-������s+(aH�j�+9��5�����5��E��JRf��������� ��~�z���In��<�R��W�煭2(�5��u_% �Y6�<�k�L��-?r�>ʵ�nȖ���>�~�++�e9u��A�'�
6ҵ��L�%���L�0�;.��Á^s[nm�R|�%�{;���}�qy��Oʱ��^Y4eM�D1Ι,���-E���]�2��T$���u���~�R:Ӊ���h�N��:�\D�j.L'��[Ĉ�����"���G�sD>����ZS&z,�Q=�"��7j��th4q���B k���41�kQ=YD�A���Qk���)ex��M��(iQ����O ��
�p`uC�tv&���)��-�S0���������~>��x�z�-dR*%"C3!p�� 6U6����j�����P�jTo5t��H3�+X��m���/���g���
���9 t�(�3�L%��I�2������\�(:a%��XG`��o_�x��#kr��y5U��G��N�@�!�aMv�!��V�;��!;�ʌ^��~�ʹ#��d��j�������a�զ�G�R�:
���1�|�����d��I9� ����}2��`������j��l%����}�,<;7��#%w��dԧ\)b��Ȃ�2"�

���ȭ�[���#o���|�+_�S��'�Y_���7o_�g�zE~�SFU]�:^hf��U�>2X{}N�҄�$	|u�P#
�g5sr��"�Wp�t��y��E���t�|퉧���Wd��w���QO?~Y:?��.PЍc�!kU�&��Δ͊�����Gmc;������:��!�Sd,��;�}�j�G��\�E�c+ԏ|��ѕ5�~���IwwO��{�,���#���O|�ʿ��/����+���_ʙ�'ICn��H��
��BT��v�@���sr�չ~�ʸy�� XM3T��.&�~��PF�|i�C1��nO���ʵ��Wj
GR,�}p�V����������q��ֻ�#S�O����j��ۈ��s�z�;�o���ɫ/�f}u?f���������.�^�(o?�l\�!�c��N�ܩSҨ������T$E�Ə���'�s���~qF%&��(qA�j�M��V��[��X�#�������6�L=uNJ�L��2&>���9��r��Rg�*���y�)�}�CJ��>� ���|�'��R�w�C�F௮�$�!�:�fT�W����֕�2۟It0��T���ܤ<<1���]; ���momS��҅���F/ZW0��c�S����Ҫ�%M�̹�aA�ae}E�{��]�u1�M�R�g��~D���/�Z{MϠ=�v��sgΨ��Q�h��*��������1��O>wА1,
�\�X�o��i�I�s- B'��_3>,sP�bg��yG^�w�U��(���XCy�F��_k�	�&.��G��{�ogʸ�etl�d����������	Mr= P�����Bpl�y�y���hq���b;k����3+[�8/Z��{��W}�;�"k9�@6��G�����'�d���^!��m�
��Lh� �8��Tϯ�ڰ6ꏇ3��2��f#��Î%9�i3�e	j�c�;��:�JK�;��/�Z}��-o�(��#���`t�V��f�!�\��1~8ϡ{���gcك�%�3?;6?}��a�2�8߇a��͌�5``��`��8Z��YO��u#r�'|�.��6��ZfnJ̃�ήH��y���"=|Q����ާ��p����H�7�[�YT�N0��}�/���w����-7�P�+F���ٸuS���{p ]�vC}�'.L�cd1!er�3�2��3Ai�u������$��KJ��y!>{4c����8L�j�è���]�"kIČ<� dd�i��O���|Z:�z₠ґAY4��?��t�x孈����"�>yhi[p�sckW�ǯReĻ��!��ypl����b��%�J�!�>7����ӯ89��*�F,[є��n�c�^�+�-C7��RE�_~Xj�β6d�����:2��IJee"�j�Ԡ xM�4�G���`k��t9M�ܜ��������]�m�%���Эw�� ��Ev snY���l��
��ī#�GtA�:��D���jj֐�B����|"��]VdUZ��Z��.r�Җ��D�SG5%�/}���
)�r ���P���Nz�E�t3@a��V����Z�#�eI!�s���i/��֟�ސ+�Uki�j�����p*�;2�52fԤ`�9p�I�P�������T�#B�T�Զy�wRE��l�의g#��s?�箾.�s'�̥�������L=x����Q�)�`��u
�6�Fx���_�j���u8�:6�VMR���#��+4v�Skx����d����pz@�>u�|��Srߑ��t�6F[@C؟(#rՔ <f�u��T�¨�(h$���l�TZ�e�,��EM��$gV.�������n`�IJ'(���K������`(�_�V^���l;�(���#��?-�yX�_�f�Ö.�ZK�h��9P� A����ZS�!�w7o��lE�!2sK�K��-̢E�P�	E��Ά&�q�}|����G�=/?�rE�j3G ���%�C��3�n ^� �s�H!��2@��J8 :@)R�o�����/�{7��:!�U��F� ����[��Lzy�'�I�X[N>r���9+��m�G�9>i�ؾEm�@A�RgE�bE���P�f;����q1V���stj�g�}Pn&A���X��u�
gm%�e�ѳ?h�u�$�<���J&��9Q��}i��Ns�̃;�}����Ч�jf'�3�X�Ϊ��:�>���� ������/2D����Yb��(��J�D��� qE~���4�򙧟�/~��<w�E]u�C���o�)���we�����|�s������Xm����`:�����U�@�_���,GV�u�@O��_��ڽ��,'2�{WV2eoR�N���w@p�����B� �k?�-P�J�F�F_�=u�<$�?
M�%8�!�7~ej��:��(���9�M��z���'ƝE���H�BhJP,%6ہ^��+�(��g�un���,bh|`��BM�Wy-��E8
��d����*�<灇��P�����0�ٛ2<�C����|BgU}�*�G�1�0��J��_�A�gZƹ��~
���<�ȡ����?�^ǹ%�O:b�_W�U?S�h���Z�cS�iMϹ�Zκ��LZ��\<q^�?t����I��Ez(� �I�U���r�i�ˁP�8г�zO��w.�q��\�%)��,h�w|`�,�>_Ui�a2s,�{u�9; �HB�O�n� ���R��j�(��v�Y��!p�~dM�ޖtZ��yk[f
��Tj��~�Q�#cGM�PO܌�(`|ԯ�^Bx@�e4K��/ۻ��Gwe��{��	����@���Q�љI�ȘU�kٯ���]��\d	���,ᝀP�\�����#2��A(;dQ{��gC٤��E��5b�b��-f�dPk���I�A�TY��ւ�0��0|���9�t��dD�}ݦ��F�Jf�����ব���N�Lv᝹�=�?-��Hɡ0�>#�� ��No�
�૶�ޣ�x5�Ȓ:�C���(�<��˩3
 �@�ru�Ba�ꬦ3��	��DN-��cWcQ�)yPj�m�ɕ�9.;8�<\߸"?ڼ*=uDk��Q �F����&6*�4�c�Y�ԲY���*�:�ջ�` Խ p���?R8c�s��n�O6ߑ�?�I��=�	-*��Z��Í)����C���:�ӑ:�:.�%T9���<�x,�G���Oun�#u�ri"�?,]��C���R7��
4�D;:�39H,z[���4��3���@���h2�qQY(��l����)R6�/��`@�Ѻ��j�g
Bjp!�nq���@f���� ⿼��t�b��3� �֢M��>ZAH��D��_�L<ƻ*><�,t�*�Sg���r��,����_�w7���Fr��y䁋�*ou��H����+,�Z=a;D/���Q�"�.Q$)6�81��)k���@�8pI������Xh��h��6#P˄(ӛo�B���V�w�]��{[r�?��xDa%8b������G��}��l�AU�����0�^z�5�x>��ÊŌ�P�Q�k(芽�@a x�c�q��������/���6D�y2͌��p��̕�0�'iչ���-|��~FU�`��JgmEv�!3�C1�T`1�5�8+���'���N�偃~�{����9��+���l�ܑ���4Vj�ZJ��ڐ%�;{Ӿ����h��	V�]�b:�η?֭? diע2�n�oؗ��b��}��x����ќ����46�Y�.���kD�}{J{oa#��+1**�X^R�TN�T�f�!�g�o��祤!u4�������2��x[�So�f�P��Ij,����XE) R�.-��}��W���]��$U���;�9��v6��'�>�����2�*ڂT�**8��Tj4�*V���F�I���3F�:-]�����cG�R@�/����)�֯Y��O����`�c4>�X��ev�/2
��μ�J.�E�q�։	��,��lD\*�Ν���N�¯�ʇ?������M��|Z�UaΜ���Lc�!��4|�ܷ9a"m�o�P��r�-�FO|�'.�+RV�2����X;)3E $!�DD6���(��2q%��寻�Gx�^�S�d� ��r|Y��[Mx�7�_��q�x�;�g�fe��wd�t���}q�8�)f�{����7�JO��p6d�d�Ҕ�:|�)�����-UR[O�YJU�M3��X��h��D�	 S�.2����*����L��iOz����	}�CP= �0vQ����2Z&����giǽ�U��C���~�7E����.���|��s� �:d�*���!@W��I�SW��Vzľ�(y����Nɉǘ��e�������:��C�v������
��,)C�����}����߲��O>��\x肬Y��Pd�ZF�[�:T�N���*�!�4ǂH�+C�����r��B7����B	Hu6CQJ����W:oVj�q#](7�C3���42�̤b43�h��,1����r��{gs1A��&U52����T����x����:�*���k��i�r}�=��u4��"��~=�����ߡ�E�U�Z('R���@�?cS���p,)���T���f�~`��L��`D��t��~�u���0"] $�qM��V�W>�IS��;����`�>+mɊ��6�� x��Ⱦ�f�#,������sd#��[s�w�Oh劺)�&q^@S۬;�����#iU(�R��V0e���p�{ǉ&�0`!c�~|653#01cG1��<��&�p��I�N"�*��T���V���+��û��˨��޹W�+d&�hhh���h>�{G�`�FN6z�*ʕi%����E�`�vx��w�˄�J��2���>���?�T<�^sk2�o���K�}��oI��3{��q��#Oȱ�#���_��|M��v�����K�?�u��-٬T	�@�?'l�<=�-�v��\~�v>B婟��-#d�,��i&�u<F���&AA},@O�
�f�S��&*���%�v����i6�ժɛﾣ �"_��?���1� ^<�D�f-M���yS�/���[7(�&�KPF�JA���,�ڢi�K/�(77��:�FMVΞ���z�]ڳh@P���	���,AK�Z�)1h��h������x:aP꺓��E���Z]Z��� ��z�����}Azݞ����g�}��X�7�f�-hG8��v��ԛ9}�|�럔���.�d'�Fv #x����Ku9����w��8˂崈��$��(3G8�U���A�N�?�>˗y�'�u���b��x�t�AƧ"�J�Z�",>�V�,����k�S��������v�e�3����x� �<���2��4���*���nP�uk�Ƞ���l$����ll������h�7olpCavw{W��wߔ~����$U=o'jsw��&o�w�.�kWߓ{���S��s�D�O�&r��җ��_}A:�5���l�Kh^Ξ��^&��_#�+���mB2�<C̠͝��`Dy���Pp΂�>/fP����7��qB �>q�B@$8�~�E���/� �����c^�(����!1��8�k��.bh[�e>3�p\��������S�\�>�����-�o:����n��a���YSH#��@<V�pM��T��V�e��*����z�?����h�gB[�o���o}P!!H1d>[���\��U �bo�B�d��i��l�V�󥡠oMAJ���t���?9����m=뇺�TZj5����d�v,����t܎.��[?{]֎�c�NJ3�ʱ�u�&������5i���Q?5ͤ��@��-��T
�Y��L��r�M/��c�\�Ҝ؊>��,�?�M�*^ u��B���](�94c���}��?|�en4xxxq�
���A�٤D/���-Okđ���������{���w�Baz< ���a�Ȳ�<yR�xAN�>E �d]}	��o�УֳЊ�'�
�{���鴯s�|�Ɂ����( �$ck>:`4����-͚d#J���w,��*<6"����,�f���uX?""��m�!Y�(�O����$ZH���&�"#���
��ˁeD��[��r�ݔ�>KU?�f�GO���Wu��cRa�, ߛ�awU� �(��^�@�TF��~��ϒ�+ B�P��f�� Q92�Z����G�?X;
��L����>�Y�Ҷ�:8h�1Tgj�q!5��8�ɖ�ϧ���7j��m�є"�Qj3�i���W�愍�&���(�z=��-Pƍ��⼧oyyPO�SI�P�x�*P?�a "˗��,����&:`G��ig�3���O���>m"��#��s^���d�����>!d��c�O'��M�vXD�1�p��l�>�1B�<d�:���hz�?�
ߘv!*cW�[�����}����A��E���Tc��h��������������X;��"ooސ��z]�U 5�ç��t_���5�}I���f�)�VR�lΕ��h�@O��kF�⹁7��Y\p��!���˟޹'���_(�.�,K�Sa�L�u���=2�<�n^ѽ5cP���(Sa���@/5Ps�>��ے�;�,�`o����+s^������(����@�v2�8�%-3�'���L�b4��RgIN?!��P�XSN9*=x���e)4�#P�+���ȁ0k͎|�㟖��O����~����?���(pu^�
h�]4q�L6����%�v�����Ϭi=w�lNz�����I�u�l��q�Bf��ĚB#�`,jj��0���\�^��y���39��{�%��lQ�� ���>a}��	��SQÌ�~�f����$և�)x��ڗB�
�N^1�=�����>����(K ��m#Y
1�`�@�������Po=R��~�:���LF�!kG{}���ڊ,�a3�	n�2!��h"�]��Þ~V����Ԑ^W��y�}Ƅ82�=���X�tv�V��xE�Q���U4H̓蓄V����۫p���������Q�M<-L )�2c�Y�ڻ����!'���ǲ��	����ͅ�س����g�1���дݲ�yٻӇg�6�w���c�:	{615X�7�-@�����Yd����^fe
��K��%���?��: EYw_>����ݗ�k]d_C/�6g�9N�����3ʕ��UR�P 
�1���(�#x)&}c��ѽ�V�䚱t
��5�v_i<տ�^���?��S0x�~D6w��Wޒͽ�F �ȑu����s���:��Z̀����$e^�X���|~
����b>؆P��β��3���>A�Y!�]������r�G��_�Yp����ex�O�"	T���I��#�F��)Y)�͂���)d�ɮ�Sc��{���lɭ���b�+���W���
O+D�5�.KL}��"�%�P3�$d�e�}�]D��!@���I%�%��UL��G��/<�ǜ/����(����+�~����ʉ]Ѕ��\p��!���׽~��!���r��4��@�Bρuh��m8%ܸ��G�����pl�Y�5KH��O_'��4z�$�l|l�ٸ�b������{�2���D6R�5�@��\o�F��Q[E`�N���v����S�'�8#gH��&Ł�e�RFZ��!h�B�BͶ����P�k@!i2�������uL�h�av�芔�#$����b�0��G0�Z��Pϭ��uSe��K;����I|�7�G�eg�(6n���V]pFC��r�p� b������hX_뭐�@�^���]mUd05�$(�"�
�X�c�S�x�.��e���

��٪q���7PQ��3HRLd�B`�A-fF)ݼ&�y�Y��cOɩӧe� ���������nU	�%#;Ԩ���� 2�C8��?�s���T��<�VC�B�?
�=fV�Tq]��I8`b	���3E2��wq���֪5�;t�SݣH8Ƕ���"!�ăw��ٴ��D�H,;9���,T,5����S���=\�5`��g#I��"0���:B�@�S/�cY˦^�����zb꺾����G�c��P������s��) h�1���P���[�g���iuڬ����{�k_��|�3_`��_�����3Qy�X �V���6�LUS���`&�8���kҿ�/[{7�}pD�����="�'�� ��~��0J�Y����l�>���� a��b�Xd�O� .�0TƑ`X��7�:<Ԡ@��;���!����� f`2O��5�6Sd��h>��,��,��,�:��Fdju���Ϥ�58��r]k#�++"2���b4�NV��n�ڔ��^�-/������
�A�59a�ń�N�����ݨ7�������DyF�b�	�i� p

�ڞ�o��졞-]:~�;������<����Xp!Ĕ&=��9�g�Pm*��0��aq�R�K� ��T��E	�σ��-�i��I�CU6f?��͝�2o& �{�+�yD�2>��wZ�[B�Z�o|�b@6��,�E<���笔�˼�����}z�6���� �5翄֎�ב�1�\1��(�fL�k�U1�օ$�k����{�u ᱱ��=._�����W�g���S�0��^�ڟ��r�1��R���8�+4_�e78�*&�Fv�t���j�f�jK�gS������-5�Q�c�G��mk��P36���ť6�� ��'{�޷,���ް�v�&�z�����*1�����OLj�ovRρ���D �N¯B�� �b���aTN�*����~l-c������-���߻�J���~~������y��!� d~%�ג��Z�^�w�z�R��E,A8-�dy�)�f�2��{[�PU_�b���� ��̍Y�������ڎ|�ܜ�|��:������7R2�Z��,�;���u��ȕ���9���.�~�h��g?<�s�y��A"4���g��Ȳ!WC��<�x$� u*|�0P�̽���dϖ�_�G}I��"v�>���� Pe��&��+7�;e�Չ�E���rֶ4�!h��D��W���q�W[�g����:�.O)��jY�`#V�.DD�}�-������6�^�F	�:���"-�k����4�
��iaaRDeC�@1�IWR�
_���@#�BP ���#efpBʅ9��!����@瑠P�|#CP�F���VL��_.!��t�g����F�ѝ�Ӕ|�"6a�}P�� ��	��ظ�Jǣ)�|a(`���Y��i��ɶ3(�^���P����>?�}� �!�����{��
�喼y��|�����/��?b���q�=����#ڼ躀>M\a-^�H��h�RoeX
��s�5�������c`���Y �	�ݟ(>@���4��<Z��.$�+�IP��-��K �t-68��u%c����	��Zp����-�Io�k)�#��G�L������`
i=1���)\X�v��Ɍ�3i�B�߽р����7�0 SL횠	#�����N�/[7o��ښ�.-��1$P�r������$�<���U����|��_��ڱ�<�m��|Oj:繂z�'ؿ���O��^��.)�ԭ�Ԯd
"bu :�g���w��?�Sg�ڞ��X�3GV��6V{�>�#�ޘ�99ǡR�Z>�a�fP��^����͉�����餔S�G���W쿋��^c���@�#ʍ��&� ӑ�
Ow�h|r/O��ڿ�,�Z�+r��$�:m]C�fB���z!�K+R���sS�d�"f�I�?�8���7�W7�,
�-���Á����r��M���}�a���(��GF�J��0N�N��k�z��1�Z��$2��ԍ����6�QQg5����AM�x�Z�:Δ�u��deeU���\������ ��w����9�\X�t�����j�+���@�ܙ#�g��E��
R�I����}ڢwtW�:�ǿCd�����w���(D���"����|�;����}Y�2'�Ȑ��������Fhey��!�ȢpI��1�e3/z��>xvz�C���ɣ�����r��'=�#��%,��.�e��Ji��2��^��y�i�K��36��u��4c��AZMx�=Lն�lR:�%����zN�vVd�����lK����)(����!����3[� ���)�{�z�l��9ؠ���`��1�. �؄�8�a}=l<��]-���Q]��� ��/�>��w|���E<'������I���&��b�<�ς�\$�f݂�β�]>T��0{�3�]��P�ry�<ʿ�T\,�b)��~Dw6�ǁeM�H��ްh� \��q��e"W:p��	�ҷL�G��G�B*��@�����P�N�M�TW�.B1�&ޤ%y���-���d�ѐ��z8L(@��j ��h8��:��nH5
:A�����w��#�l��D �;/���2�\���LMh �d��j��
�M����`��v\��ˮ��,��z�C0G�e'm��u[��X���N�!�Pe
�j;���U��jg�im]ȵ��'F�z��%b��٥!A���IGԛS��f�)Ս��"5����"�1���dJu���eÖ>@<s>�2w��44�U��Rv�ұDhޯ+g("�P�Z׻��X� �nY6�ͳ�r8>1�a�/��{�����d��1#JX@�Fp�-�rS�
:�^�P�xZ�?25n#8���5������]|O��f��ur���N�Ȯ��f�@%�dA
��n���'��j��Z� �u�F�Վ`�Y��<���*"�I��ϝٿ����9�/�Y4ҫ���	�5�6�Z�,L�E&t�rd��:������=7��b�vm2d��Xߛx�'��U����5��`9�g]�����ֿu����ViXT?ν��?t#���K�g~ �x�)��g?/+��	��?{�}T|C;�O����.�?���e�ʋ��"��[��D&�`P��x 
yl{bS��d2"@���F,X^��l�@n�u]�'��ڃk�4Ry���������t�h��,B�L�c���A��܀6C���� ʉ��t��^��!jн��{�( ��m���H*�=�CJmt�(!��F�I�Wx��b����|꘵G[�ZVaH��S�Jc�vq{D���J[���4�V�)Q��Z8�zD�/�̅�:O�聘S*NC�=C3z�����ά��Vw_�}��M��H�.�ʹ�X4��D}*�
���A�\CTf���~�^o_�uܧو��wt�M ��Ϛ:~{:5�d]�|(�4y&��#��a/Fed?���!���x-��ُ��z=����$i쉯�Bi����3��u��*��AYt:�t#�Ll���>}���/?|�e��C5w؂�[ ��G �DeCu���W����k�zk��S��K�w�]�P��|V4����0��.��*,��J����V8�'��:����<t�|���{[?�vS}��$'ds��%ПC�@�oETH���L+zZ�3��
�GL$L�j�Q� z!sE?T�	��n>޲���%������e�^�Yo��ik�)�ф�ִj*�jIX2��<���2p7��v`����>;��ė6%F�6�33��q�4&s@��
��{�����/E��:DS��|�(���p ��y���M�D���'�/���D�3��jn~O�oG�7a���l?(O��;E���_+��3�\���g��̘�tG��%_�pq�W"��� Wy�h����-JJ��������{�> ,.:��i�8X^L JHM��/�X$�B���E1c�
`jY���CG#�Թ��t��$�}�I���9�CG�ˌ]����olQ�&T	�1�+�h�:lV_U���Y=�0z�"(Ͻx��9��tiU�/_�Sk�叟��\\?�z����2k��/�G䔎���7��_x'���〿���2F��*0��H:ևF��]i�ӗ�Kz_�؀6Z��>����XG쫆�u���\a��5m����5��C�U�c
��Xcs��q����#��dM-0�B�WD����}�j ���Q����cc���@�� "㈬(�j��&Dg��y-���Bq/d���Z�G+�E𡘙�<�o%�xf�:�?��PVe�7�&�C�z��f�w|�<.�y��,2���=�A�aU���[����	{����Vx�@�$��h�@�6�)�=|�]^>d]� VhB=��������w���u2����rQf=�\!ǵ��]-ta���F���>��GewwG��u��TRC�fI�,�)YZ1?�"K�%c0���x�efm��ze����n���kc�d��e���쁢ԁ�2|>���X��3wxȡ����;ʟ���ɕu���������h�@��c?"���@�����ܾ򾴓�o�H��-V��k͠��Td߫�+'�^N�e�����j�E;�=CH�ґK�.ȉ3ǥ�׺��9q��<x�c�;�ʁڅA>��t���k��:K���E5�6�^����w��Xw�f���t݈���������ԙ�a�����@�&�jF<�+:U>G<��ى��}nEwT��,���Q`���Ӥ�CK4T��׵�}� tG"���Yiv�j$�:Q���{D�,Ԗ�@�Z�a��`Pw@�kG����<�s��˗e}eYVmf�'��Y���w��s/��=x�z�p?e��O�r��s�ՔcgN�Tυ;���!ebihѓ��2Q ?�9ϰw ��f���M=��������McJ8)mJ��Uw���_�B&-�{�`�"2��Y�J�\hPnʔ����y[ˇ��S��Η�7"U�uR�����(AW8��d�w�/��]�^0����"����=,�H��kE����^V3����"^j���/��(|Ð�����|�((��3�7�B�נϟ��9ړGN��_x�|��w�1k�]@����x|4�]*EBoz?�v��4�2�FAvSM�]�%��u�]C��VYb
�FD���.	^��K�#���2�f�ѯYmA�w+D.u��3��b��Ȍ�[�Ͼ��2�d/HT�I`���I�)���,��x!��Xt8C��R*d̔=9�����9 ,}̲߭���[�4ޝ�� wR�E�Ƃ#䟵�Ev/�����X�]c8X�g��"� ��)�>����'�`@ tД�O�$�J$4���ׇ�o���ETF��Y��^o���1C(��@.�]tps~��QDE�W��� X��F�^6Za���<�ڨ�Sp�0��l��V ����lW�Y��$j.�P?rtMA�w1���b�!����D SL,�C�	��	\F�
n��Y�l�o��@�%5�ĺF��X�sg�Ʌ�s�&�+>�&�
��d��h��`8�27w���	�<6�$���
��[5�+MDC�qn���}���yK����z�8_�e�^�A�J� ������Y�)$S��i�(6юB�
��z�-'�V�9х�N.
��UHHe0�]�Dh(�
�,\ �=��r�4z[������U
֚:	��&�l��������/�Y�h�X�ĂN��N�.63��tjR,7(|�ޙ$9O5�2˹UY���s ��w��r\FN�3�J{�8�:.�k6ɱ����eX���L*�bA����L�J�Y��(u@-LP;5#M�QZP4u�`�@�t������d���ā� Ѯ�g@Q󗡩$�
Ƈjľ���DZo�aP��� ږ�O���G��u��C.�W��e����_}Enoܒ7�~�2��"��V _���i03���t��XS�Ds�.��cB�I����)ұ_�iZ%�[h�ux�`�B�{����G�K���, �K�5�+��g(����������K�=��������r����[�������OV.\���#�>)�c���^�?�c�Z�&�dFʍ������\8wN.?��l\}W~��K��'��l�c�T��'_�����Φ��������N]���ޕ[�m�̮�}<�k��������iJڪ˾�@9^_;���7�`͜S��@D�!c�����)Uw��j3:3) =ԑaI]E�,���
�g����g
�F��LF��L�]��A��M�!܃z���AO�vƵa�ω4�w�NA�� ~�s؟`OW��^LA8"�]���|U�ź7f�|��'�ެ��hՍvK�WW�]ױ��C�@m.Φ,5�[m��E*��C�Lǥ��ҽ�22�}|(��%�����v���K���]\�DEw8Qد�՗�� E��"e	���l9 ��'0��-4l�6�^(�t���y��}���2N�ߘ�R���-���	� ˛Z �̐-�w1��O�C���7ċ-D�J�l^-:���8��3��A�� ��O�?�ϕ�����kׁu3����*�;��jS\�@ ����C���/��o�~�>�E�,�֗���1�'�W.�I<���a��9Qյ�^�5�`��FQ�:�.�+2�{u������۹����}���}���~�
���-f�+()pVߌ�\d���7�fɲ���!x=��@�AD|����������%U4�D)��,+���!��f4�ELA	��s�g�=o'~���ŗ"E���`�I({��~�Bx�_)�z�L�,�c��ԯ�HJ0)���}k�ܭ{�ղ-�zT��y�*��F�e�T���G*>Y=֦���v�j<7awDj䰭Yt>y��k�Y�0I�B*4������~g&�f�����0q���W4J
_9����3�����8�=g�U	�|��F�r�)�B��7^��ۮ5��bDb.�e�g�!�ae��2d�Ȳ���<Ud�7Kj��k�g���V�P	5J�{���xY~*oH%Ӄ��`�c�2����2�X�8�M����f����{Rg
}�Y���o��2(G�3S���?'Ǔ�))y�\/!���C<8OL������W8��͈��ˍ3$8�{��/o]��^��DV���/Y=�Wvo��~C����~d:Qs�H$y����H橗�NL��	�=��%�f��:s���'��V
fS/��W@��`9?���=���@���(a!��G�RS��_�?sF�(�����:��7a_����F������ާ�.��M�Ѭ�����@3ϨHةWI'��o��Vd��ګ�ZS�!�fw�w���=��a��umC�^�F,����߇@��D�P{� �|V�@���SH�|����G����sk���>)u��6np|��<��t�o߾-�[�l�����^���ݕ���޴I������kU�������;�B 1"�c2�$3}�'�(�L&i42����1��H�!�;Ѝު����=32������{_DfU7�9 �����ʌx��}����~����IV-�����s*��P#s��۰��z˄�fzlQ�ިb��Ҝ ��cPC����jk�Q[������R:/{]���d_Ӹb}'���7N����\�pY�m֕-.-KjdHP��j4+r��eyF�GܨKW��.�u��/~&�Ɉ5���!T�<���η�%+
H�ױ�ƿ��<}�2��М;��ak�l|������ƁL����Y�[r��9��Is����)�`Y��T�J(;Gtf��@��[�~�K�R�4$�E�`�%:�F�����kԚj�t��z����G��zY�oX���K5�P�h؝�x0V�9e��Dϗ�ϽIU��>�g���`��1+� U��V�!k���R�{=��7�%Y=�B��aG�Gw�S���nJ[f��S�f�;��mV�	��J���[T�E<��>��>�C=w��{���\.�G*�ښ�6����{2Q{V�V�X��)|c^��ĉTO���K�k���Uu_��Α�=b�*zr��MΠ�e�|-N��c���*'�?��#f���o_C�b�����Lb�^�L>V@�q���c�k8��EAɟ����<-5?����A`U��|pc�|��j��`���YF[�h��8�E�lK�)���w�^�,�������Ҡ�$B{eQ��\9wJv�+@0����];���%�ڼþ�LueH؋������Z�.+M�w�@r����[���ڢ�k~��C"��^ѭ�������@D�i��~}iaQ߃>�֯4bf2g
��К)r����	<���M2�� ��P~�M>"m�+#��b�K����7�T�աu������������*����oY'E_�ȃ*7�X�Bx6t!�T� ��|B�NM��;��?�ic_p{|�@[��y�� D �*�-YC��g���73��9��ZQ"�8ю!MV)�>�����3kS�.����[�[�If)� 2g�ߝށ��6�wXΖ����/)�j<~{�(�����������C��.�{��sκ7����]ch����@���LA�)��Ē��~?9'�P�Ԇ:��y�����{�Z7.$1�
'�y����9+�B#��^ߢڐo�	�9�pt�tJ��N�#],x}I�V"-
�"�_���7�5��k�N�<��>�%5 X��2B#P�"C���^9p �3u�'=��S��+��X��U�g��wސfj�h����pxI�ED�Q3����-=��J��.8�Hu��AνR%pٟdG�rg2��'� jP٤{�?���Y�*�pCh�Lb�9 � Ujjt�4���[}1��!�d�<��(��EB|���|n�>nN�V0Gwv+"C-���31mN���YG� �w��������u�˱9���#�g�`��&��i��v���*��J�-�,�X37#+X�Kkg�/�.�u�����̧>%��e���s�e��2�ơ�Qa�PN1��>�I>)�v����5z'��|
:๔X/fQ=�a�2[�I*1�RR ���|W���+_�-��/E�G�w�z����w��=y�g?�{��k_��|��O�^k����$����_�g�@A��d�v��4��M��:�.��,��#�}�HJ4�zj� �z��f�:P��2�N�����_�����/e{WW�n�p�A��{���� ���Kr��R�~��%u}�e��!9^�9>��k(_�U���&���� MHG |i�X���;�gX�_�/��S�e����	t��:�9��r��=iUZr�{2��K����]^��+K�q���ٍ�-���d�h_��X�U}έ��� ��CJt�r.4�:�,��7���Z�=��V\�ʤ^g
�PG\�C�e"�N��~��So(| ���Ȑ�F:��I��b�∈�K.��v�v15(��;ꩍ�O��˲��i���
�P�][��Hߵ����N�@�9%�5j;[��Z
ҏ#
35uB8��l4U3��B��;P۬���� ˋ+:>KRVp��F�A8<�����Q_�6����;B��t�kB��Ri]__�=�c{��|0��/>��Z1��d�C����9����Lĩ�g\�I���-�s�-���9�q�o� ��N�ُ:G�
ylr������G94����7̂Υ+|�@���}?�<K�Nw\x�cߊ�㜀�@�=R�fڗS嚼pnY޻���L��@֏��֚��Qs������]-��r�>P��@�d]��SKkrv���M��tz�K�?$�W ��y��ԩuY<uY���r�������ֶ�ݨ�SV�X�E������î��ao^�����9Y�1�Qu�-�s5�N,��8��H������ˤ��l��g(1��c��E�?�DGg�����G8�A�����eŵ����j}���Vf.04�p˶��3꨸s��f�犻�4������R,��_����f���OOd^�!]�=S��j���F�2-M�� T�n���� e�{8���i�����\�,���˦s���k�n�|�f����(��R*L��y|̑��uAfB�H��7��G@⨵#�wB�&Rɍ�0u1d�52{��F�g��"@e��N2�i�̤��m��N�8� z�0��h�A_8��j���(�I���2�g�ݒj�I �(��
q�afY��Aΐ)e�C�b
mEnlR�LYo@�(��@�I�!kclD��Bk�f�Ѩ�bL���3�XP�̝�0|�t뢃T?h�h���Æ�,�� d�~e�N�P_�пO�#�k���WQp��M���%"!��QQY��g�Rcm���v׻� �R�5>�Af� ��@��P
��b�����A̋�̃B�0彁:�c�'b��4Z0.��6*T�Li�;��מ�����I�:���E���¿>��/� M14j�e�s��h_�xG��H��/��L��'��%jQ{���+0o��dq|ľ��� $���.��a��W3�Z�tq)�o9�2�i�O���B���:�%��N�n��D�K��x5a���r)��Z��r��'��ߔ��-���3��hU7�woސ���G�K�̈� ���v��}Y__gm��ၼ��uٽ�!�N����32;d��b0��9����nsǏ�9�ts���F����f
��)_\hQ5��j)���WMDdxԓ�û<g�Z�Jb��Js�uw�����MIЏHՖ�sggG�},H�wR�7�v	���5 ���<u�2�hv|��D1k��q�ٖp�P���۲Pn��3�Ige9�)����t� ˕�ܿs_~�H>��O��hMf}�n�ȏ������?$����";�u�Ndam�u� *�c�Z]�VV�_|EZ�s�=�?:�:������=����q��������р5��#;���`��Ml�����(�^vu�AdmB ����n#!-��6��dA�Zx@I����V��ܗ�����cuyuI��d��%�������/���e��12�#r}����c^"��=U'���լ���d��/;й�$M��'?%����,7�4��+`B�<��e���[o�-�����"�I*��NW?����9�N�����"#�����cq�tJ��5%����R8m3"/����}w�YjO͏l���d>�?��{6�w��s���=��c�g�-������������S���X �t�
x��{����I���	����_on������I�O��6mB!��Η*���-��	����92�
�d|���"���H�P`y�)GN%��d�[dê�l�E���ڊ���O�ǳh�R��tTa#�`�2�u���ʬHʇ�Ӭ�߅&��Q1C�8r7�}��_"�P@��)���r_������v!戲!$"�_��L13�9q�8�sg� ~p�|Tw� tx��Ӡ�,��Gȕ���4��}w�Y8����@
z+_�r?n"����G����8���U��c�π��`x.jE�A �yA���r�/������'�Q��(�ӿ�:{�2�I��ǩ���|�������?���MT�倃8B.l��( ���Zk
lpF	6b�'�p�Ǌ�dd���M:��� (��Ut��.���"��!3���0�(I�aP~���ݱT��H�c��)8�k�̏�dt��B$�F���N�8�8Yb4q�y���/7�{�X�:��AM�֗�����T�	YVGwA��P�SVU X���"h���Rg|����*�S�=�+B'	��N�ly�R�������=C�~ ��g�N�Dh���?+ʥ������|`A�1�!0�Sf�S���%8|�?��m4�+���M����N�D/��9UoZVL�E�x�_�ssw^����qYK>/w-�E|���' 6��^�H�ѿ���x�'�vd�^���2��=�ȷ�ܿ}GK5f� �E��2�e���3��?�����S�*,� �X4t������F�D����F)�	c^�n�i�lGf��G��P�� 0L����ˑ�����Ky��7�����Շ�h��f�٣;7>�{�=���9��WN�ٵ�r�`�=�.+k4d��(m*?��%°i�"Gqb4����e�"(��@���?��z ��N�������׿!DF#c,�NP`�� ��5WF�S,U��v7
�@,mE5V��Î5�F��f��Vaﺁ�]��w�#?��[l��+/˿��o((\�sCV��"M����mEY��[��YWupp ��k�J���[m�lcRc��!���e��׾AJV���v'�#�a�,��ޑo�[����:��K�����o���ץު+pn��_�`gJh���t�&��Ur��ƶU*������ˍ����R��$�R���y�l"r��15G?��Y���.���˧�z_,wn�Q�@Ze��g.���Un5�#��K
$�G�.	CG�JYG�.��fC���s=4�jD|��L�ɖ����Q��\(�+�^�"*@���=���s@X�"L��M��e�R��6�#V�K��,b�$�s:�+�����=4�96�x����zu���</�oe���g�k-2D�xP1��cx�w���ɻ3���O������D�
'(xd����v�s�A�o���:���D>B���ɜ&ĩ�%�R�X�����2,2%d A�l��#�+tS=��x��췜��6U߂*����o	�%�[��'$K햂��X:�]��/r��)Y^]W�S��*�C�y��I9�����}�7R��gQ��&� �f�1S`��C�y���$��Z�ġ���>{�{0X��r��=��?����-Y�"m�&����ҕ���Z?��.��.g�W5NG�\�����J��ɱ��1p!�ʠL�G�E�"?:0�q���K����"@�1�<_����^��,v���{���oU��Z`�k���9K;��8|e4̜$��5�I��J���6>��@�f�����d�us'��:�!|�(�!��E=!�Gd��a�B6���}v����s�c&b����
�A� [=��9�%�ra�<����B��że����չ:�I�h�.�ބ��k�Ԭ�r�΅��o^S�eҕw:[��L�D!�e>��q�9=��$t�+
E�40�s�f"M ��IdZ����!R��'�z�IN��\iS*�tcE>{骜o,�Q\D�=�{���>�J�$�j3;ӡ:�6D��/��Rg,Kz!Ϝ>'�ZM�ݸ-;��2�XK ��$c�����b��"�[D��l��b�E�Ư�c���y�h��Ũ���tL	)(bʦ�	 ���M�������1�b�����P������z���e4��곺�ߓ�ӑ�U�@�`8�� ��D_�;�C�{c[b�!��c<T�:��~�j���@hc���*����UtY��c]�*�O&̨�oa�W�@�Ѵ�C~Ħ�l!�ڨ�"�l0�_�-���\7=����?���{��DVy<�M(����P��^h��M������/�@�L�Ze6�AT�"9�\���s֮�#�{³ (�܌��u�uVrQG���<"�ݺ!��7�7���rS��k�'5�L�f'B�5|ƺ��a"��uY)�V�����^�@�17qЈ&�I:�:`)D�D�|�=�Veo��S@����Z�sg�)H��ԙ�rڣ1{�B����xAH�ד��e+5̠֕�e��E��%y�r�Tvd�ŝ�}ꎺrkC�N��-��/F:�5f�Q�����z�?�JԔ˭uYC/�|B)td� :��	k����|���ͺlTk���GDl��u����^���c�;��x/2¡Α�>����\S�K�c+�_\B�:T���^:� ld2�Y�D�r���66žQ쪣klo2���q�ؔ�Q׃vCW�=/_��dU���ή�ll�@���Ρ<�L�2����e�aWz��G��P⪮��p
"2(QQ;0��T�(��ʠ�2�T��=:��O=(,��o�8V�7�7�_�⼡=�{r<9�����L&�?���bM��e9�ц@4,	��г�Rq}���$3�� �
��o���
�aԶ7��u���=&��)���_B���掞�.�z[�+R�רa��"�����Z����7,�����!`W�6�c��8^"�98,��(��V���0�}�3&z��T*��[�ta4�NO�#l$گ�臘�M�YZ�@r�>�W,E�9� ���d��ѽC˨�s��F� #�|�0�'�4��(=��gwN�(��;���1;�X��Պ��,L|�ծ�Z��J��\�	��U"��V�O���|���DZs�J%P���~s"C���L}u�������?�A��(����`��I`X�ܹ�'�5�ppO�
@�	
爀�)z��$t���1�$�]K�3����8���l�6'�B�2�<�6�-N��N��!��k��lS�x!]�uH���ڸ#s����&�mu�^=��|�ٗ��uY�7%�B�e�~���~��Ӄ�_S-��0u�i'�������D(|c�SƓC�A�ij4��Q�v��.+����5��X�����8��\ܐ/^�*��.��bѬ��3 ������;�ߖ�QW�C �d`��FV�K�e�����3/�"C5N��@�;�e���'��rF�^�O\�;=E�2�>�Cy`����rB:�w�>�f6>e�y �_�Ut�����c���j%
Kd���'.
��i1��Q�?Z�Ͽ^�3v������HA�p��b���e�9�4��U[l��
�ͣ��RWl����OBf�%�Z���|(�B����Uٹ�� �NpIL��Zo5b�v ��D��B�Жu�z�!��9֑�_bY�k5�zPg��5��Ŷ��َ�UI�H� /ҩ�r��Ԥ����R[hX�Z-�Fd�Z��=F�32S ic���ڠ�s��O'�|�B��P� QclN��*!����(��&:^�)N�Cy�ݷ���C�Y��zf}&�2X��9�}� h�G�#��Tȑ�^�D�L��Lf�V ��C���5��|	(�Sbz��n,��X�l<�#������-��X �<{�$����PmJ����H�DE܈sR���P�u	�=�Ͼ��|��~[F=���8�G�S�}�e�7�r�Յ�^^��.?���H�>��f�&w�ܖ����JY����Z:8�:L�j].=}UZ-�jI)F��E]�~��ʁ\�:���*����C��}l3�=IF}i��x)��'Y>�;y{B1!5�s��������J&Sf�Q�Z)!(��u����t���٫W����{�~y�����ŋ��-I_����������]]�u:!�3r�qt�f\ptF�*�/ f�f֣�x�hF*�0�Qٻ�{����C�����G��5�Y�Y�*��tZm���f_�?�4�
| �D��g�j��
�_���!qg�'('H�l�VQ���O3|%����3 7s/]h�eeyUk��/�1�:J�Q'�M��� �'���QM�q_Q�Ҭ����ϼI��3�n�6��#��$@�����T�[�d���'�&Ԉ L�+�<*��`��d1�>��S�}���,n.���~L:w��L�^_[~T���I����q��/\d�1��e�Uw}�C�z`H�YBʫ�湧��_���O���t���B+d)��OCkA}�8���/��R*�>Fe��>9�ٙ�P�x��$�2k����f?���"����0�)�L�����[k���w`���?��l@
q����`4�E�S�p@�Qq��\��H�������.��HQdp��yY.5չ�vgKƨ)G��_;uV��OIiiY���X޻Wί��W�~R���(��ʈH��r�P���ӗd�^�;?����rL�bg�@�lfD�U�����d:��b�nHX�W *W�jH����g�����HY��&��RA/�Zk*��n���S���vY�s�����*��r��,�]�r<bu����}������^�����ngO*i�JV	HK���� t�e�
�bs��"�p�닂MF�r#X��(�uQ�Y��6 �`8��F9���s�B�TI��{�ƣ�E�٪)�tby��W���Wh�|q�AJ%����UD %�+�L�lZ2��r+~�A�Ci�*���~��A���v��� I����]ͤ��T:G�ҁB�t,�{{rtԷ>o̬[�b�h9��!�/��V�%k�K���7�E�������VZ�89_����"b��Cg#�0p����;;���
�_.U�N��ZCx�)d�����j(Ģ�F���܄�(��&�9�?������'tm�Ju
����
5~�jؿ����o�TF��A������Q7�E�>��dD�9 )���T�k�B�ӓ��o�Xk�t�2��\�Ͼ������P �V�95��2�7�?��,���f�4jA�Ergw[J��)P�Ȩ?��AW��l4N\84'�K� ���s����'_~Uڭu�Z���!rZ,�&(�C� I�J.��Nɵ+��L���۲��?�g|��=�o ,<�
(�e�'��X\ZүE9TL�����R����	��~Z*z?�zU"��@D^�9҉�@����,}c=�Ҫ:X�ϊ.�2 �����z���jڨ�x�h�&��A���nQt��O|B�>sU��s����R�x(7޿)�^�o|����3r���Xܐ͝]��A]��uߨ�.Wjkb�Z��
�x,��&�lw��l���]����xr�<6Ͻ甓��E4���b���0���f��<r�j���Ga^�T.�m�@F�q���y�45"��|dO`�ݡ�)Q"{xp�O:i�Z����n�K��:����w�	��s˱W�ڧ,7��<ȏ��1��r�I����
�|^���<xڡ������)�cYd��k(���w�{�fO�Ѐ_�A9��J���܁�|���!5�]�ð���^��D~"a�K��1��
��*L�͵�p�;s��#3X��c���\� O?}�e���G��aɃ��+����n�P/�O��LZ�e'3��G���:0�_(ҡ��n��l�4��S�3��g�0 i�g����\�A���	�{2˶������\�e1�3�T�Q%q�(�,"�t~�d>�:w��IU���k��#]�:�������|_����Qi�St��ey�������v�'�����ڲ<�tF:���7$����@�:#u���(��|M��l�=K�(a4~��˾f�,�g8� H@����E�MZ'c�o樲^�G�Y$NpƱ��^�Z�=���d���JP�pgK�������M9(Dc�q.�������9��"�~"�����3���E����򥧮�Z�)c裇�Y��k�b�����@�(����S�)̜0 �^�l�1r%f���,��07<{d�"�eL&|I����t�R,��J���&���@(bqQF��',�v���l)�&��Tf6�=E�.ɉ:��$��\������> ��۟��+�Gc��B��B�f�|CF@Qp(�Lpj4@7|��Π8��jYẾ���C�����j�N�tdJK��>����hW�zG`�
`&����U��k� 
�h�����-�t<!�g������X����2ˎ{P��It! }k���ݸO�Y�� j@HJ�����2�v��sM�tp�݆_�7h�(Pt&/_{�?�d�`�}LY�H?k�pOFe�E�n >�O��R̹��X�g?���捌�%��A���9RΩ8z�ّS��ZP�f���߲� ��-��3N26O�N�U��L˺�42��(U� �u> ��C�� 4�* ���|�V����E�`��e�i6���r��I�_n`�j��^�ړg�y�loQt���E����	{
�o޼%u����@����Ϩ���{r�7�y�*�~ݵ��}��� ��a_╆t����"�Q3�1q�S�CF9S��N�#���9�d��A��fk��<���_���.�����W^��R�ͽֺ�_8�kp,�qOt㐠ܒa���9)Ы�!��I���� C鷪�UbF5t��`�]�����9+O�'Ǔ��G���~��� �=2c���{��gkQ��)
�A��  ����v-�ʸj`Y3���#�#�D�ȲcTuG����3� ��ð�>D�B���}����Ҏ���p�' ���1���~ZС�9���S��[��<���i�G|~�g�w����P�FKS%j��j���Cp����ֈ����U��-Y+�)�^�L`��MD0^&�($�/&e��@Y�����>��ɪ0^&���	�9�����\�����3D\ī���Sv	�Ā�2S,�b����t\�V��5��5O#�1mN�.�#+Pu���D�������j��tI� )���5��։ǄIjmy�(�g�1���We	9��龞����y�xP�a�������|�����x@�Rܮ�
��pxRk"J�*8���^bm'�8jf^��E��(L�`�]�:Y��Dz�mI�Su��ρ���P���~�EY)7���R�P'm{�ܼ{[t�$�X��y�m4���礥��5M���腅U^���z22�#�K�jJ0"s�q��g�e��K��2�Od�k^0n` ��eW�47���G�SM���1�M��'�ԧ���r�2���,VO˂��<��|�Wd!�����4�5�JM��Tsu�R��P��!!��qn�:�Z.�c�A1E�Y��zF�\A����"��S�� �ᘴ=L�<�5�2#�a�'^a�]���RrO+�����W�E��|�)�s�����E�<�h����� }h�0�g��NS����/�wԠ)p��ĵW�}v5)��ᨠY@Eͬ� 'q��Zo1�q�ѯ0%U�Y^d�P��7À@?������ ��TU�\*�oSC\���4J	f�f�z�%�a���+ �.(��=� �]��V�ɉ۸���)���}@4
j�[���Аn�$h�5�S�Y���u��!nSj��?F���fJf]��6'4SW��� �d�q�&c]S���e���if���P!Ȓ+�l�{Q��C������)�q�
4Ⱦ�2B���� �3P 2N����z��鄢
�C��5#n� d7 �\oP�p��=���	�xBH���X�Aq��y_���h�xmM�Z��~b���{��gy�ݽ�P��q�9�������������B��BShC65F��ز��R�2��Z��q2*�(�F�ұڦ1�V��H��:�I��S�r����w�Z���ߔ�����#{~��=�u猂���5���ډ��K��Ǻ�A(F�*[@%��m�9G.�W���]$�	 |r<9>�`f�HB�̺Ѝ���F�@���
������S�Vd�OX��D�̑�lc`�H�j�>`f	�R�w>�R��
��`!����è� �.5��@�c��;N�=K��؃������VzSa׋�B\B*�sc���%]BZ�1����<���VP���z�{���2mԗ���(n��4��~A�/�,��SE�@�B<(�����u%��ZJx���DF�{����ؾ�8wM�l���>��8�4�`}�S��\�Щ<O`���zO����  \�����7���]4ubRK�e:��uG֩��?����X(���9t�8�q�튊���P�Q��̮��/�3j���yA�+���R ����^����sL3����9�9o�Ü������7�вY�:μ|����P��vP]V��cFБ�bK��R#l�x;!�,<6Ip*���i���"�"ń�ш٢٤\�AN稤���Ǻi����jeLc�;:do�z����ԳB���Ҫd��*8ߘ5xݣ�:F���(���8����D/6zpr�Ta���v.�9��"�(H�gX����gXQ�VUp�d�q6���~9���@�wA�
��A�J��\��ߔա���y���/�'ao�cD��4eA���ZKP�\"%�>���B�����GjSO~�ya�н��D[+![/�����GOA�Kظ�=(!p�٬�Y������T^�2ss�@��M#(��|}6��1:���b��1�s�4�t#>+�����8G�	�O<H���t�N'9�g�\�	��R��Np���5v/�檊�v	U�����d ���)�2CF�`�S��%SF��,s��a��
XD���U2#��_R��ʠ��E��`�}� e�sf �J�(��oP�AF_8�=d�&��k��Ô`�~��J�/�M��"���B�.-�̦:phf�g��{~mM^{��$o�n�e�i�d��R/������rp�>�Xã>��@�E&ʡ�Ĕ~�3���"�N���5lz?P�C�s��f6	��R�!_�������j�l������`[�y�]]�O8���@c��?����h��}��AE����FB�T8%x��s�� �	�?
�@���+�I%�H��<1*/΅F��ѹ�l-�N�j�AgGv�t��f�Yd�1��X�5��kY���XO��7:}c�Q�D��N���a�Hgk�X���T��1���Պ����h���1"�;{����X޿��Σ2�����
�+������O~��u@���>�^�kuA��@��P��<��Is�
�l����=���p겹�y�D~r�}r<9>���?�%�$x��7���`�i|l��)�J~A��	����(W_`j;��L��}��j��l���y�m?���'dL�R�\K00+��`�F����P�Z�+++K�^Y��׮����`oOm�C���nS�+S���F��O�O[h�(�U^x���ǚW���ܞ�v��v��( �崴�>�O,�_� ю��P����1i���r	]�D�l�~��B��D!�ܱ���*@��u���̲�+�J>��rǠ��U,Y�a�Z�x%.�8%ifvC���Lk�6�����%�\}&n)���X�av��/`��d$��̾�J����5L�ga���u�����T���jY��a��8n��S��_S�IDn�H(􏞎S�@�>�����,��n�j���z���fR�^^�o�(�5��kQ?8׻P,���h��f�t�N���b��b��w>�!~X+�p�\bǽ׾����B�]V����'����2��U�
�q.]P=���u!�d��Q�8�p[���֒E�i��g�:_qINE$�a���:������s���h��5�����k_@4_�n��JkQ�����P:F+��|f��|��d5�ѸAaqyy��I����]�N%��ݹ� bW�j�~��p1"�h�Ǯ�W  ��0�����{�Q
��V���-"FZ����@ѵ�]��&��U��Vw�A8�{f�> ��S�
��faf.ciq��fEVS>2��[p �,�w+R~̳��w�VmK����j(����s-BƠ��g]wL��g�/�/\����ڒ�A���K�I�LY~����z�٭rCe��Z��}E= ���o�45���������;)H7s�ٶ�p,�QO���,/,X]_��qE�^��b�M�E�Bd)�P;�5�gO���Aπ?��Q85Ud�u�� �R],�����XiKMms�v`EA��~���|Y~��/�{v�N4p��^��NũRK�
��VW�V��[�C W��@e��o��H�,�n���EZJh��ܴ`Oy�[/Sв����9}J�,��[?������\v�deqQ�^�$��w�}�����5T��ux��O�,/t�����
��D��N���Nf����R\+���k|v��euf �Yw7�P�&�i��(�%,�ܻu�5���Dv�*�c g畕Uy��I��rq���"����|��6뺆�ƪ��F<Nu�����F���"¯�+�2A1ڔ��&��u!�Aꬾ��l�ƃt:���Y���cT���Y_g��r�ޑt�G��[��5e��@�}�@Mm!!y�5��Yv��I��=Ca~�x��o2C�������^�o�v����P��x�k`YB�����zl��
��f!�*��TNȼ�XX���~3E�'S�M�2dv-gP�@��vo ^��N�c%�� Dq���V�&�Ժ�����pA��\�xQz����=kM60H��Se{s�j�Y眺�5��-�L���=���2�Z�U�ꅁm��f#c�����(�{�?��^���Y]nKu��{�@FɄ�-�]��i4��g0\�m���D���A㤮�O|E"��9C����}C��L4E��#��3O�D {�(%��3��SJ�0|ew�3q�J^��f�W(u@�,s�v��GN14c6��q��z�sp���R�J0S�ϨI�=NT&����y��8I�h�(�q������K��v=�����.���C]'�����|V���T{/@:wm��/|�j�x���˚R�5\^�ڋo���e���U�D�|�j���fr�#u��9�ɚ�ϛK��.�V�k�&��ò\>uJ.���^2��/�
z�IO~��T/]�K/���~>�~g�9���NX�5L+�KXbtɃ�o�s8g���>:dŘ����Q"%�Q"��j�(�w�fR�;��!/]~V�j�@�ؠ-����el����JUf��xjqY��byo�/�2�)��8���1H'���n�΁B��9ڭ��D�G��鳍�خÍ�T�^RSg����[_������:���g`��y�"OϢ��ES�]Vd�ͯ��E0��\�9`�����c�|������&�& �lh�u�g+�������ˤ�Fh��]���-�(�G���:�uN`��싯��^�4��up���ȝ�-��:
��ZJ��2���>RG� /� 82��	�5Ad�r��T���r������6X��ǮpF�C1G�y��-y���	�ZN'<4P6&m2ek	��@�r�>"���QI>����S��&�NWV�
Xt|��/�� ��� ��C0r�ځ�.ɽ;w������ŧ�����Of�/���t���������U�\�e�i�0���^]�?��?ԍyI� �Z`��4+f��z���r�z劼���U����;��?��?�%h�*]B�%20��D/E����@	5�	�.^7��!@������nm���]3��n����C��FS�v�dE�)���^��?o����)�p����貦���ؐ<����D�x\k�f�$ �0ZQs�_bQdq,��+�����Rn
�������5t�_|�9w����X._8/e�" ���A�&@��R'���{������s~�:��Z	��ND�+��*!�.^>�w�� (��{��Y���������G��*�O�cV��'㉩~.{%����՞�f�s��X�/페/�}ldK��j+�������}m��l�����VPY���R�.Iy�.���(a���@,+�����݇�w��W�L�T�oR��Î���@��i�6Ij>k<�/���������i6�MB��\g^��n��$�3+8\>%K���	˭��if�\M�Գ���W���]z���I# �wmͮ�1@|֍�4-�f�&��(��ӵ1M��\b%C�G���G��,��^��<�m~Q��S�ǰ�1�
l�XHu�V��s�mL��MY�O�C�~���X�:�޲ ��!(K�1���6\���0�5)Ҥ���Fꙫ���k0PE͜s:]®hz���������� �G�Ṅُ�}"���t'�.7�HD�=�G&r�y����w6O�<��e.Kv���[�^��x,��@�OL�5xca��#ւ�DdE��QU*iYN�kr��*_~��ԙrsS��<���DjӾ���ҷ��˔J�!5�pz�Kk��ZY��:����T�g��h���σ��GT�;�O��t����XK�n2�I�SP�Љzva���	iK�<w�|��+��aG�r,�j��~xG�ﲷ_��յ�򩧞碻qK����{�X�\�*l5/nM�/d�@���1��,��Gn~���w�?�q��ވ1�3��� ��jЪI�(3;h�/��7��~�k��5ö���k@Ǟ���������J�����!����7E/J|���֩���k/ʴ�gK�T��:�̟�H��h8&�=�զhtzT�򬂞�
x{Gz�#�6�8�gQ�u�Ȧ��R�|g���I
-��3ؠ� {�1$�#�U9w�<�t����n  � ��4a��J�$�h��@�>��AO�'׍&�k������`mkN矽�J�b��y Ť\��%�K]7�+O_�p�6�r jԉU��x�-�֋��7���*�VN�s���;7n�ᳫͺ���u��`�b�󵧬�d�ͬ�U�����2���榜Y]�R5����s��x�c *r�~��f��(��	l ���	�x{��u�	a,���3�0����,��1Z3x�P~��}Yn/���HAh���	7q �F�.�F�>����[�g����_��n�}y���@y,׮\�󗟦S�����c@�l/��ԑµ�tDp��e<ҹ�̀\8H�ua~���JK���>'3�h�`�J�jϤa}�aC�(3�+ ��m��(�럺tA������oܑ��%�2�����,桮��ņ��d��g�^�$J'��0Ɩ�W3X:nߋc�ą�̎��q��zr<9��ź��R@2�/�+MA�4/Q�?D�O�bӢ;_��Sc����zo����'`	�~�(J<�����(���L��(�` ��:5�=�B�%+��hЗ\�r�$��E2Βl��P�Yc�3dr��	He���_��k#�^�΍K0�>���@�gC��"Z�1�����@IPgk v�]k�"πah���'��3�#0<��T�a�8���3�ɱOH�,�X��`�3eVmfyb-�����̮B��<k�+����G�12b���j�|���:R"�Re\�K�j�N�a��);>����{�[�x{)�J�_�(�Q���<�ɀ�`���C��dDf�q�uv5
�Ϡ�<.C"�Z0��N>P�������"z�g�e�
��ޚf�Ow����#�Og�ι���Q�
zK�20�]V��QE�;̏͜�b7�~sJ��Y�E����{>+�3�3� ��t����S���|^tV�^���W���ή��qC��ې�>Ժ:@G�����{�t=�h ����~&_����K;Ys��2�J�������l���G_#������/����1\�M���(�Q�
��W�_����2�#5@����������U�:]�����<�Qd]Xo"�x"�\y^"lm�7ޓ�5�n�sGp�W���������٤���`���Lm���L���l�Q��,Z����d

!��2��'�:ݤ.�0Tp����I>�d1s���ӈ����p�rO�>��f�>��f���l�򼳵%���<P@x��EYi6eptD�z��ii_Y��aO��>��h���Ρ�|p_v�v���Ѧ�3�h����xx'�*rΘ�r^����I¢�H��:"��R~�"��$ν�  <d�pN4��B/h`��T&c�v':��k���T@���T����A��֒�/+�J�^q^ ���E�U��Z��.^�yX]2Nj�'����v��y����M����W�9�W�p5I��Ւ��+uf�IA[�r�C3pAl� �S�[��#�fM
\���>�Z͟��粳�-
B��edA��{饗�_��Tvw���-����s�e�Idu��U���GWQ��^Z��	��@y�����(sX?{�A�{��H� ""����?5So�qB����;w����S�����G���@7����QF�H٩�B��7�s�NZ�ʲPo�sϼ �QOv��:��K@�BO��YB[�F��E� ��)A��1���El�ㅍu�hl]��߿w�b4�m��Xfڥ��L��40�E�s#��=����)c�����6��t���B{y!����O�'�����	��D��4��kO='�qE��9[+M��G�{���-F>��S���� �� "�뭇�y�����I52�$�bwlL!�w
j>��U�K؍��e9��ܺ_��ݔ��]�1���=����z\�}bȽ �
��Ԩ��S&�������g �D[��5_K�Қr`�Rb�2�L
��@_�7��Ao ��}��ᇒ���l �]y��=Np�O�Pka��S�d$f��؄$�D0��{<2y���z���p�������ܥ�����<"�Z�rV
�$���z\�_l��z���Qy7�T�� ��2ƈ�)��VK������� =ӗ��$�[y)�NtҡL*e���#te�ǡy�H0�����W���Q�ܯ�3��'19R/Mam�|&&���X�B��g[d�{1�YfpN,��;�����:�4(@h�.z&�_�����k��~$S<������̃Yf�#��g|�b|f���Rֺ�V�Xq��iI���֙����h���ލ����ԡS9���Y-7���'�ɑ+!i��.Tf���8�ӄ�%d�jr��p������?�Q���;��/����TW��~�dw@��Z��V�Ea����M��ޑ�,'�زa"�u�u����l[�:���z����#p�1Ӧ㱟�?��*���!ǉ�)2��Ϯ�E��ޑ�ԱD�@����z���ؠj�Q^\HA)��f�Y��%��ь͓�h	hPqL�����c9�/r/�X��a�r?2�ɹ��-8�I��F:�$;G��0�rM���"���"Q�c��Hz�u������k��������������겂�uF�@m��._�$����pC���B����!F�F-��iД�C �b��i��C�M�u#�;=f���E���"t���~;w�[O d܁��6�FԢ�>����td{_N-���t����dD�.�1�kC�*@�n�G��ƨ�5x��K�ڞ'�2NLe3�utz��~O�> MY���kϿ�����Ѹ�+v�ڌF��w�ϦFP 0]"�<�Pl�Ν�+O?M����C[���#�fC��? ��Ӱ��`"������r��]ְd���	<!��b���[7W��u>��> �`P�:ߛ�퇾���{rJA����j��1�P���D}r��J�1.�
&Gt|��K�΃nϲ��^(�s�RX5��ZC��K����9�jM�r���e���7;�{�lOu�!S'����[g���zX˞��**D�BŘ�}2kM��&���\� "s6�q���l[ʨ�g�y�l@����B��VM �I��R2IM�*0����'x#��kyr<9�~�Ms '0�8����"�~�S�ĲיȮڊ��t�]�c֓C�j�M�XZJE�D��@�;hN��K�Sڃ4ΙalV"Yj��w�'�d�
˰�YD
�DA]��.S 7J������~_�B�����ڍ�+��ϼSk��x�&�,z�UX[E��R0&/�[�r0XF���{�jϨ�Pr�~Z@03�M���%9*)����q�O�[���¿s���Wx������6�x���$Gh�J@�,TrS����=>����ї��F��%(a��b\	��J�,�⷗��wΝ:��g������v�֨�k�ǈ�ڞ��ͭ�����y��}uxte�L�%�k=I�u�,�Ka��̉�����>�Il [�9_�&1a����?��	޼��~��Sv� BD��ls���wƘ�p��M��5�t�<?���2Ԉ��."���ԍ|<'
�U�bs?���)L0(Fs͜\�:|vQ�Y}#��&�^豅�n<���z)^���G�^)諪ـ����ޒw�ܔ�r[�/�ʵ�O(A@)�k9��&�����ݐ_޻)�]uvt�Wpu��EYmY��2�P�N�P���� 0����쨋��m�@i�Te߸�QO~x�-��?��:�מ}N.��g�s�g���6W(s\k�	�>�qMx4=d�����&K�:��;<3�f��c�OsO��<��Hf�`c3XPv��#)&RJ�=
��^v����Z�%�A�U���>�a�:��g� �>QgV���ou|)��G]�zYF5S�e��@Z!%���ɷ� �!w=�Nޥ��E���`�i{���h#� �?���t�k�-A�./*`y��%:�o��3��[o1�p�oߓr��ڪ����ӗ/���*i��r�䎦�V�j�|ă@31�0{��Zl�j�����������b�)�O����Ͷ,5y_%���I�Vj��������e�Wj����Oeok�{7u�+՘�6 B����3����oK[���b�.�ۋ���?)����Y'�A(@���5�ώ��:qT
������P>x�<s�����Su4I�'� ��:� ��	�Dd&v��?�#�ziS���Ҳ��ܽ{G�����+r��777	�q���������r  ��IDATa���zB��A]��G6���k}��tQ =D~���k�Я�^��ֶ�P-W�A������~{g�4ߞ:;�Bƨ	ԯ���d��<�k��Ԟ��7fm5���IwW� ��Fdy/�
���/=uE�^}AZj��we�ӓ]�CX(P�"'��&������/Ҋ"�Q\�oc�\D�'ӑν��ˡ�Չ�鎝B�Pm a�z�V�!w�4�^�#��/m�˸s }Й8�L� �|b����� C�������@*�`��<9�������X�s��`]{��$����ew[���䠳'�Q_Aڐ�X}��ຨ�����=�wPk�6�u�~M�T��C�)�p�|��&d��
�kQ:�sГ� �0�r�%���I_?�ރ�uԾ�� ;7U1�=J�Μ'HK\o�%.�A��]ԋn�n��}9L�%��}�T�`�����K�Zp�c	6�F�u�A��>�LdJ���P�G��i��Y�[9��P-�ի������W�?��+)X�ӉTtkP��&S=
k�2��&��?�ev�%����z��a)�%q%iƍN=(�]g�_�4���˯��_��敕�ca����|����;�Λ�>h�{�������g;��K��r2�԰!��qC�p�e����uX�P@�|@sn���eg�>�$ ˹+�w�p�	�@�{�5o�$� q�%Z��Y�է�C���+�Έ�(d1f ������&$݉�+6�@����H�9��|��@A3�EJ�㑃 (O�B��'�1�0�l�O�ݐ�d���7�}�������+h:���-���b}ji]^]� ��e�`��	ԭ=�xJ�[m������/y9��?dW�
o}� �X��9p7?F��0A~��s��c���G	MRk~YA&-˩>���yw�'y'�ۣC��.Ы��3�~Z��l˭A� oj�7
Iуo����!\��<@��z������:Y��q�y�Td�������� �2'��a��#�ӱ(ӂ�l_�t]�X�����4RC� 3�%��������L��ҩ��ά��KuJ��Dx*��wZ����L���
x�@Լ �_G��լD%�VX�Ÿ�6
��K��sW	h������u���.�P�o����o0��������&��<-�Ϟ�F��ĥL���M9��̰�G�2\Vl[d�]k!یN�;b�4�2�!2�hf���'��n܃.�cl <@��e&�'O)x]Z^�]W��,�P�e҈eG7}���U�!�F Szߠ�\�|Q�E�T���now�b"����@E�--&���c8&��ܢ,���6%�A���w�#?y����7���"?5^�)G��bdB<8���s���y���ޮ<ܸ/wn���@�&d3�
�~�Pw-�cj��n���ײ��dT�� 7�$Nr���$� ��b]S)v�6�u֦"�\E�~��3X��y3lJ��ᩄ��@�n��m���@��DFh�[2 �R��gX	��h_����������1�&��^Cg:�gP��i����מ��R[tde���  �;�@'۰4�q)!8�:J-�m�V����At:4�\�~�ه�)߶[u�h�yxWbu`FT�:��~69C}f�й�VC)�<jUcY�qj�G;9���&��Xڭa����ٌ:jA~�8+O�'�?��#��Ή�'�H&��`G�nMh�^��ҖJC�ÕE95<-�^W��d�`G��߫��^-��/L��Ju�D��I`�t�7�o�h�S�J_�2��|�EmY)�Ն�/�&ԇ�'�����Zf}����d{wKz
DG�7����5!.�௟��?���Xv��b�gP�7M�����7��\��B�,\i�K�������gW�9\�2K��=�,�c?�#8eǘmL�`��S����K�a@p�	������ek�j��������Ǌ�u���"�tB�oƌkM���eĸ�(+��FPy�����h���篼���^z�Kώ� �ؓ��j0�}}���������o����A�f�����jW��0KC��J�xW�콍��r�L<����N�Q�y���]kf�T0N�.il5 �[�2$���$�vM�u^�S�/O���e��k���8��`����d� ��!h鄩M�|a+�R�2��gTe�(/��A��(OL�	��"�V�*e�B�๿�G�?N\�'o���Lw '���.r �*C��A!�@9a��*5e�r��ɥ�P��ʄ�h��ߕ#��_���|����P?����K2�����vA^����p��e��̭�&w7囿���L_�Ӎ
�	2��IXy40���������^3��z�w���ؘÙA-R�׽T�K8�݆Ȧ:��ݗ�7�r��䓗_���5��<� G�����)�bd�B�A"�ِ�
�lBc\G�4� �'{��|�'�9�����y��n�}gxJ���)�E�R#<�}�^q�"�rd���Tzy��Yh���@�OC�z4�`�H��C�� ��)$�&ҏz�Q$���yDK�|~�c���[�Zf�/(�%4z�����ǣsu��!��*e�Y����8�j�j�{�]y�����ؖ�����&'���	G���[��H>| �x�u�( �B���&2J�QFF�g����Ə��=����0ru�9����Իz�kԐ��}�ܹu[v�v�����M\&fl{wG�v�ޕ�3����+��~F_� ��:;���@澡�8�O%���vS��z���"�|"}��C�HO�{?yC�[۲��dU�s}�6A,"��f�����Q�&�WeswW���3�P�K�^L��z)B�f��}���ϔ�APQ2s�������Q�e�lnl0{���^��M�!�*�4�3��\�;7����)�}Y#_� 0:�f�)��z��F���V��3���u;����3�֝�L"�|����Q���H%�(^����_���sKO���Nk5�%�t��+����n���ޫ��o�U7Ne/����U���@�ņ<�y�o?�Τ'{����8aˑ���Z+"�e���z�h�� �X� 궢���t�#����[ț�aX�XȲ�`-HI�G"TF�:Y��N!k.C��$C��g����Ў����M�?��W\�G�y�O�{�܏{ٯ�f˯�����}��~�h+��2����z����V�B!Ŧ���}@�~�{��u#yU����\k��bL�Rn��ր��C]�#��)���TT,F�+UmڰۗãC��mё�x{Ւ4�d��g�ͺ�Ȯ3�}b�q���PԀ*Vq*�(�E���z��v����/~����ey�������Ԣ$J"��T�Ț�P�	�|�qc���>'��D�BU�`/F1���{�F�8g�����M!`iD��:���l��4�K��~��WE�`�#�G��,�l��q����ׅ]Bp��}=υu0��QZrড��3�.�G�X�~��t��T̘*�wlD�@��|���B������t��X�����J��wN3	����+A�(Î�Ѕ��K�����EspP�����������_���g_�ԓ�u�_]�PQ6�n&|=� �������A�_�d������>v~�	Z�gg���*;t2����kJ�Pq\ޅ��@%�G�Hn#K���8�B~��t�x��V���W��Oj�7�耧ذRx�B�1�|&�F��W�=1���k[���>���{v�g�j���3�n�z}��J`�Vթ�F�\�07%��lN��Li�����O����*���:�?[�8@� Àvz��[?�ާK�:hzt��ƴ��s�M��|��s���^��}�֕7h�`�_:Av��3�����ߢ�]�Ƞ��&��
���[��e~�9d1̀�c��c~Y����~f�AҨݠ�k����}E��.ک�8��Q��q�vߚ�͸OW�7� K�{f�F*,�<-���Zr@߼�S�8�J�����"-5��H?`��^tY_WLUfO� ێ2/��>�\���RX׺��M���-��|
�$h�z�3��9�� �3���NL~?�
;y�T��Q.��G-Q�,h0�N��f���wW�~vF������,`�%�x�g�4��j c�N��t���`��_p���6�w�2�}��u��~U�����������ߥ��?
��l��2����@MK\߽�K�T��M��:Ŗ����wh�Adf��ϛ�p�L���q��t8�R<��[t��e��y�������&��2P�Q$e�)�Ø�w9 �Br���2n�
�B��vw�o}�N��XXK�m}�)�P�c��ŵs�mw�le"1�
X���,�� �g�04@h$
�1� Z�
�r�6�$�� ?�Nʋ:���� ���x<$�=�*y-�}+Q��`,���HO��J^���N�n�����(�U� �9���n������~O���=�s�\���s��1�nK���4��wDy�H�|�#��c͞N��6b���݃� �:��e�m�Ј�0a��� ��/���y�nomА���:WgP_(�/�����l)��잖���c��4�-�؊�&i�����AhVӚO��J�T�AQ
��(j`4H��i�wܥ��X�G���t�bj�[H.Jf񕪦�݇��T��(,��g^g���/���{�M����~ຊ���������P�������q������GM���<X���>J�[�q�5)� �`������`8�,�3P�	�Z�U%Ec"S'T�2!k#o2�BЋ$�j-� ��^�1�d{Z��dH���O�)-s�9j��nA�yyEuZ���o�u�}Y��h��ZlK1��<+�L��%�eBN��7���}^*
2ͪ�?PrL� g��JS2����uD����ZX�)�e>3����(���^-��L+�AM~dl5n%�,l��HZe(���F��O]l�[.O�`Q�g�� 5�&}޿c0�V*T��i�yז���ή��w���+���5�(�=W���[���F���}��0��A���-���`l�T'��HeR�<f���^>r�u�'V,t����I��5��J�Req�񝥨~y����`���z��h�Q-I|J͂DUcDCI��,l���ϼ�^�����'^���o\۹��C�}b��x�NPY��Ӛ�&��Cx�5Ö�	�t���©�X�e��>̎�:�d�(��$VǴ��i��tᠬi���?]z]�ָC1@�X�؉B
���}�~�qQ�Z�LMv�t�ۡ�ߺN~�Ę��#a�Rw2�N�Ǥ���Ŕ�Gq��h{=�JP��J1s�G�Ʊ�����!��{����ԥ��K�ڴ���}�����a���c2f��sps���< �����>u/�*"ۈ�Ǩq��F��NȜ@x�3r�H�����,�qţ5R�ml�	�=ʵleξ�F�|v�
��TC�6�>uGl����R
P���IY�͢`�7�An�M�\M"a�����S�p�b�13�3�nPa�׸�Q�����$V�9��@"�?X ���v`
�c�c�e��|Oȏ��쥔0�m�X6N�UE{z=H�5k6�!�l�0��p�΅-}�3Is�K���u�v��K������6�ךU����?�.�;]^;��6Zҳ�{e�76�I>�y*��2B�*li�ʁ��� M�<�2����a\C��5G�
 ��}�@*���SB��q�g�b��6�ɘ><�jP;�Q�l�<m��� ���� ;�E�W���C"{�\ɤ���9&���A�009{z��-	�����2����Zc����-a5F����J���c�' ;�c�;�+xnn}z��'�ǯGv�VPz�7�z�{F/�҉E�X--/���ʚ`�ku!����A'*Q��"M��Ŀ����#��b���\�7q�K��a�s���Fw���D���8��6�__��F���P�׭+iY�yO�Z� �Gd�Ǧ�y�>�@4/C)5C� e�¢�Kސȹ}	4i;D.s��l�c��EM�������;,��Byc��P��}�y>w
ynT�
�~��P��2��4�6D^iP
��D�|�}�dۇ 4E~�{�IGr�`��~����wY� |?ǯ4(��c.��r�{B���.�� ^ Y��~#S����?�R�ٖb3��>�~����`$�[�?�8�� �>�zR�?n�� D�}�{��.���R}o�V�֥��F�]�J�7��5���mK�@u��4�S�׋���H�򼲅X+:m�Sj<A6̭3o�V)���fm�g�#�i9�3�e�E��g�)�����%0��O�v	=��VM&Z�"�*���i�ŭ�:S2�k���s91�%���Z��� A=|n�|�Wc����Yml�e���_���}�~�O�8���xq��k�����#�7հ�Ճ���I�9�@)�4P/YNO�ݵ��d����5-GSB
)�B�7A��I�.�/�-�^Zk�]
�p���r����}�;�A��]|��ؽqc��w~~��.mo��$(�o[O���Ǎ��!"��A��&}�d�H�5.�7�I�1;`��"��:VF�)����rb�����)oxt���	��$F +x�f�*�/Љӭ�Xt�R��������a�7���&��B!�Y��C-�J���ѱ���ƺ8��2|�#���z��:By��J�eTE�!�`�[�|*��F�R^�3@16�	�S�){���q�2N3��p�y��"e��{W���R~%⥅�����#W*�A���
�
[~0�BJ�d�ٜ�&i�1_Ae�o��_���;��MJN/Q���"��������e���\���[�|� �(PQ������i�7��L�5�L���6t�@�4�����P�Q�Յ%:qbE�plF(=�u$�&���	;�׮^���e���N��jIf��Ȕ8*W�1����:�t�J�0��F���2A�z�<��9Zl�I�NĀU��sK(�����.�B�~g�v��h��MA������A��@�6 � yg������C�������҉���u�&�:{V�cĀ�(���f��[aMh�����d���=�J~�����It���i��s�!���¹ȥ}?&׈���Ȧ�/4��㧨ƛ�ԣjC�u���൉�Ԡw������ߤ����؄�rpZP|"r`�C�k���ܨV2yہ=�^Du�J��<m��q��҈!�9�E�|�O�b���J�X`qX��17SEuB��Xd�
DZ�A0� �q4��?q�(K3�N��5@�4����"(�� ����3�'�ֆ����������G�p`�����E������L�l���*�$�ꦷd|�9Pfw{����,!S@�
�wy�!вX3:V�w|���'W�2�����vTi3_��;��]|�4H��|��:�Ǽ�܃���'�� �=��w��C{����E�_yQ��W@�5%X��C�=E���s�?CF��پ�!�k-�~4z�x :d��'a��y�Z�5S����^��$�x��x���d0����8�a:"�R���^������IeSB@��0�v�gTV9�8XG�1O���������l�d�pĔ��t���rXރ2�o���3���fV���i��SUadU��-�&.r��^r�
l���Q9��8��-��d���u����7*�g�<�����|���}�`��]8��y��}ޟ�y�:���/Ű�G���aJ*QA����B�'�	4���\��ԇ.���5�ZVl��5����ʏ�s�N��jf_�;�n�fi��n����[Kћ���K{Y���"K>�H�oD~��9Pk��e���ђ�xe���j�������a
*_���C}���8vQ=��r!dNxY�ң���p�z�uV����%�H��y�m�A"����x%�Cnb�@hZ)�?%�b׆�qv��}�ho�rͪP�� ���V�C�� �
�\�Ai(@�Bq
��
G��0v%��D�wܜD2$��B_��c���+k�2��8vg���D�ɳ�,���Sm6(ը$E���}�0
8}+1$�h(��`_b �5B�|�>��3lܗ[�_nRZ	�q��	}�m�G!Q���~w�e�K��d7:��k�-�f���$��C�����#��h���x���/����n*�k8��Q�J�(��hƯ��hyq��]�N��lJ	ʂ�\�����x\@���jɆ�,����ږ.�-��J�B"�p��^��ol����}�_|���m!�A�����g��0�4}c^�K+t���ꫯ��N�N>q�������.�Я�ϲV)�j�Vy�ש�Ԉ�i��:�~��IS@0��~�2}�7����0X�ku(�U�1��k�@���D�9I�w�<W���'�=���}%�|-�!�9��(��~E�`�"� < ��*�x-!#ȎLo�HOl?鉔Z� 8³`��1���~����7/}��\(3��e�(3��:��3�z��)F�J�4��z]X�Sv`z��-D	&J������7!��B�N�S*�|�+��B?z��"�L_2N�bND���� �	GjDC!rQ9_d��K���Q��a�PɳԖh
z�h�h4�Ј�3�P����_��t�Ά��֫��y��L�J� �:��9s�{�xr�U�� M$��{�^怑,�d0@D�c�2���T����"D��/�r�k���Xy���µ%LwR+�u��w
*�R��g���d��=�^!�_��4 �+��1td���	29��>e���O��ʂLϘ�É�Źڜ���2�!�_�PĶ~�{�n�Vն;hv���[;7%�*���	��S�I�_�ߧf�"Y?h���"K<C�@��;�_�}-���P���ϳ"�V�	Ct�`�kЊ�@�}�[+�$^,h��E�Q����8�âk��g���>�km:� x�Aud��64���a�v��fC�
�J��jf>�y*l׫����͓E2��qG {��e�vb|B��T�4�w�j&|m����Z?�����t<w������7�����N�'�|x�7�؍%���!4�(����3���c�ٗ�{�Vg�\�Mn�z�מ�?��ӭ�WV��ݕ������Gz��rm��W��������\ܺ�_�'���x�c	_L�
*I���yƲ���:���:d��3���o�p#h�;�8e~na�b� ��XJ�
�B�=Q�%��xy�z}Xpը"FE��l�\��p�L����ڍ�P�?VU��=�f�>�I�%�9n�
e,|�C�z�	8D�����e����2�%����ߙ:U�׊��L�d\�;qi%0Q�7���;���أ~B�E:����lzUs-ճh%�%�g���5J��A�5��B4�w������L�ѧ�Р���`�I�\�KMj!M�f�m�U.��,�f�[C�,F�~1� J�X2%�}�@2)6�U��1;���O�&��(K�}��=�2��|m�,C&#A�e8f�˳$<�lL����6�nJ�$4��$�x��C�0����"�0}cvV����+'Y��ĩj�_ꉆ[V$|α�s4ݏ!�n��dm��	新D ~�Yd��5���R�;ϛ �Q�A*2��TضHo#��R��ıhaF��@B��'��L��h������gP��\!�B���Dz�>/�����?u;]�v����2^���ݠy��@��X�N���h�k�A6i����w腍�� ���qx@��sQ�X��y�F�J&�׻��"�(K�焲�шzM��#��؉ ��G�����/Ai�����F���R���ϝ2����J�bm#�`��@)�;a�Rɰ3H�+�$��PHz�UR�q Q*AW02a;����
��]�+B�N"���Qf�ј�>��&o��v&�lfo8�D9:�<�d��Hm���"3(=�ʊ+�<�P��=�y�4O�B�|�����?�0�3�F�*��&J�p��tD�u]��E��g�0H���В(8-�h9j���$������ �o�\
�2��JcX�{v�ɢ�FE�9> ���?S��X��`���C��q�!�/ �����V�X23���5Xxso����[t���/���EZe�8� �ɀ�� !�PV����(
H=�^�d�
�d�#	kj75�[K4䂠��{����u����>?�p�h�j�g.6�h���-�◅��Ƙv8��.�%ي�e���Ve�2E��ɋ#����r���$����c��0G��љ��ܹtvyM�ݚ	؎�l�omnл��eգA_��ͤ�&d��`V���V���R�������/Ұ�Շ�mE*�"%�A��5Ӆ���?ξ���}�������>����W����w���&M_Hk�i�6w�H��$W�P�%cz���W�l&D�i��7�auG	�Q?��f���3��d����,=�������/n�c��7N��[o�~o�I����<;�=o ZYW�b��[@j4U��X����6G��涱�!=)����?�%���ϑ9�
+�D�0kA$��eU�
/6F��
	J�=rpt��x5��p��.G&
�G���Q>0�ER���pc7��_�#��gK���`ŕg*
P��a,,�meU�[�v��إ�˳�9��%`At��i�j���C8�h��_cϔ*,Y��+T�
8f�����(r��uT4����Ԕ�9�{5Z�
�8C�:��Pa<p~8�@�4�3G9�} �
�3�4����H��q&Ѹ�A_�`'��ԈAa֮�%����k+�j�5�h�g�{���f@�� ���"�䓅ȚՅ�5F����G����N����`�k�7�"�{}ɾ�������'tR:�2E���$0�`E�#;ֱ�y�	�H�5��+lz�n���NZ.,����t]c#&d�G�M)����} �A��G��7�QwD)���)D�'�12�	����cb�`�<�BVN���ܡ4
d�М^��#���{�@�һ� �.A�L�.����1� Q��}�{4�t��P�蘓h�Ei����a�E5���Q-��D�У� ��*)@�
Io~�aN&C�.;<��l7�����xH�D���snT%����2 T
�F�Y��۪,fǥJ��H�J����}�+0\����D��T����KC�;}:��x�Fz|4�/�T`/%Q99�4��X65ߖ�.K��8"�3*���ƸC<��!����?��8�BO�8�����U(���eK�����4��!��e{�]��I���2���xM���ԚSp8��xM��Fzb�T�aW�H�e^������?�5�==�@�;yƛX[i�/0��7vc��_=Z�p���4���Į�T�������ٲp�u���?���j�o���. ڊ����?�������_�B��0�xLu�r�������l�n3Xo �����N��i}��-,��C�Z��l�o*�#�)��ϝ%���6�g �Hp�Ti�1/��mrg�ݦ��IT�4kMZ�L�*�����h0��5����:�?�M��J ���N3V���&^�T�g�v.��U�%����Rm�ͳ��j$k3���z9��Q �V��s�_��^�����]:A�/]���E���U g�O�OV�gΞC�m�lS��Y��������jc��{�-�k�fXm-���u�f��;|tp���U$�UT<�Q�?8w��7������@��#�����[q��;)>�MG��H=\;t%�����#;!E.Z�g�C���|��bǵ�l/���?����/�~�g�A:�����q�~����[[o��J�������o���8��%�G����z'�"�t��H����l�}մ��Fn!J^�gQ����#m�@�^#�6�sKg�W��	������b@%�X���h�ϐ�Əd�-���G�������}�˂�=+�����xN��̰3�fd���<�H��!�T�N�O��a#(Z�J�)�Ao�m>>�\W>$r$8G�l@�hV��������k��*�/��8*#�Nt^��k�l�}�gߜI�B�J*�qx���Pށ�r�Fi+�qňШ�H�y3w[Pi4�F�+k��üAM=����4o�t��:�Z�N����}�޽�A9?�EvTѓ`�1-�!���3���Y����	���;���ktgȠŎ��`�� �=-���is�P�@��r}|�)gɄD\R�Di�:2K�I��XJl���Z�;�&J�0S�+�tn��3�L������T�l��l=�u����e� f6�!Y�B)���� ��n�ޔ��z�N��~V��3|8�F ۻ�|�-�D���3���0� �����___�� m$��ڨ�H:�i,�	��ǈ��W+4��p�,q��:� A)"% -Y��k� �N�6{~>y�c
�2�*��i��[X'�W 3Re�9�����uiq�IWv�)GƗ�.���c��܄�w����1z����(���:�@/~��ܳ��Z�I�a�FDA�%�x  óI'RV������(qv��~籮G����_�!��}��JD�z�z�.�<����/}������ @cד��#b����\n�wA��{%�F��ih�����Ya;����:՗ɠE WB*l�}��Vy�� *#PJ��$<$����l���-T�H%k����xԁԉ�`�D�_π���W޺BgϞ�����N&�-B�n;T0o���N�3��s&������=>X6���/�p�����&����w���q{h���
��;�m���_mR�lQ쳿�O�]t�+�Ǜ�����|SX�[AD��y=�7��:G�FS2\-�R x�}����x� ���*!�)5�mvR��K&���d�f� S�,@Bi���hggGn]$��;WQݱL�����%�Y�!l,�߳<�&	���Z�k}�C�U>[��(p.a1Ϳ8�]O�� ��;����wi�R]\s��c��'�����ѫ��P���!U�㢙|�i:ub]�qP:������W�}r(�x����C��$ꏳ�z�9��;����_�Z3k�ln�e��v�ɗGQ��8�Ԇـ��S.~UX���Y�.��Q�G�	*6����FM`.���j������O��/���i%�/6��7�/VW�7������/F{��������k�oc����Z�,�|.�igT�I��1+PQ���'=MN��t�����>�)s?����h������;�}vn�),z�fш$r���:iS���#B)	���޴��8rO)�`��)"r������g{Sݗg��qR���!�,��J[lgZB
!��f$�% �T ^�����$+��i��s��Q�#��c�� N����.,���~����ɳ��� Ѳ�A�iOܺJ���+��h��
�g��KO<C�ůH�D�R���]�}�����D�]�9�{4B@D��TIC����:4��(��5�l�nd� 0R�%��@�۠�4�R�)�8�'77�^��$`_���FR�`�|ʅs뢙���� �Y�����d�<ߦ���db⑂V��Y��4|�C��8��ev��N�ӕ���6�-9en��,��B�}ds�U;U3?:�����n����\��������0DU��ꪔ�lll�6!��vD ���O�� p|5� �`�	�T�zRP��>K����h����v�"8;a��V�^k��E�:�s��
岃~�z��c�$+�������"c4`��HHr�Z�����I�0g��}�Y���È���E��g|ْu+�:��!1�\ʕq�aA�Szo�����;�(*���<O�C���uj0-�cɖ ��!�Rhp c&0�Q}C O|pO@�*q�,����w���[|c�'���!
RT�H ��޿1�y�W�ɐ��뫘%SCyZY>I[i��Gے��I���B�(���o^�S'�苟NX}�̈S�F�%@;_ �����R]�ƁB�ˍ36���{ܽt�g��/�4�	������]���-)=R
x��X�&�Գ������@"��������;z�Q �F�D�/T���Q�mEܥ����j���U��m4$�8�h��`�Ѧv4� %��j���܏E�F���OJ+��WݞT���b{4�����Au!�IR��{��?-R`ۖ���Ъ�dQ�ΐg	d\�W�E�r������"��{z��?��}� (_WF����eBz�_��p(vA�UU�j��U�Ф���b-?��ģFq�bc��~�i:{�q�GR�s���V����Q �8(b!9�E2��}�5z����<���p�7~a}��:�9�\ݺ�^��}y�T���Uj�|L�Wc��6!swa.Asmc��<�"ʃ�Q	 {�¿t����jk��/�g�K:�[]M���ş�����������OO�mQ��mJӸ�j'�!��c �q��4J�L�MSC�����<�0�|/����Z|��}�qh�>\fL�+��]A�bb-3��!AR\^L3Yn(����<�1���_��Gw���=9��:aiGj�{�q
g�#�	�OZүO��<KJ��G�����y��8ʇ{��Uƫ�:Z3A�h��Q׎��c��>�zJ���:���~�^8����[w �Б~¥�y�������/�5�q�]�V~�S��?~�Tec��{�������\^��kk��%jUj􃟽Fwҡ�9W�D,p��јg��n^#��b�A^B�Fi�!� �)�8K���}�==v�Gq��v~�q�d�PN#e1 cb`"�u�'d%B�A��Y�iW���OAJ����g��CW��K�[�Dc0�G�Qԥ\��\E�P,}����[]�N�^f`"�Oi�d��W���Z%����ERb$�� �.�JƱ	�����g��m>��
z�ܹCM�.2���g�n�梯�ڀ�c�o2�KD�Rfs �s���Gғ(�3pT@b�� �ń7M���W����ϲ�{��O�<��*��y"�߰�&�zD{IF��?���!���Rw�ld#�=Lع��@FX\(Ar�����E��sdnqA*F�A����H�C�5/�B~�,���p��.,]:�㼟�i��O�z����d��&c�揾G?���,�@����.�}ɾ��  Q�5٥d"o�@��+��O���y2��a�=�uv�F�>���'�Q���f��%���4�X��`�ڡ�3*%�Fz��à" %���^#�N�=x��Z�u�M���Ԟ��>�ϩ\zh=v��@>K	e��SIO����Fg�<�|�fs�������̳>��ǟ�t8��1ڦT���>~�rf��KO[h�
Иm��Kih��;�=:T��J���h]���4PhxO�b���w{�P�;+Q�A�2��NPȶ�Մ��>�(�H�����u�$���}{gO��3����`[��6�LX��p$���(���HgV�V-4Ó�)��0�z3k��x�A1��Z�p̀���ǂA"S��`�Z�r��=�=��_��N�v2��%�K-Ah#��K?��Fg�O���3���u��`��{�!��F�j�1>�m4*��A\���a6~�K����G���lw#�oV�?��`��~�Dc����n@�52��#�z#��vv*b��;����3�,���|�������':�K>~�̅�����ώ�;��89�`%��k����X�7{����F�J;�j8˿��=h�5ǽ_~<�@�Ц�,w�Fqr�G��9О0�|��Z�eTBP � 6�f����y���y>43�<KQ��>\
�\���,,3j*�5#����s�I�'&P}�w匢��r.�(�y��Au�x"�.I�Cˡ�d`dz���������9:�Z���.��W��kiwԣ�f�V��O?�۴��H�O�����GgV�>�"oX���^�7n\���mJ�cZ��w^�<��o��g?E�.]��ɖ��Xb#��O��;�\�2�G��dXv#]7�X�-�Q�*�y2�����2c�Q�Rk�m��)���SfWdl��\K��x{*A �Hh&C����i	�`���H��=Y��+8���]�͢.}��~WJB'Rުپ�F�]�,0���Y<�P�P�2B�^J���/��{���t��m���?�/�����5��7�A�gN����0 ��!S1H�5�?�sxb �yB���k��e����{`�T��ɶae�Z��j|H�c��P�ӔMS� ��fc�?��j�%�Ԇ����F ���$ϋ��>��w1<Cd�/^�"�� ����=�`�k��3N�3e��<#������ ������^) g+fpB�I�5�����=�x��wo^��W���1��C�5�9	"'U�(����iZ���ֈ��dW���F�z1����ȫE�HI,c��j!=��
?���{ l��%#���r�®y�!��G�!��}z��d���>S�-%P��kks�w��O?����-�RT��YM#eb���T��1�e-N���sa���wonhԚ��f7���g�@W���{��}H�����پ�C�~4����q<K�M
[�m�q�*%�R�@�	4c�Y�@���r�lݩ0�&��"�`MM$Zd۵�?�x��{�ct�q�@���@uM�i��K�G�,$�+��ʆ�e���*Prm]�>���6E�V+�
��T�/�L"�+1~�j�2[XV�yS�E�f�`1�<'_�?���T2I���&�8�ЯE���lQ��س��1��d�~5м_�ҊP�U�����"��T���5x�y���'h��[��mKta�k<u/Oj������^����|���X�-���ڍA��6��L�7ު�Hv �"�<x�������\IR��{~ i���3�7�ZZ�ƅ����)��̹�;w���n_�~al����K%m+!� �ގ����|@�f�J���D�>Lb��ڇ����l���C&CoZV �����sY0�[�C���#`��0R�"�238��8y�����X�FE=��A�(�S�����i�����`��E^��9+t[L�참(�!j��z{�nN(�H8�1m2�x��5���t��h��Ϯݢ^6��'��=�Y�1��W.��`n���Ϋ�3�S�դ:��AB7w��`�N>;������ErQQ0:F���-DS}6-$���*�]U6��J�Xv^��7�p�>�<�L��(�-��\㯟��� �=e�ڠLF$& 8�`(�v�h�~<#������hp��ѣ����B�2:lvHe��R)�Q9h��<&A�I�ZE�P&:x�I�U��Ć_����[�����ή���rwХ���(�h���݃=)q�U���ve��]a���t�|{N���7ߒL4�m B(A�JĆ/�6�'@���Pʇ�ݺ.`���l�^�	mlޠ���"�>��zT�^PZɟ-��0�J5�c��2}���=Zd`���H����v�Hi�8#�/7w����kt��JP������k2ȍet�V�T�T�{	y���F2VQ���]O������`�*�,��ʠ��6ȌJ=6حLˏ��F�PzR����K�0C)#!Nj{
5�%-� ��}��f���u(���za���}>ϩ��F�J��Juv���^���� ��U��샽5��7�n���m�iw�C��?ω��A�=��h׉���|��dL�/�N_����ߥ�j��"�1�%��1��>\�i���
��QXpgf�����V��k�Ʃ�X�|냢����ȹ>̆��㡎_��~��n��'�)�՗����R��;�=��3�����
����i	,�tm*��j���>|�g�̙sғ ��=����%�� �e��d"HP�JC�?xľu�4��j$�
���l��P�>�����*J�L�$褟_4v�������:S`�,�(�ǡ��{��ʊ,*�����S�~ �" �l���������I��R�!���ѐ
�s�M�K#�9К�^�J�&`�bC���-�;tmҥ��$�`���R�ҙK�7��/�zT����������fRy�i�=�H�!9���aV��'7��:�$`��F��$=X?���^������y*��޵�߾z��}��T�+VHq�V�	��,r,m�|�`�@ہ�ڛEg}߷�5j3&��>zl��j)�N3׻cʌ��3���嚏���\���F#J�<�3��=��3��$���?��	�P!lq�%HV��
RK�e��ܷ��L�d���K�l��f!p����d��DA��W�hR��@��¥�D���g42���Mze�=)���������R�/�Z(�����Xk��򲥬���:A���O�y��{��5��)'=�y��!�<��2Ѩ�5ެ|�<(�\�}A6 ��Rɘx�g��3�,a ��������m�tccu}�*��@�3�N.�a��o�w�}��y�����>�|��D˹�frKi�*m8X5U��S�t|v�%�x �8�]��.m��ی�k�B���_cP������V�� VpݍG��rD"��]�r@ ���m�ܔ��-S�Gу�T�^ �{�(Mhsr۝=�����S
��ZD�{;���_��8���+ԚkА+�_A�p'�0Pv�B�	�4[��`G}U�S�)/��knu!�䣌���u�q���>�0��w}i�?u����hY0�A������䐝1�������ȶ!���F � ��Ͼ�}��{��C(`]��(k�۪�e~��c�Vk�$F�K	�XT� t��_��.D7x?��Q�);r=A�Ʉ������ʊh�:ء��ۿ��^y��S�����o��O��w/�E^;�pD�kg�ި�h�S#\{�9gDB��c�b�`6�[:�牨�����?ocW2�� Z�H2+%A�vr�~�����:�ǿL���?����Z^c�Z���x	��G��#mAԌ���L������1t:r��m\n_>�;�����#2;�O�#��g��(�����|<���s�ˣ��**��_Jv���qR8������E���j�
��<�2"�!J�"�E�*i�h����<�CV�׾_�� ���$��^O�Q�4"fMj�U������5�MZXX��x8��/�=�T���gټ-sEN�P���2�V���]f��c<�;��Kh��K������D�^^��˅�{�� ��Dk�^8���g8t��Zs��\�����u��%#�|��lli�8�����=y�,��[t��tk{K����cO0�r�d����Ω��_�����togs#��\�ya�0A��B쇖�#��=R�^����e�/1�B��������w_l6v�;�g;Ϭ�yig�ҟ�tXh��TT�խ{���	����O�}��De�P�ä����)��NQ|����24�o�O�����3���F֥�0��T�ѡ����P���<�D

��G��3���7��c�:��(�	I�8C�o��c�ݡ��<;�!%d�S���|V�V*�@�h���GwMŌQſ 2�4B!w1��*Uu�D)P��1o4|��GHHXx5*t�Ҫ
�EYhb�1UF)����T{���N���3�K��{С�x(��h~����'o�3�OM�^>�~ҧ��1��X�����aOE�NJn�e,H�*��jP��Njo4C�e7B������� ,����.����d���m��nZ�LE��8C�]���3Mu����@��sYc�ir6�yJ�L�|3����6O�Thx��S0Ґ(� ehz��d���� }mKG�ϟq��r�O>�	��<�)�|��}W6��L���դ�Y�a<�	�e6��_(s�M��3��;�on�!��ѹSk�������"-1 ��X�{`s���uR�)U��F������-Xd7D��=eM���H#���T"
"��3�a���G����M�o����A�1���T���	�'��d�\� �X'�D�����R���^ܧ�a�n������2�x 0!�Zo���+����7PѩYO%T��/�PX�ch>���V�~}�E,@~�Ԝ���47h-��j�n�u:��F��O�~��;{�	t̟	��`B��C)�E�*"�~n3�(M����(_�����gP��s�?�� ��<~`���C�)�Ҥ>�b��y*���'/</e�Y�~O�"�Ts�ii(�M��p��#���[#)���?,I}�_�
rߛAl��CuWf����9t������+t�Q������`��AZ�`P�����2��")�O�i�a���e���n�L*�&�b&Y�5�+m�F+��]8AK������p��Xţ�g�Q��wh����8/�����mz�xp�-��'N�
0<�ߣn�?OI���-U6 �
���c�O��a.\�#q�2��7����f�ΰ��ܲ��_�)�%��jx��OgVV�1�
Ǡ�`w{�����z�������u��c
Q��ѣ(��5eI>�~��?N*��nߦ�a��#�?�*X�+Y�}~�ԕ ,�$�;jK���f������|�#T�y�1�2���siȦv�����F���\X{����7��zB���1�K�W�yc���{E�\Tx�T��g�j=�Ð��&p���r�ߧ�Iw��~��~���8�$���>x�m�,`�{)�|3�W굹�I�?�^�l��~M/Ĕ��y�1�:<�qH릘a��֠�n[�����d ��ʎU8���"C��6$�&�)"�os���h3�ɧ��o���~���%y���Qݓ+���D%t�B�d&ƶr�"����p�!n�������Gt:hѤ����`�nm�b�u@I�":�06֞�k�8�@bPrIJ]�_��?A2�Ν��<��6;�lЩ7��n��E�s"[b�פ�ݛ�&3�8P(=`v �h�z�'�G0��T�C�g��(4Nk\��
��"��l`��H�����0Д��G�Xf�IĆ��ɒ�f2����
��/|����Ґ72Ox>�h4�I�kkkt�w�@/q2R��o��[����@���D�Kc��j�.=u��������Vi�B"����f�hr����k�N�e���؆BE�u�rA�2�\~�s�����n�U���'i�5O�����?���èΟ'r^=��ٽ��kV !�=m@
%ܰ1�����c�Ƞ0�v&t[�FAU2i1�mg<��7�9�i!j�|U�\<Sϫ���S� �VH��@R�-9��P�����6��y��9j!���0vD��%��Wg�b>l��h��a�V�۪�q�^	8�m�s¯��v����_��u�HIo����s�Q� �>y�X� ������SQ���5�(��Q����2��WhT�S�џh����Y0h���_���868ݭ<���=��͡���a�����@�-�j�c��>����;�u�ӎ�|�ڟ�?������xИ�̻���=�_������F����IO�PB؁�������6ƘKo]^�O,�ȗ�đ��<�TQxj{��EZ�_�8N�o!D�m�����u�x����Djh���4c�lOQ:���@�N�K��$Cc����H�y*��&ϲyO���4f{:A-b[���g��ż��R�I�d?W=�i%ǡ�u�WYzdЭ�� c#���1RH�Re#G%O�����-�c�d�{@f1��v&}���R?�m�d\Q��L�����z$��9�Odl5�M�i��0�;g�=r�*����:��Š2
�ISe�&��\�R$9>L���Q�
oF~��[��?�>��eݱ���;3����/��k��Rd1��AwQ�YP�^����y9�7Kx��EM�u|#|?c{/-�����C9��̻@$���2��K�Ko��^h��L�{5���̂UoJ;��#KgF i���8�Q�j�T�D�]�(�c�ݐ�^���D;�Z���@u�I6�B3�(�� ���sBt!�*�+%���Z'OE�M�u{"�ު�)��1�ј�1[�M��:d�pR��F ��TJ�
xΔ�Z�Hl��Ly(=��B���L��"�~L�΀���-w���驾��vI3�o�I!�8�`E	*��-a�Lm&���r�N�x82 qya2H5�@G���x���'r
Y����2|O	_ $�L��������i��u����j6��ի���#��`���H���@�F���-�4)�q���B��z7��4�=���1��B�jʺ;�4��E�-4������D�^�#�%����FI�$_ xP~X�2�KE�P���䪘���� V` ��)��߾}��������)]U.$Ayݒs�(K�T�đx�^�׈��QFO���*;}qL0���l�F7�>��~�}�NoL-�W�c� A"��`��c��(��u ��y_�hVШV�l�	�Ԓ��YX�����h~~^��d;:S]��$G�1��wi��9q�P��[Gk[��D�����
?�������H�}��O�K�$i"�췸�Z{����
�&!�{c��|�4A��w�Q�������-��;��ޭ�,ʹ�(���OI�\�������I1������SLz�3��c��鿎!�Q]��[Mf����crw��]Ws��;��u���� ��`c,���J{bm��E:}Ձ�YJO��})
�>9-7$w���@J���$��Pq��K^�S"���d��M��T�md�]����f2$$&_�&9Kn�@ơ*T*��k.���/�Ӆ��LX�}yh�Ю`���顆Fvnb���kT��Ku�j��v~�dTZ$ �Sh )(0\��*�J�'��AVOl�C�ޅ�9��Y\\��`H����b��lV��hmmU^�y�Z5��;�&ݷѫ���Y��B4n}�����c}�"N���G�Y/��)�S�p�<F �Dp9
���.���t��e��Q*�#�Qci��s2Pxt�%X�(|�>s��k�����֮�x����Sz$�f�{bx~
��ux`�[]�/%	���B��"{H�&�Ұs�M��_;yq��\Z�Ϙ��ϯ��͋���k�=��8���gH�5j_N����z��͂�C@��`�Y��:f�Z��G��ۖK��#'�W̷8�����GQ�s8K<��씘�ge���>lD6�Hh�'	%����� ����!h��J(�)�d���f���Л�f&Xf�?���St��pz���s=�# �)c�l�#������=���1N%Uk���>̴�*��hw����_�;���V��~��|�qz|8��k�Pe��|"��FB��KN)��L��d�Slj���q*�p�A�	M���ט&1�1��8cK�I/�� "ew�~����j��L�OS�ɳ��/h�jSOE��Ϧ��6E,%��(�q�Ő���RѠ�'���	p"m� ���Y��2�~!G��*���z���/6)��H�����}~|��X�+"�QDs���"��O�A	���p%�2y
�N�yAz��V��nXg S���ߢ4T�%a�XA#3V�O�u���S���r�9p��<\�7�D���P�󴯸� � n"�o�jBR�Bd���8$�e�������jcB}��=��}�5>G��0�dvC,�Ik2,(�n7꒹�,4i�5O��$�ّ
j �]�CW��|����%�2���y	����RiC� 9;mQ�Nv���&���g����"2���{�u�+�g>���	%HOc���P��w�}@<$jV$�a09��LgN����4�h�+e2�'��.�l�Z����A�b�&�*m��4��AL�ф��v=�����,�����

KX^8p�aw�JR���`��j	�ۧ5�SW���dd�N3�(�3��s�\ڋd�.�c�i�������^oj3���ƝԷ�9�\�X>8�����,�1���*6I��s�(���B�\U��һj��������d>�Gle����p�Ǔ`�����<	d�f.�q0
�HW�p-R���ԉ��{S�)�h��	B��ߴ��1O�gml"VI����Jp.�ה,Ѧd�֭�V/I߮��C��F{�A�dv�Ā{b�4�T��{�qU��7������� V���	�a�y���*2fƕ�c<\�uQ���)3j�T;xE��\�S�YL�.�-
F!�� ��*�w���RT��J���8� ���F��;@j6�u$8�T���h�&]i~�k|�K�`�Ü��;2�N(����|�h�n9�S��cVj�t%+�:���;J\k��Hp$#v`����h�<�h�X�'���w�R�%���W�BE(�gI�,���i���9��4`G	^I(WR- ,�?���mS�8Q<�*�י�[g���#|�]\�n��f��'�JB�7(��i4�9�w��WNz$+sWͳ���4��/��������k�0z~%0���qRN�s�[��<�C�'��~JU?k�)���l�X"��2R)�:���ݐ/芁�$W�AL_����D�=)�@���k�re�cj�����^���::6f_�	��f�AP���DK7�C�-�B�)wF��o�����*��ۑ,J�V�m����6����maż3��Ng��D.<�4-��P�Z'O�O�1[�G��
q�Q��8&$���S�I](!�Ȏ�|yZH�j%hHh�%�ZX7��h��Ŋ�n�e��m��{p ���N�d]<)��hn��*�VMQ���%H��.�C���,ĩT[�!a6�T+i��k �/d�p-��@� �0&;{�3@�#���C����[)IM���[=q��OH�����	B� UD���<SރD��SA&8bك��d@s�E`��1N�
I�F�F�"hJ"r
�*����[�oǠP�#��dP�V���"Pك�F:PB�I�f R+�S 皐�@S 9�����oekxn��a����?��`�E�ByR)�u��"�p�x�<�'4�4�2�NOXk!0Po,6i�ݢ�.����tu�&�q�]ڎ�R�ٓ�E�M�җ�5�{K��J�RE���N8㾖�W��mlmʜ�v4?7/��U/��8��\���H�5#Hg|��/R/S3�M[��<� 7��C~U�]`����^�<w�qf��Va��#�����"���ǜj5�n���I�Pu��1�����5K�R����Cn�ʦ�� ����<���4�G�n��(�d�I���@�� ��� ��qFD~�Z}����Xn5!�	M�MP�6X�r!p¥���/�vUsP�z��C�k�-h,��b�E&$?^���J����C��4���]()���4�j�@��X@���OT��M���;��e��u��%�º�;!�^틖*
�/�>�?�jW��U1ڳ�n��T9�$�� z�3-+�_	���K˷I��g���4-+��W綱�bZ���b��퇎�DN;�0FL.rt���D֖�Y2�7��0�A�b\���$h��{���"��F`3|F��TE�s��:H@R&6���+�D��������"�j�Jʕ��
d=m����C{l#���=4�R릠*c����lK��.H�4�dn���r��U�ܸ%�Gz��ق�"�UEj�}�jy�c��� l�g	��ԏ���VI8}a���|�M���r��~G�Ň�z��v!�i����y����^h�~���3T����N���>�O��D�.!c���|z4\����z��<��!쐙>0��p:#�aa��"�,֛���v���^X1qaa�i��о����e�M�T�l��gk<�f\���P�����q
���4k���?L�A�G�!�-u��3�Ү9@� !H:�GldM��dKؾ  /��`�SId�H�zz��rT�2ǌ�И2*� �lO�g��ی\n�u�h�FVE��aJ=-僘�j�E��1Q�R{��x�Y�������v�mZYZ�?��W�D���a�eɎ���@�l1;�c����� �{�������	����D�LV�N������!D䊯�P6(Hs�e0`�1�k1`ˤ���Q��a�k�J�H(�+e��i��08g�X�N6��07��Yx��ΰ���'��))����x��~�z�Ղc˶Rm�T���"^�`��s�Tg�L�����S��j�`�#2(�ٺ�AKL@�����~@Kԑ]� zǀ���-�1�q���� ���f�x��L��:]��Qw��Q���M!���#��v@O,-���e�E�|+�d���wD�3��F3��e��
��Q�y���Ĩ��<2f��kU�t��)D����FQc��$V>q63j3X;�v�"ދ 1�:�tiai�6���	�g�$���ȵ���k�V󩆀�y��%먄ȹ8B���u�7��8����=y�:o]�3k'iqq��ģ��Z��5���5�h����$�?���d�%C�7�H�& f����#��{�5�l؉���=��z�/�/(�ZZ]�^rF $����W����]__��'VEK���?S�R�R�>bP2��=�M��<�3����I
��g�l�~���7��>�v�����
o%����
J @s�_(?u�nu&�ƴ��G�QG�;'����jĩ
�^�҅3�h�ђ �{�oR�V @^�?�,�N �����"U0����V�J -蹑�B�;����8U��F>?U	d@��}�,���:�m�e&�`�|K~�4tQ�.�k����'��-.�M�ņ��p�g bM�bW��P��K񜅳�z|=�6��8��j(E\#�Z8Fn���g�C����O�OQ�l0�-z` h����ɠ�
l����F�}NeI�ܻ��8���E��^��6�h����иR�P�C&��H��lv���f�զJp/�^:ٓð��8�n���I�+NV���V�xʃ�*�s����Wg3�����T9���"7��x'�|���J�]��!�<�At�i���dˍ+޸�q��'��(��-�-�H;�x;�u� J]�V�`4� #X0�IUX�P�X�A���6�y<���.���+�e۔Đ�ߟf�&l���B��5BRER����̎���q�y3�/�vĦ�|�øYo��Q�J2%繾y�^����+Wh7P6i\W1�e�����^���/God��9����F��.R6J�ΰ����$�i!��ɤB��ቱ�1�YI2�<�b��p"Hl
[�?Nf�QN�e��K������c��LR�6���2:��3@�8i�c��%�e�	�0P�aIel2�!>�p��a��)��^������e�\��7.;y��(�����C���_^�e���+�)"-{�a b�F��Q&��JЗK��'4� G�SY[!z�������iݽ���E� �ޯqߋ���Q�>!cK�Ht�Ƽ��|������:}���T�Z�.�zF�|���'�=�ꤠ&;J����9���Ӵ�b�Piѻ�x��ř?5�,F��#�4��Q��z]U6��?sokYv]��ۼ��������Ȗ�F�@J.AeɆ]0j�aO����0��@<��.�
U�iY"Y�L�I2���������޻������dR`�J�?D�������k�M�ݥ�7d=[��.��M�F:P,�&ݐ ҃�R���)�7},�>ܕ�����v�e։��KWnJ9_���Ci�ٹ�t�E�MzZa|��I|��^��{ 't %�4q�:P��Ő�'��:m�m�-4�v A�"�~�ͽ�pG��z_�O^�U'�qC�������k��/���ɷ���9ޗ�jU��������O���[?~(7pM%8��AS�uyi	������b^�z��� ,�2����(0�r9�}�h��̮��m��l�������o����X���5�,#��Wo���Π�闗����/K��� k$u��Q;{
�dZ�8{��������3>Ul#+�������^�vC���P�Z��/Oe2��'d��?t���\]��oܖb��~Bi4�༰?cO~��H�s,�r^�/o)�s:��~[�4�i_�T� <c�ثc�B8�����$'����օ���5�q||,��},�>�: l_�_�)��U��e�8%�~W�ځf�S�{F�6�Y#[O�ھ�Z3��n}�Y��9�paS�߸��Y�2�=E�5C�	��{��:J��Z�,��P[�tܙ|�<�\%��5�1����k��̀~�\V�dҭ������ӎ�-����ܑR��7|��r\c2�i���{rz*��<�{��o��dQ`�k3h8���?�/���5y��D����[ q&3�T*��^��բ<�{*��/~��{�R�gs�gn_���Z���UG�zk�V�ͭZ;��w�}1�k�R�egxn`�mo�o�X��Ѿ�O�Vҥ��oS35��z��R�)c|<-��s s�T0n�uT�m��ڎ$�J�J3��D>W�~�k0�@I{=�y&X�����ۇ�2uؠ��Duc��?�~�g�l��J<�V2i}��!��Xj1{Ӿ��a��^�8ðQڧ��=���n���uK�i�.�ɾk��1�8���Q71m�4ce5��1�W�{��|�(璽����Dp��󡍊&�93Y*Ƿ�^�ۏ�פG��
�C�^�L[�)f��5��r>�k�v�ڔ�}֞�i�(�$Z��:G2� A�҉OÔGa��c��Ǵ@J��N�F}���S���R�Q�s�`?����+奲f�	�c]�fV1oE�y�#F{G�M�-��鰇}�=�n���=[�'�X���B)��5���0'��^lam2ؗl=����(zc!�	Z��t�o���Z��}�*[gŵ�zp �l|0��wpO�����~��k�X����Kz9�w��	j�1��c��_��T��`b�5۞]a�&��Ѥ���O��]z�o3���1Q@Ȟ�E�)��C��al�?ӿ/2=J%0\�v^6v�9�~��E?�P�3Ǚ�'a�b������H���W[ ���F]s���G
B��s�j�{-�}F
������-�����o�!���N	L$���$f�T$%4��)4>��0�J��X���1LZ� 4�-p$�bN����޽k�i~БEV�KaJ��3���
l����v��������nݕ�ߒ��e	��0��
�c���#ك���a�á�/�]�s�ݻo���/������ RH{� �G��/��S�˩;E���ޔ;׮�����t�d����"Ɓ�pM]�d:���fvd� �j6K!����Jyb]�A8�f����L{����_������������Y���=8΁���ky��{�CMi�_��k�_�'��<|pO���ɠ'Y�&��: �ش����&
�q�T�p���P��J��R�Ѹ'������u,# �)*T��\0�7ַ��^~S�Ww��?�N�%/l��/�E��ӽ=� ,�u�<��*�v:-���$b�a�k��CNH��K (VΫ�B��X#�4e]���f�!�~�ؼܽsG� !n�ږ���d�|�Ͽ%�=��(�]0C;�Lt_� ń�(R����ibVJEG�}���\�7��T����"�K?e|ߕK�՗^���X{m y6i�Z���r�}/�Y�`H5א���Wu�9�����7+Y[_��������q.�wo����-g�|�N���AP����m��_�����'��@ּX�j�HWL)��6���\Z��\/IԟJ�CZ����;�Hx��~5M�c�s5^�p�9V��N��V* ?Y�`�����F8Ǧ���h���XU��r6����8�^��v�k�T@��sǫ���,r�ꧤ�F��#�T]���T��;E����Y"��D�=��xۑx�L�oL" `�(�1���s�65n\����4�2I�k�԰��*��#�{?�d��
��	��i+��JvU�?�x��=:��8�Cyt�'cfómy�s{��ݎ)k �~���
�K�vEBI:#W�>ّ�?�H�ZǢ%&N��8SZ�ki��Ķ���<F�F��4�5RΕ����W��W�UG����1�=�奚�a��i0ь�x<R�(��zU�\{U�������X0t}�Jj��}s.���ϐ��h��B>#ˍ���p�6Z�p�C���4_�t-�c�h�̵9���Om�m<_�{�&|V�&��Tm�U�Dgk�d]�q�2�!�5L\�{R5gfm��M�᠙d{ƪ�b���Gs>�VM��\��hf�Gi����cX$���GN�<&e��"���a2�nbEsO;ٱ�!�ha�Y��[�n� ������h%62�WNi��Ϧ�mb9�`��r�Ϫ�'=^ޞ���]y��'�{�fo�=��q�f8��64PH�%��^�y�L�M_�Kg8�rڮ���8�1KK#7��fR�����p,c�4h��Y�8�����;���n��[��ͰZ����Ҟ��9�pV�&#��|؜�<0,h�
ii�C����ag9���]SҢׄ�*�g{ѳ�M#&��Q�F�K�"���Ήa_2Q{,���t�1l4>�!L'��^Lb��j�W�ɳ�;u¬�_�v���q��f��F���v�嘟����<`�-��V�v>;��>�o�2�7)OL�G�uW�(�^Dy�����,C;i�'%�<�=���4�x��S�{���,h��/�3�/j?��klA:)%NdT�T腍�U�SC~��4"��TL'aݓcC�5VJ��d���2�1���T��G�+���LD���R��v�J�����ʬ����R#3�iQ�X�E��Yܻk9�4n�k�f�(<�-�'V�a��/���>U��Wn�"�rAj.�]<��>�w�ޗ�p9�zA>�ɿ�������㙑���}(��<�G�;*�L�*������/��G�Ȩ�Rz�t:�F�pU�5���tH����hD�6�L�%��PUGb^��m� Vc��A)�-5$G�0��pM6������q4'C��\�,P�',�ZWI�]f{	�[YnH봮Ժ`bye]n2{J1 Fq���Qe�Jf2y�]��)�	{�������U8;�;y��\�*�����
I�e��%<���b^�`#���FC6V����k�>9���)�2Ľ�i�za����#
g�t���T����n}�.�[B��{'~pi�'����J�.H5m�k  U�̹�? A��ё��2������6G�2I�bN5��5�|�Q9-�Z)U23��N���XgYRd�
 |��)�u8��|N*Nƣ�f���ʺ���u����֫_��[
Z����Z�/�ve�\�+.��'Xh��pj�r�D��Ԣq�(�hA��<����;�#������}����1��"�5P�qb���i 8+�//KߓO&�8�q���Ι�Ӏe�cӆe
�ر�X�q�1 �* ��v��\ґY?��[����*��"Sb�����Spb 3R���1�$�9)��^�	�!�S�Z�j��E���@k̮\�.7����{p������Y`��lf��2kN`So��u�q_�?}(o��2teM�2�1������c�O��E����6VNڝ���'Z�mQ�H������C9���+S`�X�θWZ�0��Q�S~q�ܼz{��q�	\[���:�`ѵ�Ñ��j͍c�|J��L�B�F�5���)Hu�� �B��\��Gc�u�L!!KY��(ϥ���7�b�_�. ����kqF�'�g�����ϴ�wn�|�ͽi�|�+_�~�������-��Ǐ���4{�=�9b[�
��x<Q`�df��F�����k�-2n�g�9����]ٌ�>��Nl���`0�g����e��^�s�����bI2A"E���WT���1N6a�3=sݴ|�2��4�a]̵�B/p�YW�[����L*gd`�cj�����z���
��L�LUEj����?v����uL}f�i{�j�M�( ��̖13���Y�X�ee�$je�(�>�q-�F�����y%��X?8���N�~�e7�Q@��<�F`���=�o�u�Ao E������Y�|>�}[�m�ͨM��
�،�&O=G����<dF0Ě�X:��ާ�^?�mP�f�m��w�������`1���QJt���"k���,53~�i��:�N���r���1h�|�{�a~Ü�v����3�Β�@L�:oQ�h�N�d�$�r�n�؏��'�P,��t� ,�'3��9Y%�Y�o�Is�ϕ{��؆R�r�8������t��L¾K&���d#� �)�M@D,�.��K���k)��������ꮻ��i!����Y~���ɦ~����q�k�S,G�Ӕ����͍���&:I*�k+��Ϡ!%�g؜ґb�(%�w�'6���̳��6�j��X`�N�ԉ���z~�iɄ�|�<7�)��7=,�|a�s��g��|,��s���	ǎ�X�:i�x��3/�4��V�Әt�F�M�2֦ϡ6U�,�u��`L��̰��S.^0W�GUV�Ma/#�3:�C��g
I�2LΏG� ��:_�n������zQm�~c[��joC��~"��G�~�z2��M���i�`�y��5�<F�������~��|�K�� ��?C�a�@�Á�t|>�'S81�%g�z�vA��Q+3��5SiV�k/� �f.���Id�7*L�n_�@x��@2�)
X�
Eg �Y�vus]i\���e.;x���b��)���p���1l�S��'e����h6��yd(�ٞO�����X'���Ky�U��_�r]V0��8H\6�Ȫ#��׉*č�c)T�p�8� �p�H��z�
љ������+w�Y������q��)���T)~���։�����˥�W��ɮ���X���6�C��+�ƪ=֌ 3äinnm`nFRkT�`����PU�f���
ʐW��Nb賢v�Uq
�����-Uʸ��d �G��p$%�}�>Kp ��򵬫����謒j�b�O:r [6������t�@�#�V[3[�Ӗ\�zI֖W�s@�hN�J5��D[�+ѧ�g4?:Y����-��,7�T\��J�*���,�x*�� cC2Y�ˀ��(�lA�Qd��N�P�Zh�O7�+�ε闉�C��g-�t�ƃv �jM� �i߳4s`�kb�`g���QaVl0Jc}E��Ui-Ջ�1QNx2{�����tGFH�^Y]�+׮i���]k�p�%��ƷRj�f�J�G�n�@������ԗ+X�� #��;�m a�td������Zjh���Y��J���C��	�NN֪���XU:^��23�'��c֩Q��:��~��:�,�}yyM��yUf~����m�\Rp���+�>�/{�C��ڃ��1"V�ZmQ��XFG�}��\S,��JoPПHPX
���i@0P�Q󕗵�m�T���d��D�ws�Eiw|o�_1�2<��|�IQ���s��ӵ�'� 0��B����o�Z��郖\�V�wR�7�t��P���R�~�b�2��b�.om��뎂�	�3��`,�X_4��e.;�z%T�����N���Q<��A[�]i���#<�9�d�ry��\��-�rY��<�ӓm Ζd������Θ�*��|�0�<�(�^�ae(����c�:��z1����E����b�b��������R����}��%�Z��ϕ,SJ�3�6c�SC�eX�b~BۛU[.96���^r�ό�a������IC�<�)ÇYW-;um@�¸��	3CgLl 9W0��jVi��d�K�j���l���љ~�1���[�Lh;�4[��G
��5ʩ�{� zSp� ��8VNeژ�9ӝXd?�X�4�3 W�\��槊���b��ɨ3�E�[K�`e��u�Qa _Ÿ<��@�؂?:���ͪ���g�8&o.4��Ɨ,���u��Ga�w�_�/�t�=����6����_�&����e����h�T�	s��	�`>�j�S��t�ʉ�$�{\�<�t�Q����zI^�,���/U�21&�%�l���jŴ�e|�r��e��l�ȓEz*:[��$M9��&j� %�)@p�2^61Z�'F�<s�l!�{�Y��*-&Tu��u8)�?�>����b|�4j�,ba�xipɂ�4[�cvԥ@�9�����A:_`���U�s����.��ߓ~�U?6e�6� 1�zں?�<��w��[���\E.���hab�mi��3��`}�ZQ P<S��L�J���} �܉%��1I3֝eLM����������'�ݳ~�E�Fժ�%i$�N8i]xowґ�æ�glM*u�la5��F�k-���Is6�C�TQt���i��'�n��e �J�.>��j<�<_[X�L��� �M#��C��@���~Kܯ{�G�Tՠ�:�1��M�@֪��=�j��ܑN�-Ov��gB,Ei�����<mvNuS���T9���ɱ�2$U��4	C�AJ�����Q�G�� ���z�q��T+uͮ�B78�Qʔ��4fX73��9cF���O{�<��9�|}c�ڱ�,�������QX���i��Q�Y�lU���@#����:��\���)��VG���L��r'_�
UHGkD$G�H����}���!��P:!k*�FK��R>I�S�o��L��$�2�ϕ��h��V�ylT'f��-_���ܾ%_z�-8}�`���c	s�3� �"l_�o"Fd@f��c�܎�#Y��u���T�9@���1`Ć��H웧"2��Z�BZ�c)��d�gFc�����i��A�����Zэ�-Te}�:|W��Hm�9\D��:k�߷��z�(�pLO��f���`��3~ֶR1��[/�"i����A�-} ��~K>=x"��&�~]N��x�Ǧ-J��q|C��s�E�:F�.���T�y���}S�b4w1.c��r�k�y03tQ��B�)�;k���ϰ���t��?�sBF�x��	f'p^��T�
�j�36۞L�JG����x����<�e{}S.l^��v[�]�f�B�$҆0�+Ņ-b=s�V20 �9�e|��׽�s>_���צ3�ɩk�0;��*��('�9ɞ1��2�-���p"˵���F	�p���S�ZI��4�"��U���]ތ���Q�4���^���%�Ϙ��S�Ba��
y�;��r��\�xQFԓ�0�����ּ2HůT*R��������wdzp��Q%�*f��J��W�:��ь�{�1����~o,��\���E����� �݉L�i�+�'�a��:NLoֶpV��M�ԝ�Nn�v9ۜ�+�U �H>~��+)�t��n����[/ܕ�`(���c�>.-/�"��%#´�<�>�E��Ն��獪6��5�Y����J��]Vz+���6��`{�:bbut��E_9�9*ag1?����?�������z�uJLۘ>o)e,�����Yi�0�~�RJ�9��"� -(�b����!p�	'�'��,�9��,vXƜi�a�M��Lz/ι�c�Q��!@�ʹNj�����|@?�g͇`�:kf!�#}��$"T�-6�]�[󘤊��4���&�y��.�溦6U[Qh�Z+��%3�=��%����'�~8��V����6� �=��~]��[���k�?�q?�=_��48V6����}#��"JR��4'_��#���8q�2�i�M� \#s�4���[�|�򎭲Ws
"�"#�{��E�1��n66�H�e�^QA9Cĝq
xC?HW#d.<콦��8��T`�K��z+�6#�!Z��G�L�D����v������.��]�h-U@��s�E/_L6�O禶Y�-@�z�8��Ϧ���y5���T��zG�	�$f^���Mk�R�m@�ysJO��,� ��QGl��k$�;�L���M;![���'6�����j����4�d3$G��Yw*Z��C�����5�U��	x��P�J3�g�>[{��S�GDH琇✅�\�yWk�(�X����z��ic���}��+#Ja�}� ns��F 0Ӻ2#;�F����F��y8$ix�p��مS��%��Lcm+�,���l��O����5���H��' �2��Q&�}�/�~Q ��qO���;�{�iv��:���y���_R=8���!k��|S�*|�Z�:z�D�f���N�S�38'�U�J�2���}`�)j�i� �
nW{�� ���I��T;��P;/���t��%un�x^U
]S�������Z=�.)K}|�t>� ̒�&r��Y��5C���h����~���P� ��/mi�ǆ�����-/Uj��D�3y�M61A-�N�G���=�UǓ��j�j��b�:?�Ȇ������\Xݒ�$�K.��/ܑV��sLEM��ď�L��WK2����yN�OO���j+�nmΎQ -�<H?�`�s��xӌ�����3C�J��i���'EpLe��ey�s�� d09�Zd;� �4�R��XY�@&���TY[�:L�I8�̾�LV�H�ab�:�gaO1�n�]�ݑÃC��1LJ��Lڜ-W0u ��ɉ��@�S}���O���x����BS��#�6�u;�mh�&������y�����xc���"��>���% �ʁ2�A��� ���ٓ�|�����I����Yw�M�~�� �Ś�r�Ӷ�c�}��l�xS�S��t�١ �x�����P�"6�g-_4�Txh��zX�Y��I6����ْ��P~jJ����涼p����ڗ��Ӑ� 8�%͊l�=���g��FD+�  |pe�"�#�,QUdүg���Y|�62g�:��F,I�V���U���4���)bm�>�f�i/�`V��Ĝ?��K��=R�k�e�y `^�V0vYic=Up�'G��fˀW_}UV6����G�qry���
��JLO�LN��s0t-�n]�Vw���r��-I�����R��I�(���� X�&��5/98�y�E	X����a�,�x�׊yVW�Ĩt�51S����ėl�ԯ��8,-��h ��=�bqC��9	 �w�2�g8"��Şfc]+aT]��y�,U�ƥ���,] �{{�r�<2=i��f�U��1�i�f�h�غg�P��._���N�T~�w(�����V��P6�[�:��9��1��@�@ǜӋ���Fҍ���ȋ���3��7��3�Hi�Z�Z�y����f>��~grF�L�Es]� �������O��<�b>s��o�A��>Ty6T��=y���_�dA+&:�|3��N��1��)�p�f�MQbC���Y��M��i$���iL�!u4�:�w�(��m�ޮm}��}!�V�2����|~~SnD�9�C��5d��:ʜ]!�y.0J='~�%�Jo��Ա|��Hr qE����ihM�X�
z�B�`(*p# ���O4�9���v��m0���\i/�~f
���R����Ӥ`��6�3
h*T�����|�%�F����Aa_����^�N��06Fn#�:ws������׏�@;i�j&S��6&m����L��պ��X@���~o
�R��Ă¹��D�T�qU��_����oӠ���%f�k#���j}��$�,]����5t�H������������40�@��(� �*pP87�6{��6`�d��ɟ�u�ģ������y�ݳ��-ط�_��f"΂�H��YoJM�cf�f9ƉfM�U�b� �/�Y4g&��-#�e-׀S�s��'fM�4��͚M ��R��+��g݆�{FN��p�Ĩ�g�V/�̳�=�=,�`s� &��P�  Lf���!yg&-o�t):��~�RNǣ�7���<��p0߸��|��D��S�Σ@#c�}�ZG��4_��8��� -)X�E�seʶ{���ཱ?�ܑ&��~�3��&���x������c\�9S�1MfZ�8f��Y �h{:��#^*V �*��/� [R�T!. �P�E������5x�-����Cͦ�&�TH�t�3T=Nth2�Gщ,��֦����S���
�;�Qw��'��*D16�NuXN�Z���q�Eqj%y�S��pmE��l��qI�i�t(F���+�"��� ����1��=��%�;�>�N��,Ù�ӜS�[��f�)�>;E,4kݖ�X/�qf��6'צ Isry��$O�0��`�$�JUi��� '��
�]RMqO�i�g'��ɵv�V7�
m>M��\�9�a��~�,Syx�ǥ��*�k��(�
����Q� ����1�lU�F-�tǹD�/�X{ V�zE�kd�p��fP��*��k.s�2��L�O�1#�`OUJ5)f�7��k�q6_�^gs��2�u�H���>DGAFb�Ƒ��K�����i's ���V&�ܫ�pu��1�qzԖR� � 
���#�ȓG�a� ��U(��f�a���U9n�T�mH#$%�e�rY�R�n_���
�<�<���m�c�R1�����<k�e��e]�i^�(7�⹡��34�ن,@N�ٔ�ISpqcNzi,�vG[菆}���bͦ��Q�4����j}j��@ETL{ �hǸ�]��1�3��4��<� ��f�Q�5�,�%15�eZ��h��WFA  5S��}���r�;����v&W��+7��vA:�M�R�K�Sc�/�c�`�E���K`��k�s����s�kq��o��3=k���BN�j�g�猪)�C��oR1gY�1/����k0[��Ҧ���LU��l� 
:)2���VJ�0f�(����/H��"�&#�wx(���N���:7b}���O��gf��r��k�4d OOZ�pʸX�1;Hlcz�d�R����>O�K���i�p�� �ql/��9��YG���8g>������sNY����!��rV&s�l�?�b�&j��*�KO�m���g�#��K�g�R&SH�%�$�X0�%M���mB�4���M����M[�jĈ�����N[K�yp�䈳H�$���-{���������/�~�`�<�Y����ڃ2���I8�&38s���ܮ��B�us�`7@��z����ěm4��-�}'M�}��V-��<N���qm�#Rڌ�X\)O:����0�Μ[�t�1��@ZSg���:�z����ɐ)5�ܨ��尻��I$$p$m/���-�R:����8iݡ8@��HRbf���hչ��������=�1S���z�8�Թ�t;+�%6��<_:gr��۱�.52�����r�S�"����}�Y9�����c��#�2h�������:�v�L��������
�l;�
,]��`�s�X1q[g����Z�aaU�d͔O��E�O���X
 8��!�h4�T�,^�"��d�f�5��8��J_r̺K�ί.>����FfM1[�y�s�gTIњ�v0c8aS�/��R��e���,Pvk�QxF���
N�`4��Z���u�`/�²�q�X'A	z��������#i&��:����NxD�C�����G=����z�U���X:�c#����Ud�Ͳ�_������X[],�Y�`O.=<K���C�GH8�3����q�vó*kl��cD5�d"��R]�;w���˸?�LG�3�������i [�&[*j-��T�A�%����Dt�G���5���y8�\wAp 98��j��0J&,Jg>�M�M�,�L��'��p���T.i͙��P*`�XԌ6�7����yt�l�tK?cj5J�h�v����h -�ҍ˲�k)�%����7"�_@�� �b牶�5�B�1�%����L�X/8a���:��t�Ŀ��i.2����^g\���=�J.c�&Si�B��`�i�<��"�3M1�O��JP�/��;��KiA8+Bcj�MO8װ�icE=�65;-�WUU��+3o���?���:QUF?훩��4L���<S�F�Ԃ�lI hg�Xz^�x��-gJS5��f���33� 8<=����)=\Wf4��B�))hI֞�_����H�ÞL����H�©����H�e�T5�I�Z�L���\m,��8c6��M��>�D�ߟ|_VV���_���p����0�>%�`2�=ϔyC����uo �L{C�08^`��M���d�5m��_�/�f�(ۣj1{�{�	�3�1�7�$]+��_�g��G{y&�ĺ�m�2,b���@JX��](�f]�����nW۩��#�`0K�ژ��
���U��N�P� ����m�6¼Py�:C5E*�b��ݎ�G8b��6-goB�_1ͽ4��j�Ma�\`'��iWVW7d���|��\�J��X� �g�
=Q1���*l�D�k����4s���i�'�eB!��֚�%P��� ňL)E���p�G��>���4�}�5�=Ĭ7���)�x�u5���+!�v�Kkr����]���D>�ݗ��G���M�9-��o`���ꙮuLR���O�l�ɞ�I����3��XY#��Z����B�
�X�|�,a�M��8ag=�L���9��f_�,^kn�~�s泝�N֏���:w߾$g���c�R��u[�*�3V�_>����L��F.r����l����$*�dr���~�a�p�җ����r0��Y��M�ϸ��t�L���� ��$Q����k�X^�x*&�w�8==��'�(|;c���FTt���Y~��(:_餥@�M���s���{�pY~,�|�I�~���/��pe�������q��Ь�c���hn,���:�b6�9P�V�.�Dlt�l3��hi���pw�}��[���q��cC}:���jO��8gߵ�[tl����>��K3��~��6�9��g�?S�io��k��IVA[���߹6�C��57��S7��8b�X}EG7�(г��0.���l4�<}4���H�{&:�EtL���nZ�]�`�d͛�|�E�����_� A?5��Ɋ�=������*�e�����4az8Pݡ88�Y�0�T6��cvf8�F漉)[D�uZ����F���m}��}�U#���ZmDS�9���k�h>�*��ꨮ:�bǄ@,9ߐ���\N��Qw3΂�����[P�ˑ%�˅��p fHq&����_��p]f8h��� r���@��fG����Ɉ���*�����[��11i��154�VU􃆟M�' ���W����♬:ӚU�L�� )�щ� �/n_�f���Pc�̢�a'}�Y�H<�Z��aS�B^�]�*�v�����E���lT)6���$ P:��8��1�ŕڊ�JU&�P^�}G��<�!�؞�s��ؗ��p���p���)&Cy���u �, �؀5R��Y�n*��<�g��'*��Î���;ӧ˕5|���EY�/k{�	�=��al\Q�`����x(�vyiEVVפ�d�=���A�T~��;��ސz�,� �{Z��*� �jG�Q����j�����ޡ��0���0vc��ڟ(=��9�>�➌&�Y'���ّ:a��c[�C�_�Sz��Qa�4���) �;�T˜����"K�r�s�01���G���\O��h�<gH���~��T>�bjv� �Qlm�u�S#�5U)5��13B
C%9Wi�m��(�ܵA=��*�V.��|��la�� w������Y#����Lbz�� �60���y��U�����t �=0�ǘ����eF�ǱYv�,A��e1^���7�~W����{�G3�1�;��!�n\���/��~�T�2�q9f��C��
�^k�A8���h�B���9�v����7~���	��jh�j%���Z���	�l��C[���I��=+]�U&��{�bI���*�.0�@��o�Mc�8�1��0���{�qHB�5�s9��b�G����im���ΰ����3���;�(�������~A[\�,���斂O\�ԆS5���U�y�E�8v�'$�M����LRKrxВG�v�������2���}(�g�� n6�MD�9�{\�lq �X���GX��GH�'��܊d뺸�b2��;,���d9Ao<�DE�����#����������|$��Ao�k�%y �s�sr*�v�����t��ϋ���NN%7�R��t#J@H��5���o�}����'�eh�H�*�'F��/��?g�9}V���$N���I�:
��ңR������gg�Q�5z.A!6;��5q�85�3�EYЙ�{N&9�<ʙo�_���g[}�4��&o�H-��w�O�FFI�l�E�JǔXiY2}O�2��`�1}�Y�N�y���cՋ:��Mp8g`���u��P�6�|��Z�x����7o\�vo8�����|�۽=��Wf^R&�=����D��� ��SP���&gTER=H�����Iп3��+���pT��^�'�s�ϧ<�PM�v�4�N�"���=�.���F,W��m�ڋ�Z4��i��G:Qg�D(���MfN���4�f����&�45"7<xxLE^�]ͺ�����#{�.��6��&8��a"Y�!��f3��u�[����&#��������#3��{)5@��d�	���l3���"�����A���(��"��
��a6��>��?�,�G	V��4I��t��j��E��H;i%���!c<�a�@��/��K �Æd���8��.˖&t���p|S �`.��P��H��\��)�`(�a��c/�D�!3�>r~N�X��YVa��<�a��Lf�8��{F�8�^�Ū�Gw>P�¬����2���{ƳP���&�E�KG�Taf��Ԏ�k%���>K���;�lC�H;x�g���5�}]y�ԘFp˪��� �������d�8���/d���	�;5�Lƍz�B*YRd��G:'�QG���'�.̀��DG��'��#�������?�Hw2��L�D��a�{�-��3�~oO6�����$��D���U�4BZ�L�ج�HA;3|��_��/�R��$��� H��b*�d,WA*�����#��C`����T�+t�ֵ^G��q�b���eC�0f@ �H��n̗�2Jf�7�Jκ'{�\S��{����b���ax���XVJ �F�R�F�!c�p�53�Ah�Gb����J�Y\k�V�ְ#�zC0�
�ƒ�ץ������+�vO޼���{=8w}�Uk���Q���`�G1��(�^w$�+��=j�>�{�%m�;:��:���K�8 |���ڢ��I;e�4'��/D�� A+�V��!8ִ^�
��¥KRf���P3��LQ�]���!MѢn�5��-����ʮ�~�CC�&}�u��7�؏�i�y��{��{JE�4,�vy�j�J��J���1HS�ǜ�o�dF�D)���Q�B;��&Řg6��%E_k{��6�N��:f�sw2��P�lkS��IQ��s�@����ڤ�zK��쵧��A�B�1W1�t�;{ݦ4�}��?��7�7ߐ~�����\¾}��W��+b���V��ז���J>>����q�%������ޟ��o�!7fw$��M<��G�C��Y���E��9��h+����8��l�Ǳf;���V7mVʇM�����<�N���{��U֒���V��������ʾ�U�$��ȕI�TW�d7L�x��#և�)}z�\�xY�����o���*���oȭ�����坟�LV�V��������X�1�#�c�xc���&�D���{�k�0/��r6�Q�z��s�fy���0�R6t|��sL�=�hG�&gI��Ku�"���N=3��7���ޡ<���D�����"�P�8_aۢ��lU�&K
q��&w�o�JuU�O�WO?�G�c��&8{�E5pg��ϐ�7�"F���T��bf<�8
@��Z7����?�s�@�I_!�K����ɀ�TYS�Z.^$��r~��7�+���?�ı_y,�{La��k����X?��!�/�?sI�/�|iW�p����Q�ڶ����LOZ�d�^W};�>�����YAǳ`PE ]��3����^��L�����֧�o̶[c�Y�w����q����Ug��'%ɮ��6υw;�dk/���8���m�*{���ωʸ�}
���`�uU[d���5磻�F�K����6�kr~0�Y9�w{��B�3�`
Ns�܌,$S4�'6�Af��i���m�r*JZJh��M�Ʒ�,� R���ĤbSCAg� 4ͬhA�����bg�/=�L�\�Ѧ��\3=ZDkTS3�΍��{F_�)�;u<�(�im��b�%2�����fŜR�x8i/��L����U5'F�GN��a4~X_A9F��T��a.�i�X
��jf��h�*�� �t
 H35���h2����+b�z}\�	YV�(׌�iia`h'�B�OcYuqN����A`L�%\��e��R�h`��@�%8ޓ�@�O�s �͚<�Imz uW��p*8K q�aW�Jk2�v�h,ƫ5�t(�Y>����X�_6%�}���Xe���'Z�EZ#V�ƒ��n���*��pG��K���ekЕ�18#˙'`�����rvYA�n�y��AT�AJ�f^��YmW���Q��̙-&�1(�~�ܚ`�����'��ȍ�M8 y��SEm6�ÝS���O	s�ջw�K7�ʌ�t.	�O�Q�'�v[��KJ���w ��4�]y\��Mu])a4�lAF�ߕ��}�Q1_GqR�4��zҐ���W��{���񾜌;��1_ӱ�#���0��JQk���)��_e�|.��g�T�al '>J�Y�,�F)�{�f�����c��	�T*-�}�[ob`���-ŨR���:(�*Sc����r����u5U04�H�͘1|7��R����Ē��T^>��d�	���А�9������LARh�|��-;����k�\[V���ǌ9�=o�"���j�\+w7ƞ��ەޤ��멨���β�\+���#y��YZ[��qE&p�^Ƙ�~��*e�:٪�Ʌ�M��>!8�v�2e�˜���<�`MRE��X�{l����:�¨�4B�N�k2s�1��i�GAn�^��Ғ
�xS�s2*�1�~^bkj\����]�3�P�4��v-��"!�7HS�80�6���
��`0���f����6�Z�*̀�hV�3��"�Na�H桝?_
�^sl�vi�U|�5FSK��t-p��3\�
�������3�k��4�W�w+{�����6�S�gFk���>�;Wo�Ѩ/=��b/�������H�NߺqS�xn��J�6��_�%��I��:��Z�DN)&�,���Y�#���r��@�{�y��d&�N[��<��%��;փ��S�h�3'���?���U��
ϰ6���#ح��K�SLJ�\���`$�GR{�H��/�J�YU�����1�Y�c��Y�j�Ҭ1��γg��ɟK��������?�Z`
�4�'�@���h=*i�l�A�8�T�2�5ġ�1+�];*&�k�S�/ɵ��q�hV����?�g�B*�	�RA.:��`��\���̌�� �9�}����3$y��LB�v��W�Af]7ƥ;�c��q�|�2�ΫV��#{��Z�w����cB��X��rcc[.66 ���)�~�w"����@03�k2���<0J��Z�.j���`�"�`�U�5������*�R��.ڋ2Y0��g��z�9��P.9����4×�K�2w������I�e�V��`�w��2Y��Y ��g�~��D�j=���T�]�*q�b�"B������CU؜�tb���"m��L�D��T�Կ�~�_5�U��!��c���MB�����Զ�],���	����І�Txkg /<��;�N���W�e����ӎ'��+'����QPf#�	��h����\g������&�oO���AcDc\�pz���~mg��O���88�>==�ޏg׃�[����9�����.j�=����Y������5��H@�1F��5Y��5���1��C�A=�b�w\Up`|�`U-�S\˗4�P��Gb�����'�c��Rā���+� x(��#��w�(+��ю�7��\V��ݩn��)6���!��O��E'���1��8
�|8�y�s�J�$�٪FQ�n�:p�}����A��u�Ԑ�LI�	!-��;lK���q�M�N?['de's�.6䕋WeuuM�ʯN>����/��^�-�Y�������١\7� '���G���S���#9'��BK��M��F�6+��:�@͵|C޼}K.�x�3����0��9�E�ܨ4䵕mY͕P1�t���o�3�n���)��:��+r��u)0�m�r�lO��M�ڧ�q����s��)���Z*��BIV�#��h�ΦS���1x{&���rA#�����/|�4�R������)�������S/��LL�Z�rG����|��M���ѳ�G��s���������K����\��H~��W��^�#�JAEM�p�E�V
zhe�3��l���+���_zMtc���'�ݦ|�{ߑ�QGk9rX�wo�$_�yW�VNa`j&���5||�k����u<<O�x�JA�L�on�|�������q��P}0c�vK%R6/�C<�a��xO��N�P�8����Z.1G�dp�0H�ϝ/�r��@V���t:3*m�q���F��쩕Ҕqt�岬m���?��\�rE~�uGa�<S�pXj���xZ�H�JF���)�Cqi��#G���ӧrayM�)���ALkNJT�
4�s��`�U"�z��9d��3Ql��,Y�+� �}sf�OG��p�v���)�7��J�.�lQ���!Ն5d�&��>o�
Qe2�5�;M��r`��<�jχ��*�f}�v����ג�nJ.r.j�`_�'����Ǐ�礷ז~�+7o�V�`�َ�eVN[�KT˴Js��Q�Q���|��f���l+g"1���8��0JpJ�Li�r���Z%��")sO���߅���:�N�ӧ�H�HW�Ck��E}7���B.#B�1��h�����9������=0['�ux[S�8�H:k)�1�ƚ`�;鎳�Q�e&�ƛ�Y�oEs��>��ֲM����H �V0s�7�I����T�v�c�)�D��K��(�#LTvW锤R���1T�%6 ���}W)変QX��E'b�������Cy��ؗd˴�e�gq������B���գG��O�OmS!JÞ(m���&�	3u �#*㻿���~�~Y{ι����bV���,����h)��)+ь�hL���p�����꿹��3Y�-O���w����rq��F�{�ʸ6cOp���y(�������m_Г��Rk�<Z��M��`�53�,<{	�j��`�\�u��>��:U@�z���G��{�ܹ��V0v9�_��0ʕ�-h�n)���@�A>�n���˳���^���L,g=�b��N�d��P2咬�o�OƠA	k���1��ӱxx�N��h�{5a<ұ"#�,�:{PR1w}{d,>�/OƧ ���R@&��ȵ`�s.�eZ���)�V��uy�e��u��p����p�M��X�>y��,�e��C��=QZ%�(I[����8��?��Ğc�q�, ���g�<G���U眉=q�qtR0j2����-�Rzz�O_�0�|ױa<%����u�b������������i-�X(���V#dA�u�sGĹ{vRb���8s'���'�Y�r8h�;�|��ǿ�<n�Ѹ֖������������?8���M?��aw��<Se[;Xvi}.Chb�Ihb�g��w�Ba$�QÌ�	W��~��#,��Q��܈�i�[y�<zs$�9N[F�yߌH� �}}��lz%iDYq@��Ôf�+�w�Q�F?#_�|]�mk�����&��kf�OZV��L���#ǣ���.kp�3�HRa-��T��<�X��`b������?�p�w7oȋK��l'��~�|�ޯ�p�%��޸*��oh�����L��#��=;^��d����ё5''��]���ܖk�M���ؓ*���S���'ҟ�C��w ��z�vu�0:ۙ�������l6���\�G�q9�d��+���T-�2	�ڏ�n�b�!wַ���WS�6�����:�C ����4k�>�c��OT�3�Il�'F�:k� �3r��*�/]��ٺ-��Q��*Tӄ��X�]��W��7�k[7Uf��;6���^��M��G���@�p:3^U.U���%���Ifړ�������Jmw_V[)u�r��1��?���p�}��Eb/�B�Y��|82��c!x��R^�jQ�)�+k �Y-r������Odc�B��Gj�rX=���k���Qخ����[RL��D��r�E�]��%���0Y�~Ɲ�W.ߖ���=��h��ߘ�����ӆy�YW:
�w ���~S��u�A1>���%�޸(��P�����C!���=	.ߒ�8�K�c�TЌ�[-̉'�K��cD��F;FγYC_��d��G�˓ݧF܁�,�'p�E��c=)����F��{����s��[���b/3C���Q Pz�S�����=Y�5 ����HZ(��==��ڤ86�6��z��5KO?�����#�NǨ��zm[�0��%s��Y-���y�LJ����o4V�����T2�`��{��f�@y�}�H2C ��,���t�>��*�FJ�L�����!�vL�LۊD��iXN�9��sr�����ʊ�m����|��1�����E�zv��� ��@�t����XF%_�^�����p�ve�j��K�a�O�}N.�N�̃�c֚IgБ�Җ�8�<�
P#Rf�^�~	���28E��@�[暕๦�"�I�U�J�r�	�z9�3(�Az�
~D&3��[j�M�,�}�&�@����g+�IL�*zB�F�՝��J�Pm�"�.
x
u$� ?ڜ�A,�na�V��]E��W��t�I9��k��̾���8��f�٨=�^��8P6���0;��oA�>L�T%�I��M�N"VI�L�jq?�lG���>�qb���};5��j �}�Yq���`/�-I2���_��'Ӯ������s'�-�_�|q����ш�"�Z:���뒁��_lb_��U�	 Y;W}	z�,��UЇw��~2��A� ���l��xbmѤ�Q�6m�Z������hI�f�9��k�����@
^A����8_V��
E�wqe�=�f�R�}�Yc`���A��*�p�����e���M����K�0l| �w��UWm"��:rM�,K�� ��i0�Ns���:�q� v)d�Ҩ�
\)/UdW*U�E�Ӿ�ǰ�����)2t2�s&�ޗ@b���k�Ȝ�W$\0#��/���u�`ޗ��&��@*8�_������u}[�cO�ѩ�0Fe��b}Yj�C�p,e��j�"]o,���F��u��W+r�����U+�sϡ4`�5m�8ԖA���"�$i��НӌSZ��:۱����]��Hh��7>,�p?���me�X��������?�|f�3M'��8��-��es�>"vο߶���7'�{Km_��#iG�Upu4��f.9�o�3
�0��!�f)U�B�t�|��}��6l��|>��L&c�,��g�`������[���eP-2l��$�O�'���ޣ��'�}��֓����}z|r�`���Y��٨��`�p�N�wѻ2W~.C�,��Q�șx�c萶��c�W��y���h�����<ّ/�H<��y���t�f7����e�2.*����Yqr�P���N2UC@�;���BM��<���w
g<_�%8��F��������>�t�P���YY�yr�3�g++�#�͡�aV�m�K 	E�1G3��,�\��H+��~(+3WQ=%��kyٖ�Lp���}��ٮ��DJIM#5����	���n�ZyE���rР�QG�jz����/X��r<i/�W�|}y�Ԓ��F̫pJ�k��f9���z���t=6��������|��M�T�=8	� s����3�p�0ڮ�WKeqq��ͤ'tx*o��t� R)=�
?H�hAQ��U��\Ȗ�K�nɝ�>� s|oH�#�$�Ey�j%�����K�We+S�	�f���9�ۮ5�dr-�'l��p��o]�&��_�:�͓#����<�+~Q�T>O�1�ΎQ���ٮ�ȖW�,�Z�>��~�%�\����V�Z]�Ĉ��]��[�4s��<�N0�R�#Oww���Uͻ'�Vk2�ً�p"�ܚ�dL߫ � 1����Q��`c��@�=�/�rU޸�\[ْ����xS�bV�;)9%`��	B���-_��%�c|e�u����.����_����+N����ޗ� N߸|C�6�w<S���ɚ`}����ϣ�~�F��C���Ƽ�q�hw��<�v���<ّ����ـ����L�7FJ�pN&c��= �HpH�HH�$U�V� L�;��-ɼP�����V[����`(�9�Dk�<�֤&��I0���9�H�Z���S�dg��p�2�	;o��g�g�.�f�T�'�ӘQ'�M���¬:���h��%u����/w�6��*ii�X�� Hk���3yv�T��!gd�9F�.ν���q�NfF5�u<nF����Ce6���'��T�u�f�ju�Z�g�C������ކ��t<��r�.+�/�8�6��{�
���y���㖇�6s���V��$iV�9��bFV�)�˪D�hpy�!I�H��,`6:M|mN�|?ΫB�B;e	�9I���*a�I�3m�g!E�W�F�BI!���G4�
���]ݾ ��(�s[�5��l�J�N}9�T��(3�
z�����*] �+e����D��/����4c�ZG����t�j�u�s��V�Vk���'��<���Q�� �:�J�g882{�5��c��$h�8d�;�HC�-�\h=�њK#�m�H�_�����+.�TG�� Fg�r��˰ew.ܐ�򺔶s��d�P^�C9��!��g�܋ B2*8�:��-�Z#��u�L��&��q�s���c :� ��W���"+;�߶��cô�*@���KbDQT���l���@U��0�iեꇬ�#�goM?�u���v��"�/���Em
��y���fM�dǙ��r�-�������n���@� ��@��0��A��*��Mf2�L��2��p8$� 	�X�ꥺ�-����Fđ��D���Ƙ�8��3+��XN���?��?Ǻ��T��!�=_�pP��*�`��p. S2�F"��,9��>���v�j�A��
�@X�n��82{)��<Fg�.�;gR�fE��k��|���ZJv��K��5B9�XA`�$���c$��Q���	�iw��D���Wث��l�ĉ�nQ�~�
��ƥ+��h���.����u�����Vy�b����]#��I�ӧ4:y)���\ ��5��4��CIJdLNŴp�XyϮS�~g��Ҫ���u�r�s �KR'� t��~P������}��i��c_�;�h��_�s����sY�,C�3� �{�~Pv����i���ښj��'�>��gM��&�F�
SH3�*�ٓK&�>`4 �!H
P�	��B	���/<�1�L{~����6�� �cY��������
�E��{'/���\�=7��x�[���_:���x�:u�w:���>�/���x�C$i�[�M�Ӆ�_;��V���>uɈ%�.�� ��ѭ�<����?f�V������9~���g����i��q`*s_��R@�F�uT+� ��҃�t���9��t��N|cUj�^�����L_�z*$�����Jҍ����"6��bJm�Rm��2�h�l���9y�9f�t.����/�Jǋ	�N�>��)]���g�����7�(����/�°���Nz�yJkR��k�@��B(b����P��}�UWi��u�g�苣�}��o�6���Z٢O�i����\m�Ș���3����vV7���*��;������6j/Av4���}g�*��w�6��;=*7������w��ZdsF���
@����]Z-��	��|�+z�N�bIq�@7�ȁ�h�؊:J��J�?{��t��B7�y�̍6�N��%�?�r�+<���_i�1����_|N/�G��·ߢ�j���&m��2]�����5
�)/��݃t��!��RXev��\f�0Ecq�sB&����y%��5�x�FM�e�,}=���+�N���K�4�[Wo�0B�ਛ�h�*Ӊ���)������Ac�FU2Q$;�1x����H1z�?��hHŽ*﮳1���O�}B�g��֥�4��`���k��`�F��.�g�P��cd���~���tu}�&<�Q�۟��8���7�C�%`��[�O�����y�2 �n��>P"��� � 9c�7<��:Pz2ȡ��q ��%p4H�Qg %8ۧSv� ��!��h���32P�g�?w���1�� q��	��h�ʹp��.��"�ʢ�0�{>��>m��Ԭ4$k��8��h>Y}e��:��
����.�}E{�Mc��Jm��$.�b��**��HZxH�?P��>@g��U�`�1E=݄BO�q�*�8/h��}��X TBLg4�9hL���F��%"��(�1����Fõ���H� 1���I7��R�QO"��h��H�=)�EX6 i6�V�N��6}��lҠ��y��|�l��pإ��=����hު���dD�aϥ_&�=����^�^
��\2��1�����u�}��S�@���ؿzZ�cGt��J�P�p@%LBO��C�%���`{y|��?� zeB��ͣ�·�6��y ��tXg�Th�(�9��s+ȳ.�Z=瓄Jk�vj���s�Ns�Q#�+Z,Hcu�,�x��:�Fm�{J f��DH m=d P0�L�=��!k	h[���@_g�!�e��_�5�� �]J�=�6l.@���i���߇�TzJ�ʅַA��|0M�w�=
u~���%P)#i��C�����U��׿I��ݠ:۠�v�n^���nΠg�s�H���Q��-��u�E�S�(���k�)�<��mrI� 9��,�ҟ���?�rRD�+��������X��=���  �Z�D�)՛+��= �X�<�8���F�S�ٞ���
c"05c(�����B��,'�%�h�X������`1Z9`JJfu��ooC�r#�4C�v���c^��,�}ۀ�(���ۼ_ �y�@��v��k+T[��=�z4��0/}�p<3���� �i�G��P����E(n!>��W��-
�;-��ǼvyM-�I${��ZigR��V��u��u%��>�6�eǇ��?�1�y����T�!���TDC��m6���c�~n��J���Q�_:j��~>XB�l�ߒ$���iB�[j~�ʻRs�3�{R|�_?�˒�I���m3.�5[�����-�t?�J*���Ɣl�.Ʀ�)��H�xK�_����YU�-�ہ@�
E�Yh2Z�m��~�t�%�GY.�\㲈d������v�6o�D��M��D�������/��1?Z�ع�G~=�>e�o��O'��������M�6y��~�C���K2����3��%B�7%�� K�l�V��v�\�W�[�0��7y���I����'֮I(����q���w�����;��ٛ�=jDw2UJ^�<��~2�{D�̛��H��2����͢� (c6��z}[j�fUj!�?�{�/h��tP�{��C��Wt����P��+����Y��3p���0�P�S�b�,}�޼r����&�������;,�aZieЊ@M�>c�("��@��h��VS�`�g���΁8�hr�z�)�]p��,@�=�N�]���=��5�]f��N�Vk|r8*�J��oܺK�B����8���볃�oš���y�ݨ��J�ǚ7P��y90���:�b�*~#_v��jy*�}i@����%vrg�	�Rxi�*aA3�����P�W�2[�N4�g�cz>��&�g�q+\e�T�:o.�qLwo�э�K�4�c|�>�ߺ�����_рi����	�d@Ȏ�6f��[��w�ַ�錝���.]�v��<����j1`�PcCD���{רT���3z���8X�B>5�Dx6)ϓ���<�7�����Z���������E0��ل����3�(ׅ~OR����TUlԠ��*ui^��(�xL�dUm7We�����l�ʛ��3���oӿ���*<���xؓ��=�`(؎�9���ʨQ1�GcaS�~�gBB�ُ�Z��J��2�18~��	��@��!v��D��j 얭k+T��fj�<<%8͠{,T1X�&Ay=���"��g��Y���]�hd���|,�7QG�)�(��(^�q������/�A���;�3��]� �^�V����#v��A9�*���G��1U��@;eq�X�*n��AZ � �3��-P;a�737*h �p$���s�A������� � a[u�Ϩ[M�o��#�l����ԑxG�FmM6(h��j3Epa�sh �gQe��!n�f�O��ƶBKh�1M}�Gq*t�)T!! '���!� b����A$"^=�G�h&���#�&���Dv�S��x�`��T#� �v����$��A�����]��|̅�`"��A:�RR��'?�*�E�H�N��� ��>���V�* ��@�anI%��C���jH�m��k�#~��NU^��f�6+Ze�]c���y�RY�p��LZ�&uEp�p/����{�DlK�9��j�kZ�/������<�|>;PoݼE+�k�E�-]�RV��ܕ�:�4��y���$�%�N��$3�6���B ��
5�2]�|��A��Bl�����i�Ң�	�mJj�tB�v"*�́�H���=���$xKΟu��̩_v�-Rt=�2"���;�oۈx�?�۷�Ǡ�c�����MS	������]@i�����[��v��*���􈞞A���)j�p/�E��賏к~�J�`��b�)juPz��uVfo!���F2�N-}lmu��.�1Xo����%@�֨ӄ��h�р�^��:�$�xvF-^���lԧ���ZQ���󊰫�����B* �[�)|���@�F&���xgh������ⷝt�RS�JU�x�8~I�aGS�7��W/�P���^+�z�y�{�;��t�������}:c������4؟���K��b��t�e�c'���;$�
t�����I�e���U�_�Y����O�����
XR6.98B�۳��g���.o�1�x�WB*��qt@�h��P��Vb[���Ǎ��X�#� ��b d�|.�����/���Ny��3 �h�6�b���r�.��xNU��m���[Z��4v*����|�Ǵ�8.�\�듧�����h�J����0x5h_:���Ť��$��ø|1�}/B�@Q����R�6�l������/�{��;6�,�l}�ճG�8]}�4���_���}d��x�����V�?��2�Q�h��x�
��[LZh�v�'b`C/Է B��k����#^JB�&M��){��mT6���봹�+}�:�>���1}�ާ;��'�������o
���@@=��i�āz"D1b��J�
���G{����W��Q)B���
cQE2\�@>�`���U�BqD T����G���bv�G<�?{�����{"�����F�Z�*�)*�=�Q�q͛ӄ0�[�.e%(S�V	4�
�ݹFך����|�ycs���� �"Ϳ�Ⱦ�Rs6求Z�|�����N�iAd��T���>���#SxR+&J��&��d)A9x��������������-l�4��Z����bZ�E˃t2��-�kֱ��{.mo

�!��>_���i\[����7(����gO�v�Vy��>�{���oз?�m�[Y��~��_���{�T�1۾������x#��y��\GS::9=c�9�h�ʎ���@լ�����&�s�:z�N�`D-�P��3P9��i��Ҹq��3v��S�{����x��4�D������z"�R� ��Ju@�A]�~%*�S0������?�/���ì4�S���6u���kMy��G<ƝU�5J��ZL�*ε�D&�F"�(X��6��a
_��F��h�q l4��FhO�'sD6�N>>W�Ѫ�&N���x%^�M:����bPЀzd!�X"m�!Q�@�b�qJ���I�����u��V/T�I�4��?;�U�M���g�
�t8T`�tA����O>���RS'B�����QJ�)ʄ�5�('�'�<�]���H�,i��K_������� ���78���6!X�Z�j{��Jmsb�co��Z�Xj��T2eb�=��U٠ r6�Ȉ��fR�[��Z_��Ϸ��lC�Xq�N�L�e��2�XEK3��"���K���l�oꫀ��\����7�x�籍�!�!��<Ó�|~Q�O���s��)g�&�^[�`T�!o�H�����/�5�C�<�ИL!����~��%��6�������o�`��@��aUʓ�\�&�v��(H�"�,` ��Pa����c@hwN����ZE�zhm����B�m'0�l�# !��)�|�9T���O�����e=���d�y}F�Uxm��%R4�
�<_#���r])��~kD��u 3��e�<�"�,_�Iټ�Bmհ䊟�����t�r�p}�zKΫ�����p2F�D-Ƽo���ɤ+�
�;�ۀ�)2�V�tU�O��fV͔ʋz���b=����hfJ��E�[J�"uU{^N�sw�iˑT�>9�SA� �g�/h���~���A�/e��v����6���{��
����P���ф��)W�8�4�� �1;�H� ���ꂏ��"�=>���n,�(�:t�����Dޠ8'���oK5�mا�z��UD{�Z��{N%(jЧ�e��XeP �~��"ꨡn�௠���FaOj�{/έ�4�/��]�>�ssӽ�h��E��˔P��ra�ԩݼv}����-�;{^�D��"�0��[Z��ʮ�f2]����B�I�:K�P=P�d|��b��(�$�D�D2�b+-(D͠�2�I�X����9q����(�ʳ��`PQ���JP
���'��Q
�z�D��Uyk�������?��zy����nI��y:;
�<i�f��φ���d6�ӓd��iWۼ�ӹ$q ����s�>X���Ń�A����r�:�o@�c�}�������q�_�:ţ����������?(�W�W���䈢�u�d��,�݌6P��0�ڱ1f�@10�7	��B��� �d�-1�bѱs�]�һ��i����ӡO�^ѣ�	�*�F�P��V�U�b�6�7wߠ��[��#�&̜����yq��ȓ�^�08��Y�C[��4��Sl���:��~���GCj���3[����z\c-�!��^~n ���E80��c!ʶ���v��7�@���Ȭ�o�:�1���G (9��NqJm�r ����YŔ�\�L�_�Mv��3@fǘF���@��Q�nA��P����0�҈7�Ƚ��@�$�2�Y����Zc��Rd��	!�������gCi�>�~hR�8j�F���
��}�D� �O{��xuzL�K�U}��6��gfFe��"|P@+�4dpTz��v�R��}~��tx�R6Lԩ���o�ƍ�<nSz��Gmv�!4B�<ϧ�z��*���G��  s��E�զP)�fD�f�Ny.T���=e`ycgO�B9;^��ނ�*v
ؙb��/����OI�@� �>[E;I�6[����_��?h���U�-����m�Ц������"�s���Pm0yz#������1���|��	i�T]�Q�T�sty-������MR�9i=D��� �P�f�E �5����c�~�p`_�1�+��$��U�Ⱦ��bN�قL<�+�r&mV�*l��N�}���ĳ�fc�F��X�(l�j$�8���;��B�CT����9}6�����b =�пk���F_���)�\sE�kM�-��#�WZ�P����d<m��,H�b��]F�a�}Jm��؞M���U3�s��g��Kcr���n*�� 	(���r�@�h���t�7}��S�����`�91�)����v϶�	0q����.AO�y
�;0*غ!��A����%�&�%Q�-�B-�ݛBQR�	����Ua�<Ml�Vq�mT[(�9a[��P�+%^�e�K�]Oy��iz;DMRK���P�EYv�s�r1��d<ɜQ<�4���}����� �ԋ�����`�'�Z�.������{bU�=����L�yY@`�L��q�:�%�=�1*�}V)ȀDsZl���	ve;��@4���5(�<���L�_�5�NQճ�U�U(�J�\΄evŷ�Y��q54�%���4�������]>�Y"Q���^s�_dm����Ԣ��!�s֖,�Ua��7�爊+ɢ����4����Ȱ=S�7<�EU�������-�sw�9��A�#�)�������*��AC@;��$� '�/ID�8�}Ի����D��TC01�!�t`�6O2.Xg4і�R��z�B��.%m{#�m�{�$�ca��p��@`�)�	��-��t1��A|Q����1��Y	���@��T�t9����'�M�8P�e�}D�ȁ$�Y�2^_��+�/��s!f�|��Y�������O��#��!<�ǋ�}�Fi\��1��A�bQ�Ee�sz*��yY��ԁh{#���!�Ei��-��̨q�*��sD9쒯%$�fA4e[�M����|��s{��5t�A���	jg��X����%eT���dZo�J<�|s���k���'���l5.���y6�&W;}����^��u��?�����i��{G���z�o���Y0��q��s[ӈd�炱�-5��%B�8�q���T'G�j�f�\SY���I�$���Y����K�%U���n�����WI'��������g'/�}9��C���F/�P0�Y�iL!u�� ����zX�k+���e�n�Z+��a<I�B�-6^P�/�͵zk�
5������ӣ��xڦpg������0��A����.m]�̓�W_i8l��\HK������x�!��\cMd����j�s:��Z����\���3џ����V��E����i�R!j�EIO�P\#u��^(�AS��yJ�3��q�������xe��ⱐB^�gP~B�x(�B��i� "�C)��E���u�i4h�%�;zț`�6{��Y�yϦ<oT��b��❃��A[E�;l
�A���^�6فC���P��ltB�JB?x���~\�U�Yl�A�6^�/-*���BN�):��BJ@KEѧ)�w|�P;E�ݦ���ID��8͖A�$:a�b7ӵZ�W49��^��S��Rz`��n���hL�g�tum����ҷ�w��f�3�w�?~��|`3�`F�N6TPy^�Sg�����g`�A�|��[ݦ�dH��'4/�R���5!b��r���WG�E�h�ڢ��U�u��x<g/,�*s�%Zxm����#�ߔ�}l�?�iȕK�E���\�?׌��u��l? ��u�ͳ�I���A��Ll]���L��0�F j_�N%���"z���l͏�up��Ǡx�F��m�d�˪�4-�o��IEL�Ql��!�BM�$�+�Ƹ���M�,�Ȇ�
AId굮W�����`(�Z ��<�!,j��3� z��IO����4I@��니� �d�<#���e���r�������6-@z�	5�g�i���L@j��0g$C+�yږ@�&��Sk�S���)����㛻��P�"D�/Ԇ�^���R��p-�l��)qۦd5e�y��T���A��䙣�'���61�E�
�Z�m�����N���$Z{����*��sLl}��-)e��d��نkȎ�C�5��\3�j���B��������تS�^�?��5��(����l���o��z&>&z�����ԋ�b��Y$�Ej�
� 8�2�=zt�~��D���#���:��Xc\���y+�����!5�O	`�=5�-��G����
��9�-��J�֚uQ�=�Qw� ��v<^��Õ?�zj��D
�ܙ%0���K4R�7ϵ��A�y�!K���s���j?��Bڲs �!�p�y�Z�}D �X��	M����'�l@A�WT��X�_ԙ+�pZD���Em[j)m�I/��[�<�\{�t6�
����CN)I��g��hŠB�zK����@_ Ϫ(ʬ����%��^��^��}1SF���S�R5HU��G�t	�$�\3�?�Vέ�+�W`[AIYp�z��N-�~N ���ZM�g(�`�(����I;$�!�6v.�J
z]��4X�ʼXC({Â����5i�ȹڻep'wb�;��ʿ�9O�H3D������e8��{�^�x���+�U���{��r���a����q|Ҳ	�3��F}�rC�n�zD~O5U�'29	�>�# ��AfГ:�.��c�W�K�A���Ƹl��:�����Fc	���`$2Y]���b���������p��ɠ��;g��ǃ��
A��>���p�˸oAՠ�k�Xx���?��w����x>�4�N��F��u����ʸ�&�<@�g��d��~�b�����|�p��A������LQ�3��ܯ���w�щ���+c3������Λ��-)��F������gӳot�����|��e�����x#��j�
�>�c�^�Ӈ�~�j++�� ��r�>=�����=�<�3*�b�Um�7v.�ݐ懇��������6����i��@ѴuN������f����>(�]�2���MK�:G�R=��[0(ESذR���{���]�M�hf~�;�`@���槳����eک4�VJ21��=���J=�'2�a E����C�	��|.�&�4<��:� �	Y�;�Zk
�B%W��489�WO�Ѡݣ�暪��J#(gh0�vȀ҈3$�ҌY���^D�1��|5�n��w7nҕ�)u�^�D�`A?��#�dt$c�#έ�/�f�1,���ф�y�a�P��\�A��4>4��(�HV����-Hh� 6��)H�W�UZa���vkCh����f��4�ߨ4D�brڥE�N���^ߦ��9m�P�;�kW��s*��es���x�,�v=v�N�]ګ�э�K4��J���BM�5P�=��iR$y�� ׀:=�ZBχ��o�����?��M�񟛷iҡ�ÉdIE*���Y�م�cd���,J�mD����&+v@1u�����&�������δ�r �-��W15c�i$VTl|<�1��Y ��e�[��IkR5@}�$�QB��6�������HjאKlỒm�j� . `#5dn�f5! ��R�asK��m������3�=�S�l�Q	{Q4-�֩j�����:à$��p�}K-GTA��a�S�E>�i<��A�}H��:ǆ�6a^�
��-�B)s3�1w�qꊦ�Ͳ�q�lZ��6!�B��G`���񔾮��+	�N�'iԖ�y5��K�M� �2Wp��·�����4��[�*��	�Q�?^��x� d�R�V�<������h�N.��88��mGQ6Q�'~VB��9/��"��eT.iI`��r��J*n!�z������Z�Bg��ڃ��,��DV���5.�@A���Z�&���n̘3;�]8�R�:hI馈�#�Xѭ��ba�9|�%u��X�����Xl�Һ1��gD�%CKk8�d0ՆB>`���j��hAU�2��b֥)��d��q�9����J��.;�]��aJt+�G���A��C?�%�_�u���Z�rl7��,��5z-չ�}j���:�x�[;V���쏊ƀ6&"8�:{s3H��TDMa{	�'�@I�>�Te?��p��ֺy�䎿�6/ �ݯ}m#v�h;	��w�#{��kdׅ���G��A<+�Bl2W@� <�H�x�b�hlBA�h���-nV��B�?�G�O��ҭ��S�٢�G4&D�v�e�7rg!�T��c9��,HfH����6�6j��7$�@Uzq����F�j�~N��y [��E ���=�5o8������2���wn��5�������S�v�� �{vJfK*��k�su��,h�e��-bY�F�=���̰�E��0CVJ� ���\�ڔ@E�gi)����Tt��,>�N�s۷IڕxZ��1I��	C��Z��b�d��ߝ�}�����ړ�Z��Nk�~�X<-�'�<�_�����'�|w��/w����|t{��o�(ޛ���a��2ߙ�j$�����;+��.�zz!�^vV���O�zpC�U7���F�q�D8T^��l}����qR�Z��rd�u�?y�hxԾ��Y�?��/��٫������qV���{��� ��k.*�vs��Q�����hg��^�Q�$0 ��l6�G�z��I��ZQT�D���͵Kh�^ѧ�W�*�0 ��� ���3��O|zrL�8��h"M�M�P��4�=�qp�l('I*t��P(#zuv@U6r�b���x�6�-6rP4���C�R�V�����Uzkc�j8l4����1@�������a�^EU2��Ǔ�"�Ev�z�Dͱ�G�@�#+�Y�pF�9M�d�F��V坍+�6h�i�،�{�J��#�Q���Gt���1�PP�t���g����3Zc�� (L�?�K���u���wԇ"��<:��?[�{ApD��O"!�W�řD�"���ѭ���
���W�S�����4��#Ω��� ��R�7�q$��� q����k뻴�Z�hP�ӝ�7���w$�^rM>_:YP�ϿΛ� z��U��@�O8VB9��wԫ��)��4��7���EIuN5vj�?vE���;!D"�s�sPm�TfP�f��ٍ�:|Ioo]�~�ww/�g�O��\Z�^��=i��TJ��m+T�}�#��c�+�P(�:�~M�i	$�%�:dD�`��n����g7��(J̯��9��C�|y�'e^75~o�T�xG{l�ʄ� �Q\U�ĘJ=��-S��$3�l�N�3�)N6�	�Q���ZY��pN����J[����0u�W�tb��\�Z��I�T/��=���k�`���֠�7By�,�Jj�OX���|Ю��-�6��9E��
Z"Cmb��u1�@�+�z_<d�E�FA1N}�KfM(���~���Bc��*�u�f��ǰ/T6@j�P]�9e���~r���V���f����xN�;?�J�e3��-OB}�8A�Q�n}��\�N-v:Q�}D_���f�J�_�Mw�����OF�� �⏦���LfZ[΀[j����k;���R��� `�z���!�5��GD��q�Nd��
�R��UYz�š:����SUH;1'e�0��Tb��,��4�W��hD�(`�]pW�ғ]�P�I���mE��җ<�y�H�K��)�&��H�0(�ZF�+��
��_���Tǳ(�wC���"H6]LQXʶ���A���x.�"��`�9�����о,�u��ӥ��q�?���\2��QҾ�%6�����kT�?�jU�;��D��m��{���R�%Pdd=a_Nm��$�W���픺
a ]������V�5���l.tzdQ[�[.�I����h/w�]V'�S�e~���������.tD!+�6?������7�h�T�!�$ `	%R�����N�5�`3@�+�s\���"a;����D[{�L�uOܷ��,��h���.s�?_ʲ�X)�������^>�����W������%�W�"m�|5�9':���}�q�uk�#��.���R7ٿ̅�_�ZhGku��~ς2����<3�u  IIDAT[�w��.��S�,��/�	�VQ�$㝰�06���y|�m3z�BUI���b��^t���S�������gW���eӀ�?�R]�y����b/��>��ە����QoZ`Q��Q��)����7S+S��w��Џ������P������xV�f)+�[�|.�c-1����p}�h�Ѹ���R����g�kQ?�`=�T����|�1Jgwk��O�'?��������N�9[�����_Ҭ����+O��ֿ��/��L��-
������a<�9���w����F��ŵ���+�LQ(�C���k��Ӱ�"(�2��Q�)�&��8�7wv��훴Zj��K����qw�*�"~���x���30��3=��c��:�VD�P*r���f�MQ� ��);���B\��8:>��ƪ����ڡ2Cԉ�I�l��!���'����EJ�&�DQ�(8_��`P���[�p�gSq�ZP=O_ҿ*���`����2��#�G)�0�خ����D@gBsK���M��*"�v/ѥ+{|�4��b�`0����|�������'?�r�i3c��ƋY����ݰ,��#�zĀg>�� ն��b��( ��.(mP�2ZC�n���g0kꁴ9�ri�������J]I�ⓟ��BA@�w1�&\�^j�zB�r��E�~$�h�T�ԡI֪^�񩱃�cl�^��H�ClT�������N�k���h���Ju�y_�MA���h=��I�Nz]��m7V(����є��|�%s����|C����.7�sg���0���^O�"�����}>R�d�𥞫�s�3������@��D�_5�^x�3<�H��
�Z��p�A	�h�h"o3���h3�n��f�F炨2Z1��:"2�,5�(�X �� љql 览��`���.�T�p�)�����lk?3�w,T��@��I�Y`e��2*�ɳ�����J�+���NԂ�Y�5$�ߗ��$��=�"S�����z9%��p����F��2��A>/�hZ^VZ-sQ��<�y �[	G6�l��QC���U�_����j�$3dך\^�.�����J�����|��ؐn A,dF��fBK�������"c�Z�VPQ:5 U�pd.V�q>���\�.��9����<�4�o��.]���*�z��.�r���}������Ԋ��vs]Z�����"<�����穡�P��c7�mC��*dl�ľ�pf�4@&�w�w	��U��F����,#X���/���F��cK3��`hkk��P{�yz^7 ��-G� �'}~Z�����9���s��]ҵ��(6[@��{�{��P�g����s��VE�UĖ
Z:�h6���D���A�P1E�rg���	?�2[���7gNf��Φ�
t�2�뢖�S�S�z�36v��K��@������'��������F�4�BGQ,�� Ռ��B_�ʘɪ�$$u�x��Ћ�+袞��S\ ������Y��d�G�P��l��|>a���"S��E����6��C�P��'G�k�,
�yc��G-�@YZcɾ�Q�T���3s�[ؙ�KR�?j6R��T�Tp����p�w��s6�3u��`��Y�~�d]N�;�.��� {c���.Ρ��x��� گq�����;��-�T�=�¯�z�v�|���0��匢�e#��/�7C5S����^� M�2`����K���-i@Af$0 ��*��g���dA��-O��z�y�{����!7����%`�/ے�3`��^)UT�f&,�4&�:��:�[�Ѱ�gql>�GӢ���v^���(�N2Ȏ��������ܘ�-�B$p�j� :uQO�I��<{0|DA�'�D�
Q�%���W�`#���,�~�}����/`�?z��nmLW�+��0������מ�zu����7z��FT����'��^g>���	�p�S)J9-?�D�y@���`V-hE�20��ΧB?�T�;/�c\]����e���wh��B��3z��)������u{r�|I�i�=3F��4�.�c"�N> ��j:��
��8Ѩ�����:������c�bܣ&JQ#I��I7d����}���*N�3�(���C��)Igh��]kn���@���l\�ĳxLSd���e�M��UW�b�A�Vy��,թ��	�]�|O�����8�(B�A{�"�-h����c��Bb�eO&���Ao�X���E����g�����+:jwęE6p!�41���|�������"d�PL�M0�'��Ǹ3���e�\���*�GZ�M�Vũj�z4c穴�N��OҎ}�.�nKh�ؐ�B6�4B�(m�פ�y�7�ބ�D�g{��<��.T�Z}��x�����uFԼ�E�.?��J���]Rpo����d������a�.�V��N���)���P{6���M�����u���w郭��sD�~�)�P9Kiu�!�> ��ӡ�4l_���N�,��e��6�'��t��u��ؠ�W�Q�B/ڔ�a��W�HQ ���d�=�BRA��>;�[�z�ukf,��檶�(��J�y6���@�*�o��Z&D�a/(�Hh^�R2�k6��0����c9�V�v���9���@�F�z<*l�%�"p/ȃbz���Uf:̞�7���M��k��A�D�yv�d(�A��4�� �n��o J�%q��TU���4�@�T�v��=;�B5
��qmC]d��A�ؓ?O�Y_��B(t�����5[�A��./�zj�a�����6]����]�`��"0�) ��	�����O���#]P���
��ߤ8<�1%�Wڭ PO�O �c8gU�?�'��x�\]ߥ�2����������}����ջw���.�VW������)��G?��3�˗��U)Ik�R�J�|Sj�!7��8�Mگ�R��ңL+�#θ=9��7������m��T��g$�4:8LO3O�t��`�5v�t����j�dl��߇�!��ZP��� ��N��Z͇�^�S�i� �(�u*�$s2���,�Bd4�7O�uI�tS$�}��n�D_����%s)<���&�(���*~���)�㈀��R{^9����s�[��e��d�u.���:g�����`����V�^�I�o�uo�7L�\�C p����:�{|��L ��Md���@��^:�{ϟ�����_Q�.��ɾ����N/E���g��@���*������v�;o���cA�ց#�/�Q�ц�5�͔0*���Z@��ml��G&��&`�����u�y�@D����B�Z[���7�s�S瓚�,�?*��!k�I�e��� �%���lf����z�l�._O���ǭ��חa��$�ޗ#1��]#^�љs�u����-'s\˕��;�깺Uz=
;S2�E�sߵ�f��l��w�b]x�ʲ���]�Ő!$�a�.���4K#_�,�sȹ��
�ˀ�ſ��xZ���(�r�m���Dַ݃|8+�&-�b�/j�.������eQgw6�-�L��6U~}�Y���B\"�䋈�P�H�B���N�-�hCT8��̱�s�(m�iQ�k��o�x���B�����?�{��~�T���ij�}�$`0YZ$qy'��A�_+^�T�k]�^:��*�ETIa�@$J��u���RVϐ
�X�"퇗���<;4�v����"3�I��C��n�A�]�+~��G]��Ѥ?�2�ލ Q���/;b����B1����4�M��
]��K��+Aْ�H�A@�w�iK�,6��_i6�1��F6ʄ������vZ�U�B (|͠����(Q�����
&��#j��t��r�Ȥ\�إ1����u^-���Sy���
�w���@t�є��� �����3��Տ(L�NƾU����?��>��jt2Џ?�9=�T)!���t�C�[j9�<"�����%�Nf1u�*A���+=�\�(2��L�l��F�e�"���;*�bڧ������}��۴��'B�͖���Q����+y�oS��`�A���m��n2���8���сd3Z��ڽNW6wh<ӽ���˃'�`��􄯸����u�����J���:��{��\��d}���G����Ɔ�n��3p���xl�� ��wF{����~P+yn��ֽ
��{���u'�/x}�2�h��	r����?����s��ml���'G��ez� �Cڇ�(WH����w������ �3��?�OcЖ��#��IjP@�E����Vѓ���@&1�%����;0�*%F�fz5K�l_*_@�O{�Z-T����?���.�KA#ɢ�;��ʥ'F�����"���;Pn(3��Q���I�����>j�� r�K��S�3�l���+@v���BJ�*6�s�7W����#�B$^�@�p����`hl[�d�u$a�Cߊ���ۃ28d�i-S%I^��J�H�����Ҽ����oQ%D@Ǎ1j'suf�R��wGŒK�c�M:�B?��P]̠v�m��f��e0)�l�������ulk�R�"�VY���,�x.�۴C��	�AlhB=Q�ӡ���i:��Ez6�J�������|L{HM��w�~�J�MJuy���O�V꧊~h����=�[ː��L윙�՗ߝ��hpF�d��Z{�UPk+^����k����C��ZB�nS^�C��YO���_�?�2z���"��66sv�r�X�٭�kJ�Vz��c��|#uu	7&s�1"�o4����gs
��r�/)���Na�䔹1q�h�.�B���sp���~ʸY�ʟ�̙%����������> ZK��A�qIIz�e*�e-TRޜ�e�:_���-"R/�m2�x��3S-J^����'�̑π�{����!ȼ��q�mY�Z��_ٓ�]�ۉ�S�j&�g[~�B5��8)���C�I�W��#���~��c� j*�l��� �M�-K�ѵ��\ɜ�U�	3��k\�o�U�}�9!�'�_�|�e���q|I���c����+H������s�Q����:p�֪�Yu�=f��z��_rY�?hf�l %K�^����F3���@H�;���U��2��{YO<;�z�b��D��T�W�=��{6�A8��ס��e���\�.��ځp�D����lm9:�}R�`"v��X�<��	6�֗U`�g���#q�,�]Ŵ
�
2AX�`�	�E@�`I��h[(7!E{����* ���v8+���;M]Z)9i��1J�¢���Z%�q���$b���y���;�d������ʓdN�³O����qq��8�aI7'fR��T�~R��C�	�yO�-B�ZoDe�m3�c��<��y��2�#���jo�ƼJ;tcs��`g����^�ʥM�Ŏ�����E�n�J��g#�
=3`te��N�!�*�7vʠ")�<��hDO^���_ *�CB7e'�����Vy���%;0c6��&����H�a�DtE�O�A��}����xJ����6��[tc�Lf�����gO��3���G��6]in���m�m�q�V���`t��L�z��mģ��e#vt'��2@�Ѱ��@�S�W�>�(�/�s�-��� �U5
\jG�FE�� �/R>V�����T�߲s���
���G�7��a�Υ'L(����4,z4nӥ�>�\�Kk��X[�
 �G�!DC�Ba!/�|F�r��ٺBWH!�_�M��wB'�}�ϯ�`� �Xo��o�:L'tR���:	�q9��G}�1��^�25w���z��?��x$�c��[�; !���쨢�%�(J>d@����Rm�V*j�ٝ��6m�������������Zc�6�6���˒	�3z��c�dpD��)�@j�Z�v���[�B��_���G���p�w�&�_ݡ�Qi�_=��NGfF�X����Z���E+��������t����-���W�h�/�vX:�P��t uM|%�K��-}�HE`�0��y����J���TU�P�� d�"I�4�D���~뷥�7�"$�	톐�ZH�d�K6;�(�U�D��pF LPGX�e<,B�M��>S���V��-p�U�����jo@Vڞ�јP��qn�t�<���v��7t����"�o���XG�wN_������ݦ*�sQR%m�X@*JkҘ~. ]�_]+��f�x�,��-#���dR૪�w��'���F���ϻ�����K`�"5������U[0��K��Dm2���b��3�D$��o�mه_{�
<����'l/S�Q#��e�>E4O�~^��p��-�ty���=�ST+ҟ?�H�C"��d�p����ۓLF��,���ة��x|���E�ʄ,X�\�P���n�o��1�;k����KߣYT��[g.��T-�pH�=M��j�v��u�,M��:�0�G,�u'�7}��I���
��]� �L�Qڤk����� �r�����,�Zz�b:�~{wCyv����l��s\�����*x����dW��4T]��XlJ1V��dլ21`��N`�
��Wh����̊��l�^u:t��/�R�-�ZƂ�嬐�o�_�hdN�g���R)�`�����'�Ϥ%�8��f�}w2xd,,�C��hJ`��/���'>�S0[�P\)I}s�$؟�Sl���h
6�P� ���2���9� �N|K�_�ĩ����>�|ȩMfbF.a�A�D�]��|0���d�1��'�~������}2̡�R��:�־~(���T)��hK������ʵ�3Y���A��L����^��{�>��`4(���TQmV�)f�p����c����	�Jl���. e��k	��0ٚ�Į�M�:	[G�4����{ b��HYٻH{	�W�]k��t�Tb���O|ߖ��GZ�Wt����b"�d���'�A| �k5�Kg]t,�W;���p���I�Z�2�FwB|i��J �p��n�00[)��a�,-%q���b $R���㣃B0e�	��z5 �J<�gJ1�'��m1��a�������m��zlp��c�WC�����5��V6�f�*���|�x��fK��rA#�P��E���|6R����zyt$��b��)0�ڠVqGz�I�.�����y�F�&=QWUr�Q	ƲLN����VU���Ǵ�Ό���B��!���$4�� �$�^PË"v�GS�b|F�WB/���[e����A�s>�O�Ag�����=J�N�f�f�m�W����y;�=�t�ٴK�;t|�g�U��I6�����1j�
�hޣ!��Q�P�1�7�d��Ά|3:���J��PH-��QF����Vԭ��.-dS�%sQT�b�^����*���)�����FP~��p��F�)m���<�Jk�{�:���dќW���l �0�ƃu�]z�;�tV�#�Z�C���3���)}���WF��
�!h3�Bk��*��{@+�����9;�I�gP�`�A�wnޥ+[�`�G�63�D0F|ߏ�g�?�O��m�bgc��%ђP
о`�1�q��1~|����]��.��������ྙШ�J��b�����K�}����2�x"у�1u}���LDe0� l {����j�*���5se�5��U�u�q��I�Z��j֑D��@Pb�kͬg3Q\�
'&�z���Ed�m�����8����ˡd��ٗ����f�l }�J[mЄ���_Њ_R�'4K�;D�t	���#'N��l�
��#�O-T.�0��M�6��}n�A26�S�O�{�33�_>$������!;��v$�VZ_(���o�d;�Eb%ڑyC��P�����
�ll�s����";�,q��p�� ����S���%���D�MX��E"6�B���yN�}A�ӂhi�k�Bݦ듋n�M��+�T*F��}5h�~����g���&6Y�h�k`i���Ŋ���F[���)A��_�:���+Ta����\��@��Ӑm���]2�IH^���u�֝w��x u+��FS�7�\;��1���\@ε#���h�X�e��Y�BN���_�ZZ:��AV��Kۻ�_9�I7e�\V�MB���G{ ���du=����uG�����/�B�l��'<[آ���>���S�uW%�X�)�A�^�����u�;�#{����\8U��J���;�Ჱ��6�񳣆�c���68_.��}vzB���<�e�шZlJ��&Q˻�j���j�fQ!���e8�����Ŗ2�֞�i<���{Z7y�B�E3;�2֤N�qvˎ�����/����x����I�T���J�g�r�����Z�m�:�N��K� ���Q;��Z5iŵ�1��>*Ȧ�&������`����}Y*U�l�`濫�v3E��,�BҌ�����X����ts��hɆ�197G�
RƎ����c�m�--��u�7?�r�B���螻�0f��<�����%�飲S�k�h�^ٌ��{�X�o(k|�����[���$^������/N���Vz�y ���+�� ��>�ϲ��n����y�������V�g�5��Jl��Lߊw%I~����2���G�?Y*�-�vб^b �V\N !�sZXt���͘j�?��:�K��16�[�|_���G��Xx��@�6�15���M=^��c�'�񖊞UT��cm� �7Gt��2@DC�hM~�ZD�)cmB-���S�t�v:�����c�؉�j�d�Z@��(����)���T���ҹ� E-Eo$ s�}��;/ � FC����V.R�:c`A5�g��!�i��t@GɄ�y�{�#z�<�>��S�bPp���T�}�����3��dĎ�����_<��������W����*R�b1�=#��>����_?��ة���C��.ˢ�b�9}��1u����1��I<������e�'-�����.;��b*�����B�ƹ`D�`��|B��5z��_����R�N8�d������{�L�옝2�=A�g���aq�,M/�BbX�Y�(8'c��'��j�J/N_�����l�g͎��8�dHDnO벰N:�҈΂M z��c0M���@��=�(IL"S|�6�����'�Cz �%2.P-*z1��d܈���?�+� &�"My\а���Kzg�
�}�M���>�1"H<_@!D�ה���A�á��Z�Y:�(��A0�L�8��qDO�m��OŉE6��}B����c�/p.�;4�i��0bl�bCl#��C�ܯ��y�$�j�t������-��	;�P�D̷�L�R��tJ���1�N&�5�$�:�h<>�)%Dk�4Z͇�u���;�%�fPL%Rg�g�Ji(�(��Y�׿�{
P�X(P���d��:3~j���H�ˮ�kl�����qAId��1;����*<g@y`ŕK���S��4hT��3��w^�0P=�+���%��K���T«0�E�s�tc+�l6������1��l��6 Q��4�*����.�/��9�}�?�JW�EV�
C��y���y��o�6�&��?&S�ҹ�7!ȄgQD�T� ����Y	�Η���=*)_�m(��؞���U�-g5&<p�x*������x�vR*�q׶wh�P��g�R�;{�譽��=>�O>��NGm^�E�$#8!��d쳰s�t�S�	�A�D�1�b7�u�
F���_��T?�l�����_���2g3ۖsǒ�3(�6�M�kWuP�t!����<��w�D��q��l�9 �k�e��J�<!vۨ�@�{���=u���XB�u�5_$�7M�@��Iw�&Wδٯ�f ��4���n>O�������t�T��>�6)X�����T��Aq}E�
�3��8�
�0��F�v	2�b�3Rw�l"�6 �LK*IOS�z\�"SB��-��@����x�,���N�L�'{v��ST�S"�ie��!k���1�T��f��@�M��i)3�S�Sϭ}[~$�:�jE�)Jy^�u~^S�m�"IQ�N�Z��p�k#��?���b;�"�;�)Z���f��t�8Ǧ�_9G���/�.g=�a��8�� -�͓`�k�c	��ĥOf��� �k$�T[S[&�4H+���~f+<�H�v��ܒw�&�I�D�<���=�l�2 ����y��v{瀇��.'�l��E�H��á�5����/�'R1o�q�y�~R�����g���?�]��=��ٿ��ڍ�[�y�lHx�{K �?�4o���'�j��/�p2��욖����KO�����J��0���=Ah��v�a�E6�uQ_6]O��}M�ba�:U���,dSa,�г����2aH�3ȆIqc��-�7�p���,���
.��ie���4Wsp�ר7���v��H��Tзl���0����E?|�	u�LjU��)F�7�*�Wz��s�F5<{I_,^���M*|�l�R/��qO���p˼d�;>�ǏڴbB�����n=��8�Fl_�D'F�ħ��TBO=d�RA}Vg1���p<�#"�����8�=����c��^(��؅�N�g���tF��1������ڣ��[���RWFBUa������,�$;eo-ED&�o<�l�BM��3o(���,�}֩'�B"��c���%��sd� b1�E1��X�pOj'��vZ��6�-���@<��j6�fDe����� CY]H�3X*1 P��T$�Ր��M�^�p�է�a�wj�{��YWu@~^~�(Z� ����u彐h�Љ��t� >`������9�J��k98=�;7oѥ�:u�S���c8��l�#���M��*�i�H���}���.��
��e���]�e^ ̈́C���Dw�bI3b���� ��������1*|�
��7v�ioc��OO�_|N�|?P�%�?�rB$E��b�'<mzAf� kݕH9�m$�Ɗ���ʠ1��!��y�4�S�KF"���sG$�W'
��o�=wi:�H_��t�T��ھD�Y@(`(UUMl�Ȧ�܌��g�!�o���(�v�����7Qz���a�RY��0\/h�����J�1y}li����u ����{�KckT*M?�l!;[+u���ީ�(+T�U��x�m%��a��,/�=]���Ʋ���^�
�\�C&��/�!H�o{W�#�u\�KU����R$d��a�ŀ^��O��R")��tגy�97�9	�}c�쭺2�nqN���ۡ1=�@�`!m�y�K+,P�+�5赚".Q�|ƹ��������z<��嵳[�x��?������G�`�s~����|��������/�N�迾���֗7w��a����èU;˗l@��me��)4[ɍl8�����9dK����F&����tg�`�k�Z�����w�й����!�0"�V�E1@>��W���1$i�A��h�u�Z��b�%Gz/E���ZH"Xe�����h��T��Zo�'Df+Pq�4��,��[�9�>�O��� J��TH��wou��=ݞ�k�\[l��i���W#��}�<A������GX/�c�,w F0H��O�0h?M~ �2k.��Mm�_��j%yj�b�,��g�t��,�}�H�I�
n�m!���!��e�9e�x�f�ՠ����i7��yis����}n��i�$H&P�ؼ��%�3-`QU�hK5�Zu�����r��B@�U�м�+���X
m8����F"��i�l݆Q�2���J��"z����q5�qӪ��+/�v(2�ךF��=�P�I�S"&3�lϤǋ<ӺțW�t-$'��$�����j=Ly��]��}�+��ϑW��F!}�F܌��vm�N���N�Jc���Z��I0m�zd�%`LH,8 \L�ꆋx�Жh[�z+ď�<�uBh/���5pmsjD�S��v/Fr�}i�]r:����`G�1E7x�)-PN�Z1����qdވfJnF5�ֵ�'{Ů��	�L[�48Z�'�%�M� W�fTY�����~��Z搰�ⵢ���*�k�t1%�E=F���$����5"�7Pې]���pX����_�&Qĥ\__ځٶ�g��@!��欀�hnX����ۅ�.�PS �l!x_�h"�n*��s �-c�&}U�꭬���f�EM
�,�^5\A�I�	,�9� �	��J����*	�� 󙋂zPk;�ԛ�2燊t7�øsg?B\ᮎ�=�7^L �//�� |���g�S���9���
/g-�~�K��'�8]Vc�H7���:��A��\U�z���Z���kaދ"��n�g�^dȑ��͒�q�ݥ\�m�[���7�$gx��{CA������0�!U��m�'��	�9�Ge�^gX$  ��1�k<	@�����w��&q`���u�4܅�$��w9��%�����k�y^�T�r_?�(s��������	�~ɦ�.�/h4�<{b%��Nt A��4'r������e�j8�<���6�#)��&CARx���Q��<���0�_�3������o~Ԧ�T�X��g
�O���y�:��q��OR_�aqV�b�:��,^h%�Cm��}I�
�A��g�%.:��sx$ie����7��E���jyM~��L4��4��Nf��dhZ�|V�+3�F���Q$���	�ְ�Y\��hF!a�����b#�l�z«�����YY�2ԟDր�W�<��&u�ǔ�顝��F�@��Ý��z'Q�"��c�/�9�̰����V�l�K���3hc�k1�|��t�� �O^�W��,����Z�	����N���2�1!Y~-�v��<���k���-"����ߝܟ�7�W��_����Q��r���x熏����w��GQ/�y�UFe���dȚ=��{d<8(�tf1/�O^��v��ؑ��X��6�Ǟ�&���h[����V8�!���<����`����ϴ��3c�Y��s�z/��$�*��+�M۲�MWW+J���i�R�8ΉzrS�妿�rQ�zU�� �a�N+S6�Z0'������poؘ^;a��� r!7շq���)�G�2|=s� �8��3�L,��<��a�;7x#(�TA�r�� [�Z+�'piSWʋʆ���J ����$�{W����chEQ5��7���)����V�)��������!���c�����mH��ro"�$.lޒ`��p � j�L��jyw|�8�qڹa�y�8�9��,K�W�A	�9#77�Y�_�	^1S}?�X��umric䣨_Z�3��<>�u�-B�[�����Ŏ�	�<������Y��K�"۔T�Y�V�&\�&��ur䂹
��{��qy�>���W����n�f4G���G���� r�F�W�C�
���B�9-M����P3�8���2<F:�Ҏ�H*��Fؖ�~tU��
�)q���#d�j��>r�,)O�.=��(�Bs�Cǲ狯[th5*�h��_�0洎�;��Ӕ�kB�5E�90�#�uJ�/4����0'o��ѳX8��0���a۹���kl�(�
�֍,],�8�u@y���Y"ד���f��k̣��Z�^Ō]Y)��d .a�f�U���SOr���!5
.@N�*����X�	�AסU2�X}��Z.��ɟ��m�$Oj�l3��F��L\��_�Y�8G�&hm˵h�.�(<��Sw���Y��U	t��g ����ź,�"�γ��$���R��T�ڪP�<Z��p��`�"o���h�Q b�B�ypO�K�^g�C�6��
h�-֓�ջ��@�>9?W#t\�љke(m���5*Ip�7e��e�I�6#��]�qs�gժ�i8����V4�����o��~T���N�!�6���63i�JP��5O�/W+� [5?���oW�fb�X,��蓂���^}��2DAe�ߥ0���ڼ�P�ȋ@�P��Q=r=	v��ѹ�����*�)h�M^�
�;2q9K�x#K���1��׏oݟ���}0ܯv�$�w�
^���c�BB���y�,$�@�yMk��@�K䓨75��e��G�9{I�`i�����`�0��q+x��5uҼ8�@T&E��C���\�{��7����� �^�Q�Q�7��"H�9n�L��U�Q^��j����''Rd�`0T��U��a�B+7f���N����@�@6 ��Wx���V�|�t���#���Pe����ei~\�Jk�J���d�.���ħ���|��!�E�W!��ה p\����îʞ�B��ɇ"$.�\��U��fq �x�hP$;F��26� %#u��zD���{ �
�(�c^/r-�>�� �W���we���9$��V��49�fK2�$��@`e��~6�|5[�6�O ,c��'*y�qT,kn��2MSENp�@۳:� `q����*qr��Y�^�u�"������,�e˔fQ�?-g���ߔ���\e?��۲^.>�=�Gw
�A�fy��8��_��-��x��0:$d+� r'�L���Bh���-��E�d�iϥ�X���\U��x�aDA�	��k0�7�E�l$��'�&�
ē�j�0ŪA�-�1h�t �B��Z���r����/�E����y4�!m^�k֖��'�a�J�U�U�V�c#-O�F6��H/�Ο����yE=�jow	�5���[q���v�/�j�C1i0&���"Tֱ���&S���fG6��)��-:�^#QE�-� n
���B��?շ�zs�p�و8q&�)��%���ap�.j���5;��V�U��'���8�֩�Z�_ �2���X8���9s-"U�`a�~�l�"��ta������p89_d���Q�J�4a�?�o� �%���<��<s�6����0��I��;n;[
ʧw���,�-<��ܢXϑi �Z-K��h|ۛ��*{�x�ă�4z^ ���k���D���L�x��ƬF��E6���s���{� �E]�r��>��c��qa_#T�1�uE��k��u+V&Mټ�)��.C�}l�>	���g9Ce
ae�Ѓg3Ö=j*s+��̋�&�aU�*gҸ�eu{gi�-��N�c���h��������|��8��O��ݾ0ʜ��k8�|�0p쇈b�C���,���o���pT�y8Hܭ������-{���v�A��W��̥@��_ V��W�S�w�)�����#/eZxY}����Ͻu��<ἀ��	��釹��ޘ�隂۬���`�y?�S�Qئ�P��x�����(����� {�e�=6�T2[J��8afn�d�\�7�?W������}^oǩ�^��܀:���o��
n+˽�&�F��<B�žEu��[�Yg�ׁ���^5�ު��p��E5i6�,)��ŷ�s��X<N[Ltb9f%e@��=�I��E�D��I�D8�c� ��ϘX F��U�~EN�� �ױ�j� )�W3�&e�:o%s-T�k�ǀc/�)f}=�Aq�؈�5$�Y��0�0+I�]���,��J�gv��+����m"-�;�	`/����fȄ�e���`�G�3y�pZ/QO@���*
^�T�<�/����<`�QH攙ܧdP9��"D�D/XX�G�A�r����X� �)"��pC$� ���MN�1�QI�Q���,p�8�g��G�.k��e��T����?��y_=������z-�2T��ʃ�]�2?^C/�J2R	�h�
t���?H�� /�~��&�l�T��$i�*���� �$dDm�r��\�.�W�������KY��\��/?������Q��ܧ���#אѣ��L�y�,Y�=�>: Of��X��H3�,7��px�\5��#C�x5�g:�垱>hCub
t�e��(3���eXh�`E�D�؂T��eeGZe��s��cN��"N0�p|���D�-g68��BY���'�~RU)�i<ꅭ�AR�Nn �>�VB��1PDB����1"ǃVɨ�b�����ޑ���C"Q4�t�p7 ����wb8���߹��P(��#�L�G-қD�'"D�B�n֓�y�t6B�F��E:$�ג\1����V4Y�5N�vb6�_*Cs�HPa,	K�q�~�qY��W?��uS���vC9j
�x���Gu>��U�V�����	�w����Ҁ��Iǧ�2%((-l���ֽ���������*GP��^�S.8�6F:>iS)��8��`aU�}Hq9/��T��!�I�.�T�2�۴�����|x��Z׺����x�~�,#��]CǊB������;3����0T�#�J߀��My+���,lk�z�N�� L���̓�X������O��H��Q����5Y��P�S�2W�Y���p���x�r$��8�O��j��g���W������R��H�/�H�v��4�Q٤���Y�r���i��awC��'@w �fY?��iX�;Y�q�z��[�^w��tc�Q�������0d�;�?��i
z����5֥�Ky<��x�1�1FD�݉;��G�#~^���P��T�{W/�nk9~r,_L_��ͤ6��w���N�w\��ߺ�(�r(u��| �[2,aE����{��ǣ7��ƕ\����Ո鷪)m�ilЯ�0�����	ݲI��[sQ���yX��`�&eoW�I��H�����X+5�D,5R(���0��Vg,���������/]��<����z{�Ͻ��*�ڔ�o�ܨ��[�^�z�~)b�٢�Ϗ����|3��YeT������R_����7��;�y� �@J\�X�4e�Ȣ�G�Z�d0��V���TL�Ǔo�b5?�H��#h���JZ3�6����-fz	L����;�7�
i�Q�Fs߬F�Rf#`�\s`�K	���/�%e�]�2��)���q_k1� y���)3���x0���#@m^F� /?j�HÐf����NC�X��\rXs�I6� �\dJ.�(��	o(�T�`�-`y�d�A`�`Q�5�*al1�G˲sC
��%�^Pdq`&?�eEXUK�V'�Z��&�ʞ��(��7�Ќ�(�~��nA9~ �(�2��YMh��
"��Q�t�C� jv���eG�#�55��h���ir���\D���T��d�lX�s^g�� `��(���c�'����eM9����9�^��(��z.)Ÿ�@��E^5�����@B:�� Eq��ߍe���p{{�������S�B�y����s��?��=�� �
^	}Kϔ��8�	(���\��9�i�ů{!��S���湱��l�F��6e�-e��� 7�iҌ��P��(�@��~q������~��e��\,��4�D��#�*�eI2��,c:!f#�3`�'���`
b�hM<��^�#��N֠�r�7!T+��'�#�1� �&+Ęm.G�7����\a �f�Xy�G;54a|��@��e�䀷�қ���ȇ�ϴ��z�� ���ٕ�
�ê�f�a�xd,|0A�R�0�s�8>��M �~���>�JI�M�
э-^�9���ؐ�X�@V�rIN��yx�pr��'j�Ţ^�`��p".��U@�Y��M�����n��p��e�rZ�j3{G��`y����q[�<t�T�9�����1g��P�ZZȝ��g??��]�n:��<�a����4˅g.�Lp�pc�#w\�x���T=w�,��x{�3 �nB�)��<��[a�q��d�]�yئM�b�mQ��@��<?�!�<�X �?\έ/8<�u7O�ţ�K����rZ�q����a���ܗ��;9� �F����O�k.����E� ���kh�S��u�#��^&i��ի�il�cT�yx��MĆ:"�xT8 �\w;Z�;{��t����<�d����&��g%/3�#���#�6���ݰ����#��H@9�B�H6"����Pxk��DEr�Sҽ�����=y��D|s������J���g������>V�����GJ��|���߃,����\�k��BhJ�?����K�.]�t����!��B��$�5��ҥ�/KץK�.]�t�ҥK�.]��tBإK�.]�t�ҥK�.�T:!�ҥK�.]�t�ҥK�g*�v�ҥK�.]�t�ҥ�3�N�t�ҥK�.]�t���J'�]�t�ҥK�.]�t��L��.]�t�ҥK�.]�ty��	a�.]�t�ҥK�.]�<S鄰K�.]�t�ҥK�.]��tBإK�.]�t�ҥK�.�T:!�ҥK�.]�t�ҥK�g*�v�ҥK�.]�t�ҥ�3�N�t�ҥK�.]�t���J'�]�t�ҥK�.]�t��L�d���_PN    IEND�B`�PK
     mdZ��$�2  �2  /   images/e77f5de3-b891-4dea-bd4b-a791874bc34b.png�PNG

   IHDR   d   ,   ��U   	pHYs  �  ��+  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x='adobe:ns:meta/'>
        <rdf:RDF xmlns:rdf='http://www.w3.org/1999/02/22-rdf-syntax-ns#'>

        <rdf:Description rdf:about=''
        xmlns:dc='http://purl.org/dc/elements/1.1/'>
        <dc:title>
        <rdf:Alt>
        <rdf:li xml:lang='x-default'>Untitled design - 1</rdf:li>
        </rdf:Alt>
        </dc:title>
        </rdf:Description>

        <rdf:Description rdf:about=''
        xmlns:Attrib='http://ns.attribution.com/ads/1.0/'>
        <Attrib:Ads>
        <rdf:Seq>
        <rdf:li rdf:parseType='Resource'>
        <Attrib:Created>2024-06-09</Attrib:Created>
        <Attrib:ExtId>a83a9794-4a4d-4c22-8a84-66c76feccbc8</Attrib:ExtId>
        <Attrib:FbId>525265914179580</Attrib:FbId>
        <Attrib:TouchType>2</Attrib:TouchType>
        </rdf:li>
        </rdf:Seq>
        </Attrib:Ads>
        </rdf:Description>

        <rdf:Description rdf:about=''
        xmlns:pdf='http://ns.adobe.com/pdf/1.3/'>
        <pdf:Author>Firman Abdillah</pdf:Author>
        </rdf:Description>

        <rdf:Description rdf:about=''
        xmlns:xmp='http://ns.adobe.com/xap/1.0/'>
        <xmp:CreatorTool>Canva (Renderer)</xmp:CreatorTool>
        </rdf:Description>
        
        </rdf:RDF>
        </x:xmpmeta>!��  -�IDATx�u|g�\�y�y�s���3`�X��.6rWZ�%�D��%ْ��UVp�U���!��*˥*�lKeI)��(R�H�\r�؈],�0�ɩ{�s�~���׃�{k0=���;���~sc?p6�"D��^υ�� ? <��.�+ B�)ݐ�M�������T���E�4=�E����IO<wh����`r���+����^��ˑ9.���#>�|�CUU�ÿ0�&�m5�˹��QC������._2�5�|�6�(|O��N:T(���c�bVG\+�Bh�K3�y=]��kb~�cD�J��jȹ+�¿!��|UXÉ�r>
?gp���G�kEA�DiV9i�`�V� ;�����lm �`wh�69�x�&/�m>�q�#���o�A��y%GA�����,{���<e�H(�W|��4-:َ��?����,#
.��v� z�+!��9Pa0�jk�%UE�uzxm�R�p�n�)%e(_TTO�NL!m����������jz�c�"h�@L-r���#��JRO*��(5T�У�#%��I�BNI(��ӸbH:E�:��,*�b���n��C����x�#���KJiZ䅾�iE�t��k��?���k�l%�����o��=�uՔO7�J0H#�p���g�<~�U�l(!��i)�?�F"!�FUz*�)�-������Ӓ��ص�\%��Ⅱ���._QB�E�5�+iN�0��y��8?P���<y�Q�B���-e��R��7�J����d��w��`&�O�u���B:�/���]�8z7
#O�\y�@L;
U/����1��pa.��멊������9�"�C�#���L%�'�E����j���` 憮��ux#�W�D����<d��7��G�%k��U��8C
��Wǘ�g�F�0
L3;$$0�4�A�/m����	Brrj�K�hg�]0J�F-�.g�@f��a���K��i|:%�|}��2��!��vu���{c�#�����s�B6�C����d
O'1�.�y�+[���u���ώ���2g��b��uS�>�@�\�+�1�k���._h� R%,���m*���"�/���봼�]E��.'�i�F�++֯|��+�3����w����؈�^��_��ԏ�����l�~ٵ�jwڇ��������a�n�t�I,M�I���Q�,\��#aŏB�<��k!�=����X��&K����5tB��qB�Q(��j�ҽ�94�n"ed��b��asm	�fE4�8~���8<6��݃�H�R� a��̧?����ׯ^�G��� j��%���i�>����H���&�@�M��}��q����4F�)�D"�}���D�~3RYW��'�k:�_�mu�l1�cJ��:������ �A����?���f����!�|}�	}�f��\|%h⋵�0�.�b6����փnY���@WS��|����ip�rd�G�S�e9��a[�Ik	i�FI����F=K�Y�����2'��Wp�j �H����k�e���Mu����w��=�N'N�Dy��͍u�����S�ݕ���41T�o]�%�xI2�4�g��7��>�+���=�~v)��;d�� as�~��f���2|�qm�F��/��*
�*2E��z~��?�o���3cM��X�����Qx��;����7���Џ$~{����a=d�E�Lg@�0�,�M�E�eTuY���\�'.0T`�`le-���2�i/o�����ӹMl@'��r�'������%jP��X�<6{ӓ�����-��q�2�I�r�,����}MOOcphvφE�*
\�F�u�̙����ī+��ӳ��$����Q)2��G^���%	kQ�����F8��P��`Px���M���d%3m���s���������?��P����c+�ՃPq7���̞��dO�#CO%~�>��{�s<�#fHĊ�跛;X��#H2�h��eJ�ȒI�G�'�0���?k���r�����rX��B"b ӣ�Z���dYih�%����M��� 3��W��3x��g��[E��E��E2���qi�.6�WQ���
~곟��0Q��?���<���I0����N5�r(�;v��Y��ge4+�I8Nv����t�,���ƽ�Z&��1<:u�,���n�� f��X�.�'�h�����r��B�_�5���g�{�<2�65G��~c3���vm���`0;T:c�<��#Xkՠ�˽���:�¢@q�?V�Ę��sS�'�a��{m�dz>Z�*�
�������5�^��Y��X:�p�a�_��Np	��H��L���ܳ��������)�F��A���#��;=3-��1�B�������Hߪ��(at��c] t��ƔU�e�Vd��(Q��)qָ�`\
R�fQl�n��?�6q��ka�X�TyY��kw�Di�0ΌM��Z�� �L>7L��/DP��2��tR� $4y�:�su����GҌ0n%q�8��T5��z8�X#�r8��c��E��碻u.�$�*Z#R�,��oͣJǊh�2j%���6+4(a�4hvU<u�f�t�!�&�ݹ���4G	?:��t���*b��t"�.Pwv�$׮�7�	c�t���Q߰�b����Tc���B�(���{�t������V��mZ����V5��u̯]�V[�Ev*`�P.3���*�NGPc�L�&�"C#	I
���!��Ay���6.���5@F�����8Nn��s�0��D���&�ڸ��f��R��)��j�$ Ȑm�6!$��t{����nr�Zm��Bi��,�Lo��`����Z	-�*Y���9��w��mbjx3̄�7�#I'����x��G	C�̄J��B�󃋗�sd-�~qW�o��]�݌"����� �P�һ,���"أ"��'�|���Ls�
�W߀!:c���K�hP�n��(����8,mv���Cn0�fm�Wq��@ Y���"})YX�<h��1ce������e���tX�C�s�8�.�R�?��0���(��)�Wgv��i���Q	0FG��
X&Xo8y*֧����F���[��+H]t֘Q���{�\Y�9�\e��9>����^�SO?E���d�~�㟠c,	C�|�������ŷ0��I��c�dk'�kT���4�e81��:*�E4ru�_���C��P�x�q��C��1Cm�����ǆg�Ԯ���cu(z5N36>)[e��2?�B�0����!�8p��'2CLy#�o5H����|���m��;zZo�z���c����)��.�9F����rS)3��EW�{8���YG/K����]�Ӄ3$&=4����,uE�)���DF�:7����6^|�e<Bx������$k�'�Wۻ�����������C2�5:Bc&�$�	���>�
Q����˾��X�����&G̺$���;�V�Gf!/A�r6�i�}�C�h�(\[Hj�fP�|�
����W?�'wN �����-M"��,O���n\h���%��fPJY���kF�y���*v�Ԝi�椳��(�.oX2�߱+x�����m|��ne�~߹y�B?r��5���箾���Q.�QQcTUl�@���T6�B�H���/`e���������߸�����H�u�hm`tp�Y`�@`�$-?fS�q<f^�QT�&�pPܑ�]���!�hl���1���xG��r��I���U�j�@�|s��Do%�N��I�+$IA�uyى����S����Nࢠ�*�k��Q�����x��Q?�4������C'a=�M*�K�U�r�t?5xy
����O:��y�5t��Xq��LAd��{�m*g�}7����#pR��G��l��MR�����V;]CT1�`
�k�(�I$Ho��6�n4���7ajdc��#��2���*�q�Ye��Y(��4H>��~��E*��t�]"��#����1	:�E�����QL��0�U���^���dI���Q�(]P�0^���%B�d��'�Ǹ@6�xIz��A���
#wW��yq����C�Y��S^BF���[a�DFé,r����,͕Q-N#Oj�J�}m{aӖ(��&����$�J�F���2zUoN3��#����k�7���ۯ���g�Is�K�j�qx���&�ޗ�}B!۔�;����@�ل�5.��d�^�@e�G@�/
c�t�*!SQ�;�VUhsjû[�Zm�Mbgy�Ȑ �$q��}]Bg�J,r�g�Ϭ�D]���Aw|��?�ה)#�}�J!�J�Ɋ�l�������نk%�HyǓ�%z��Ţ��GR���釘��8�"|�X�ѯ����gJe�<%)���>��L{]l5:����g��b���[dl�FdS�CE:���G���5q���HsnS��O�y�L#�d\s�1���p:C�!UO�xa~����I�����/(�l��B/����<4G|^�bL�_z"OB�㒞
�����
���'����)L�hDD�7^��  (�/@�塹�%K͠��`sޥ�z��}S���DI������2}J��G�cXu�X�G�gQ��c|p�]�nTt�� Y2�IF�`l�GC�Ɂ�!y=��EJ��c ]J�zc)�f02q�K;�;� \����.>=s��^��ׯ���$q7���E<��F�ϱEцH ]B�(�ɂ�RuK��UUt4x>K�ȌP��"�E	��}�+�Z��q��� �Y'J����n��~Ch3S��m��UU�U�8��/��s�>� 6o4Zd�WP�CO��MC#S25EV���o4��i��^�YÛm2�b
�ؼ����s'h�oVW��Z�7�i��_=�s���>��+S=���� ��˨�C4Y����h	)FkuX���F!�Ǻ����>޹y��dY���X5vQ�pq�YB��ک�AF��&���!�X�@[�C�$�v�o��"�c�!� T�;A쯩���0sT��Ş�pj���o04;���1��o�P\�Z�r�Ua���Z��4���~�ݵ1>2��ު��DJH$�%�h�13�y*0o�����=�L�I���dEF�z��%�~�El���n�ё���P����R�~�[�-%����U8I�6fT�̲� �,���M,l���lÎ�K7�v���E�g8MB����<߸�R����	�	2�B
�Li�B���vy���}I}��2����!���]��.A�������m�%��(Q+e �N��z��	m
����2X�E�G�{8�\��:��a@�R���O ���:�k�)�L��~��y|gw	��ć�2u��� y*f��8�/�>�Je��ܠ�h�P8B�A��5C29�)��s�9�c�����?�,��u�;��$Q����P%=e¥�2D���E�_tX*\���Hfa���-�����Gb��޶�(�"��X'�X�M��_����z�����h�'=	9G���q�l�jz�[h�=� �U�Ǌ0,M�萬�x(Gہ�������_�g(���l�������B�_��@���f\۴�e��|��k����W�00��� � ��2�>�hч=�@�ۯ޽��e��F�+X���{���f����4�j �1�cKc�uFR�F�p�,�'�d[6\��q�Ϊh����θ��-r��Fy$�T�����(���^a�(޳x��»��R�xOEԢ<-��xg}��RG��N"�B����s�l:fW���^��G>o�����6Y�@{�\Z�
���F
�R(�3�TO�ͥ��@nY#)F� #�+T����e��W�qj��$�Y�J�wO�<���7��;o`@��"n���L4� J���0�LH�������t�ڢ2w��2�������Mf��]�y:m����tO��7��Ȣ�5�����K���~�V�3��T�z�{t$�l0&D���X�-U��E�`�P�αy�N��E�4v��ع�
�N�k�-k�>�	G�Ҩ7�&(2Iy	�M�����Lz�ө�?��f/�vpvh'萧��$�.��ƉJ�� ܀QaH�QbԎ$h<
��R	����%�T�^�AJKc����4d���~��E<G�	$�0�`Dz,�"��6<*b{��}͆Q����xI:�?O�(���/j�l
խ:#��5�~`?���QãP�,�j?������6I@R�T�8�����*�aQ{�c��t���9���lN7U�*]�qh{���'lLN���� <����D}���urL�Fq�c���Ù1�{��2�E����#G��>��_œ:�tʔ�)H�>5=m����ܩTq�(#_�k+��o���.�z�#���~V�:ov)2W9_�f���l�٢}OD��X:�aM�N��!Zd���է�aIbC�W��ɕN9�kߋ�~�A�S�v1����Rm�@}��kb��+Ȗ�fЂP�NDӰ���b� 	�<�US0<\B*̖�qe�UD���G�������Z|�`_��·wW�k���
�����ad�nu���V�_{�꜌JvT��d�@�8�aI ��=~g}��k�nu����.5��qe��O������oB�E�$�3E�.�7BK8��\8E��V��/NT��E(�C�� �4���p��d(_���@B�@Fg�F_�~�v=���ŢR���n��@���A+2KL�:���ė���ϝH�&�i��)��D&�@��@�j��$��c��$�����h|���,2�A-)O�CKk��>����.�`����R�t��Ǆ��lI4 �Tq2������,r����>:����S�YȘ��e��,RU�P�R4#�_0��0�D���`��k�u�)C���J֣q~���Xe}��n_�\�}���3��ۧ��4�3�!�[D��W�=b��Њ�o��(L��#�O���P�N�΢~��7��j��Cih�&�~5�|������m)��F$]:ר�<�KX�K���W_,�0X�/|��>6s
��W�M��$�S,�=.v�<��tȏN?���u�}|^I2W�7b�@�����d�_�̚$����u}�8���Ds�?����r�G��vz0�4а	'c2�T		Q()K�*�oe�|�L.��.��řq .�PU����v��{!�[�ã������z^��R���w:.*-�O=$�;Κi�w�J�Y���0\�,�c�'-��ޣ���,'P2H��h��a��btdZRAU2�x2�8E��on�����!d�iu�4۸�!��McQ��R��y��Jͯ�4�<�$`���Ǵ�<*��n����
�����=*�.R� %-�-9�j���yF�ьT����{f�jS��!i5W�Y�%���=,R�)+)������}På��,�>��{D�=.��V�qac��J)4���I(�GQ����=��I������.�>��pRv���M�B��t��Q��;$��T�>�RcEZ�v���]N˵elu�(D#��(���`�}i�2��a�/��f�5j�cv�}�}R�?z�9���x2�&3�ˣ���=y��e<_ۄ��d�N�8�\fB�B�N�WF��Y�8b��$JJG��"�Mj�4��ɍYM%I��H_�}A�Q �-Y���D���@�.�w����=&Nkb��i��?�diC%#��޹+������q��{�Md�4}�;K��`f��t��4����@�t*a�6�]�e��#�5��j�
��:iI9�Hf2˽؛�֍�M`2Y F��7>��\{	�n_��Cf2���я��L�)N�����]>�3�G1[�;ﬣ1I�sT��S���}n"�Z@��'$��Na���Ź(ΙƷ�8�<��P�b��n�i�V�oF�l0
j�"�om&}�C4J�y�@(y_�ms�p���j��mbc�����6Z�E�'��d�1jp��tF�B��zu��6f�O@���ޥ)'��K�v�hy
�'���8Fu.J��Y�uL���#	0��W*�{�*Fx�CfR���(H��i�(������u�T#	7����8�������M|���!Ɉۮב͡}�Y2��˳�
6uz0�MB��5�x'U �p�0���u�{=��4�����y �˗Y�d�V�'�o��QU��C4-�9sjA]�.�^B�Fc�$'�ѭ�392Cۆ�qD�Lf�K�^SÇ�2[819�+,����7"'z���c��Lٔj�b���j,���$ɏ`��A��r9|�G��"�*Na��l᭷����D���O���qְ�x���)e&��YL�bM��\��!_�"�,�Wv���*�`?:t����^�F��j��Iږ4�FW&ņ�)���{8�#T�R�I)�[:��J�!��Jǫ��@���}0�*���P�]S���a�$��4_���M���$d�	�!)/�MH�`5�&�2t����cU���H~[0�7[�iO!$b������F�� �P��SN$Oܥi�f���i�V��X�Zv���φ���l����s[�
��W���kx�N�R_Ü1�4)��Vv*ȓ��mBV�|E��g~�\
����a��f`g��[Cؼ�h����5f	��ߢ�̢Jf�Aj��2�~���^+x��+ Ol���?A�!hCy�F�������5%�7b)�Hvd����ZGy0��F�C"Bh�Ʌ�4��)4���Q���&��^C�d���B��K4�Bo9U�x@J:��`�m������$��@X��.C#��V���Bc6���cX��W�MLf�����l�l���� �S���AH)8����\޸��|��&�<��4�v���<�NT�r�����������O!wn �|��פ�|�'$n$*>��s��Z���ϐf�P�n�ߒ�����[�Z�2!O�FRS��\�l.
�)I@W�㩁f�ݵ��󺊟$D�9*N+9��	�uk�TC#e�NC2)��i)�[�
2
2qrӧCD��d2e�� ���V	O
N�:O����#g��,�J��q���-Y�fF�X�pD����A��oE=y�^g����'Ҕ׸ګb�ك�w��g��h�|�L�Dm���Ç��H#w%y���2�D�#wK0+�4��FKr����>�^���9���tF�������s��C4`�����(�Ӈ�iŧK����������O���a]��8���Ӷ1@v7R*3 �����5{S�r�$%y�7e�P���%-at�sD��i00�0�O��Ҵ��7>�	N����uk��#n��ҳgY�F]QW��Y+����g��mFK�<��S7�"",;�L��m�����Z�:;��MlըC�?��O��W_���,�����x��>~�Q��}�`�Q�Yd��`���Pr*�N��{j��h�İ8Q��6Gԇ�8���>>^�. ������ޱ����0�V�1@���z�B���
Un��im�����F{�m��:����C���@2S���/�&��	Y
���������>�e�����ܺ�?n+�)�HIq(���{W$����a�HK0.1�_��A�K(�kL'�=�WŤsΐ�%	i8,�]�)$Cێ��,�P�Vhիة�⟮��ݥE�h�z��s��RW�3����:qc�V�A�fN�Uk�c�"��(�vk��!���Ū4<�/W��K�EF���߰S���~�U�"ʄ��Ei|��!tx�m��YR`
?������1�(b�5Z�XJtܵ��s�n�b���l��͝����6�f=�6���.��� �a��OiC���g�M���lR�h��9)M�>O􄴃è�������B������	X,�'R�h�u����xB�A����{�sq��e$������~3
#j[s����8��D�Lh�EQEJm˓Q����c�F"�9	+�Bq[��!LW<�7�H��i�"��q8�bg���q�W��]%fD�����}1Q�����.�F�c� ���ap��i�i�q$7�G�P��%,+���ɥG�Ww���џ�򏿶�ˏ\�6Ԥ���M%1�1F�.���ȆD2 _�e�N8�7K*��Ė�5Z�i˨�����&�1��&u�L���
z�fD��m��8꠾_ų�'1@u{��+�t����_�l���Q�c38�Qk���?���!N.�N2�r�(��ݷ��Y��8^o-�HfP�jm2�L�(����t �.ܥ�F��zި�0Uě�K�H��O=��@	��/0��z��8��<��{[(�G4鐰hF��ߑlEI �5p�Z�ׯ�-ĝ�a۷H X7<:T�hV7���>�YL'F=Út2����@t���_���$K�u#��p�>����7|�����aO����)^�Gx��%%Α����6�����''�U3���K�b��$G��E�>�Se������n��qt���eܴ[��l��n9!�?[��Ì���*�g�fP����<��;�+	���wz.=�#�5�Vs���"�v:0���X_�_�:� V�V�KK0	��������.��M����U�P��F���u��z�5�n�^߮oc�㉦�H�t�N�'�1I2.��$|��,��!$X�<��߰�?N�~u=t���_]5z��	�=Uɮ��'��Wę��D�'��,_wj5m�r�v�q�V)YNʄ+��w��+'�O��G�d�$��t��`��~�5d�©MH���C�<��u�j�
�\"�NR��>��N��QHg��
���X�9=2Sej�4��;�s�����5�fY?�X�kP���~t׭DfF�tHF/���l**d�]�o�Ve��Dv֊:�}ꉨۮF��Fz�u��ɣ�Rm+��H��*hz8`��%�8s��S[�l��y��9�h����HO	4Q4)Ɨy:�D_K��W�{zF5�:$V�&�,x�����X�� T*��(�HC��Od���}�o��š�w���T3*�`�ʮߎ�)p��z�q� N�G���He�H(�*#�\�����B����G��b(G
C���i�©�@�3͠�:4V�L�F�(����U�(R#��:�.�w;�h�n��甹�r���a��w��oF�*9� Fx�N�{~�a4�2C1������������L��&§͔�#�f�Ԅ���ah��Bj83̶L:-Ŋ�)��>
U��4�|ώ�V��'�k\��u_wIgԌo��Ө��n;�ޔ[�=�Z��oqd�7!nB
���V�8!"w�žw����_�����F$�e�G���xBd�@���B黲_$nG��l���|�'��}��P��.w��N n��c�o�lz�<�&OF��)QY�54��.I�x��<���CdL��*�+�JQ��qR�l���j��cJ�򋖋/w&Ŧ�hj&1B��kKB��m�ē�@(�[$�Eq�9ݳ�6l^��ɚ?�GB    IEND�B`�PK
     mdZ	C�@�v �v /   images/e975526f-cfd2-4a7e-88b6-747cffbdf2da.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  ��IDATx��	�]u}�}�]�ΒI&;	Y�$l�`�F� Z�B�Zk�hťj�U��>j_h�ԥ},տVZкP6ً��k!$d�d2Kf�����{��~�d"�v:B�~|]����N8����E���p8��pBw8��(����p8G�����8
���p8�Q 't���p8�8�;��q�	��p8�� N����ppBw8��(����p8G�����8
���p8�Q 't���p8�8�;��q�	��p8�� N����ppBw8��(����p8G�����8
���p8�Q 't���p8�8�;��q�	��p8�� N����ppBw8�F�V�qT��6f��T�8�F��	't�c�̇��޽{��v���޽�3�����oԧ>-���پ��Bkkk6����l����U����G�O��;gΜmg�qƮe˖�	�^y��zzzN��;�o�>��/l۷o�1a~�J���*�B�`���9�җ�t$��Ϛ5kdƌ#˗/����,Y�����o�����E'�����%^�馛�y�������r�]w�x���Y�|��\.��144�H�=�g!g!�d>��~g�	�U��bY?*�ё����)�����o�.\j`"���׾���~���:okiiY>ӊŢ����aNQ�[��O ��R���m�6�;t�m���{����gg��c�=���;��~�����1t�)��X�b$r8Ok8�;�q���]ظq�u�֭��{��s�9�www�ķ2圶�@~�"���Ig��2�E��8$͜93��NI6�x�=!ܠ��h��gϞ�?��OG��?�f��|�ӟ>)h���¥sA�µ�����������?��0n�����7::�|aB�T�9��޺u�Ж-[�����ypѢE_��W?�x���N?��-g�yf�i��6�+F��i't�Q���94�λ�{VД�B[�cǎ��d� ��@���|.|���3"f}D�"n����p���]��}��I�V�iӢ�;w�l���E�z�G��枌(��\sͪ0�&D�t]]O����55�A�y�x�Ms�-�!�½��1#�;?h�a���aܗmڴ�@�l�����o<�~y�%�<|���q���M��SN莣�X[��N���>v�-�ܲ*�Ya�I��ͷk���m��Z)�"Ai�"L�y�0�e�L<�ly�8)���z:W�:G�����s���'����a��_5�{e߾}���fhҺ�ѵ$,`j׷�\���:F��:Os�Gs�>���膃��_����a=f�s��ߣaM.�>���7���A����ի���+8��e���SN莣
�ز�ׯ�y���{��^������O	$�d�ܹ����e�G��xƌ��Zd'�7�."D����]�Lۂ���lr׾����85�H5����y�-Ov?�я�Y/�j\�O�4s�E�i>��Z�8p 9^��v́y���'���@��8l/�{/��g�����ܻw�+��<����䗁����X�������=���0~9r8O	8�;���I=h���֭[�������|~ض&���@��w��Q$���Xi�"��5'Ĩ��[D(��>��ȱ��7ڵkWr.fu�f�ٳg'��w��E�:F���tuuM߽{�����R)���L6Aa(̭-�e�_G���'ג&�o]���z���ߚ�,:F�.!F�A�O"����c}�f� S��1;��,k�f�����]v٣W\qŝ��o��W���N:�{�ڵC������	��R�~�_�������?���϶m�^4k֬ŁLj��dCR"3��4mm�-\�0�'�}�'��1�&�	H�<��E�"�={�$�@�V�\�Вu^8.���=o˖-3ü�+�,}?W^ye6�m�w��U�bii ��H�>N"h0��o�äN���[�&�߱cG��.���5o��t,����&���lv��UA�yI��7���n]�fͶ/�P����������ii�;w�lSp�����5?��O^�=/h�����gu�',��TD�B���4����_\D'�U�V��K�|F���?�c������"U]C�w��w�Ϝ9sVξꪫ�x���3fd㡰��Sl����1��{�w�ϟ�$���w�o�X,'6����[ ��}��6�R7�'��]��9k��w���}�SwE�r[������1����෿������;������y����Hy�c����x�C~q���g?[��7�y�֭[��=;��IA;\�b/�K�$(��H�����?h��~Y�Ej���`��!��ڧ�E�C>t4���3a�9�ׯ�h���g�V
[{>�i+��T�X�(gF������9�}�|/���m�щ�'�M��ߚ+���.�o�E@�a��uo���
<����0֙A�z�ƍ�<���׼�5��=��'���w�g�p8�'t�S��/��ҹ\p��(�Heuض2���-��4�X$D��k�(,>lA�EN�i�և�1������=�o)B �o��mD��^,Jj���85��p~����t��Ҧ��L�F�s5Wi�:��^h�)���v��ah�6 r�X���k�xy�Z�z���"�]n�\X�N��>}����7�߿{�w�s���t�W\}�e�=��7��`�p8�W���x�AD���|e�����6m���D��e����;!����x���	��Υ�o.(Č��֍�+�\���4������'E���l`���:v�����2�ׯ-{w����p��֫ 5��B5��_�.���7�[�׹�[
�p]�s�������[��7�=��f_'��M۫����}ױR8��c8�#���l^��}�G�x�+����A�s8&N莧d^��?��c����Q �f͚u�4�@*Jfm���Dd#���퐯�>ti�-�Y�2 15�-3f�M���� �m��o���� 5��k~���������[�+ h�Z�=�b8�<�Y�5W[]N�䷣�k^v���G�gN�NZBV�;^�hQN��a�3��w�w�������|�_���}o_�p8&N莧�6^x�^p�w��@�^�p��4Q}��j�w�ކ�Wd"�$���� ;�nFA�	�\��:�M��Hp����T5W�����4������3�����NJ�y���ڸ>�>d
�\���龵Z�z��F�<���1�cz�fyH^����#!g߾}ɵ�]q	ܫ��� �8��Z�x��m�v��>��U�\r�W>�я>�u�cr���xJ��o���׿��͛7`�ʕg�P�t"�iB"y��R�a^Ƥͱ���j���Q� ��+���YǬ�k�oL�"c'��9�V��	��b�� V���l�.0d����X�� u�O�%3o]K�j%lu���CkC���G�����X?�������\���N�������p��.���8_�m���N�_;n��֙�~�����]�{�@YȲ�gmhϘĩt�F	)	h�h�h��)h�����N����-�J�|�ܘ@3k��6�گ:��IK#�s=���HS#�{�~��%��Hx��}�?�ԏ��irG#'�^�;��Ӯ
m�P���/�Z�a��9\��o|c��?���|�������N�_+�m����׽�����(���@Y�K��T�L�o�ةc.X"��b����N*� q�?V�eV�uS�=M����sm��rYB�L�$%�P�7�wM_j�m�	A�{�į�3�?�hu�Hy�t��Z4?��A�63 ���ۀB���"6
|s�~�ο��nc}-�7r8�m8�;~mP�W���?��CZ�x�ʾ��&v��4S�H��e5C��W�5��@# '4Hr�����~*���C�D�[��@T8��f-�̹/�!�M��R�v+'�5y�����0ZK��m�|�̇`<ƭ�UOL�\��/4sȑ��s<in��P��3�܅A�{g��Go���K�;����p�������@�G>�e��z�;�/_~booovѢEI@�HH�"r�L,�NAb���&%6o�߂՚m�yז�!qr�m�v��ncr��)�b��l��u4�b�&XX��Hs���Q���gK�jL|��#Q����F��mW%h@ܸ7,!��~���a�C�����s�1�������~�nݺ�^]�����	��k��_�u饗�q�������Pd�>�3.2ЋR��w��&H�d���	��� ���[���IC��0��Ō)�b�H��=��V���lK�����G:�+9ߔjmo�Ց'��딧��(�+���P`	!�\�d�ڣ������� ���;ϳ��!`!�y�o���%�s�}����뮻nO8����p1��S��Bϼ��/<#�Ņ�ϙ�V�lٲF�u��m𛠗?Aph�6���Ar���5i��Hw|���m�������3�Aa�!P�k� >��A���k�%tԶ�&r�e�|�5+�`c��D$���U�ڱ�pH{�|�ߴ���B	Y�Ȗ�e���i#�w��]���ϯ1�3o��}햍7n���Ǒ�	�1������ׯ���s�/'y�~�E��]̻h�h���!(�j�6��i�,���O$��y�G��o5kKxҮ��o��>�Є!HHXc���6�|i�D�Sڕ�=��l�<~n��D��.��x��)��P�q����K@���7�����q�0DnS�N�c���^x��_��9�#��cJ!�|�ڵk�fzn�@[E��Fj�S/F�9	y�5�E;G�p�ͮcEF��5�s<��d~&M?dM6�����@�̑���#?��X���ky��õ�0��q�bT���Vn�Ρ�[�&������!׽�[�:�!wR�[B�賎���!L�4W�U����a.g�v�m�׭[w����#��cJq�׶m޼�ܶ�v����ac�f;�WҲ z�	A ��smAk�G�&�˞#�I��p��dR�0U#4�zl��h����}	��-����F�D��#. L��s�-?���j�"j*�铎I���6�cޗ ĳ �����Za�q��袳ÿ��|衇~~�D�c�pBwL)��������q�u����Q�C52ҟ�	�Ӡ��de����Y_�5��:"J�v޼y�x
>�_�Y�A@0���~�P��[b�Q�2Z.>f�]4�.dc�`�,1�#؀t;'�Kwfc�-i����A��ö���n���µ�6v��7߼(rBw8�N�)���g�}���3g.����$��j�����A(�G7�g��)[�j�
�#N�����8K�V��� j�!|@fV���s6^��PY�[cI��@�8+��h~�!���B�+��bQY�k!HpM��ڬ�0��D�T�w���{l�����pLN�)�M7�Բm۶Ӻ��:<FC�%os������*@bh�h��p��&qK������"(4{����q��_�(|���A�+�,��B$� �#�X��޿�g�(sޖ�M���V{��nl��<�������F������^��7o˖-�o����y�W�Ǆ���2<����4���K�k��tA ;_N: ͦ��s�C�T��O٦�!p.h:�c��v�g}�6u�8s�T��_��&P���\'�x�"M�qu��摳6�MDMљ���}��<.��Z�s��pݶp��{����pLN�)��?�Y���J���V�P����"*�!L�˚}�>u����Ai��-Pi��9"�&te_ #!�a��=����Q3o|�:m���m������6j\ � �Ĥι�5�c��fr�% �޿5�c���X�q(rc����Ρ4/Q����\8g�}���,"�p8�N�)î]{��]��Q��K�s���l ��� ���/n�� E�.U��AM�:��ӂd�K8�z��>[G]��?���V�)�mǼo�~�~�Q�V� �=�& �0>V
�ɚ��k�����k�x#�z�t�S�!��k,H>>�º8�;G 'tǔa���i��m�Q�47�r-c*��qBl�peM�߶x���4nS��ʦ؊�������k]2��eL�%�=�>�v�� �"Ў�j�ͩ�o���F_uK����ɺ��`)ptCc��6���,s��9�\j�cy�Ei���@�"��!���&̋u�>��'Ɵ��ӓ�Ǆ��2��[FK��l�uL4f[4K���v:^z�j���.b��m>6Z6�g� �9�@�$�Z]� 1[�����i��oX" ~�[@��j!s"����R�DoS�l4��_[$K�;Z��);kc�sn�kz��9��r��}NuH\���a<Oz�t�cpBwL	�b~�K^�Z.��;�Vnl�%m|�4����Adh�T�o��;�ϧ!0�Q��F�CP��!w�%���\n�͘���toS�8_kA}vk��<�Qs/8�	�Y��b-��M��o{_��%(k���U�P�[����'�����8��j%^عF�Ti$�ܛEWlp�%뇶� Z(�g�������(�t�8���J:��h�6����k��<��Y�;sl�6�B*��0y��_o���Q�&� ��>:�>}�D.�� �V~c|K�v�_$g���6� ��N�>Z�Z�p8�N�)C�Z�Gq5�=�;�b�͖��MG#O��� p��i�C�6Wڒ�@0�v�����le8"�1�S�5m�$&p�CP�����}۸ ���2!�#�@�9\��� ��&͝ug��[B�=�f/y���|·V�_�Ά�����8�0�)C�\I�.�/��"ύ1C\TDK�7���o��}���՚mJfdL�D�3�%M4x�Q�:��7�g��YS�M�BP��I����֍����R@�6��9Y�c  u��Clc+�H Aа>xk���k؞*�5���7φg�Aq��	�1e��l�P�hF���� 7�F3� ,1���~]���[2��k�H�In��k܋ɍ�Y�)�q������q���k����Z$��fނ�ƚ�����@�3�mK�JC'���~>�iK�
�>�i7�wX3��e�?���pLN�)CKx��w�n����Ң֟�Y[��a�"/�X Q�K�#�r�m��̚Љt�CYZ�F�&�L��!>[T��D�q�fq��x�Ւ=�n���qv�0}��h�܏-� ��x����^l�t��I�����X��alI�F�9�q��2�3+�r��*��Rig�6��x��hq� ��m��	���	n�Y���N�i�҈G��&ӿ���Q���׷� !<)�䬫9�T(_*XS>��,gɤ	c!��b4��o�g˽Z���~�;Gl,�%������{�V�c^�5A���%Ϝyvڏ���ʫ'
�@Dc��%�E�c���`S����
ߦyU$�I-�js��,Xm;���ߦ�A�h�cZmX��K���%pA mUM48]h�J'2��'�H�%�N��������Z��{�<�>X��VrC��k3в�8�b4���`<k8��o�ᶢ�|�Fa� ��f���#��c�h!a�o��m�k�E�ګ%x�q�s���x����t�h����C\�祑ҕ��u"�u���t56��wJ�R�f<�vm�fo���˖ӝ={vC ��� ,	̉����x~�D�c��mh�[k����a��%`���[��q8�N�)C6�)g����L�1Z�Bj6�ZHG��`/Tqb�,L Y��f�Ƨ��%HJ�J��wM�����b�$�o����4�̙3'���M~�4R�-`}ܺ�r�m�4�O��T��=������;y�6ͮ&p��NGK[H�Dn��1��m(�cc���r�e�~������2�q�^�K�i�%m��Eh�i\���m�&e�/�cm��Z�i�:&J~��Dh"O�HWD�M�k[����MSfd�����<��B���� Dls�1�acq���)���2��1�c�ǟn��V�N�Ym��V�χ�.x66+��1���3�>N���	�1eH4��Xݚ�1�ZMB�o]/�Y�)e�ը5��q��bh���Ș 2U��\�M%94�}��%��̙3�cO@����g��[��֣��lL������I>�/��v�o]������>~y�)��v^2�c5�:��{]�Pz���qpBwL9��JHx��hp��LY����m�44qұL�h����~\�nƵfmL���˛�`�G�K��I0� @碁3&�o���v/��ˎ;�@y�` rɩo�cd��X����܋��mZ�-�c�,�Z<� r0�L��~�������oBk�Aq��	�1e4<�/.�G�xr����
֌��ڒ�"B��Ԃ�?9���()e��1�D�u�-R���#�Lk�G}4�/���0L���)k](�dɒh���ҥK��s�&�v�ޝh���e���@5���z���N�8K�s�6�}~X(>��!����&0W��A�o!����q�pBwL�ZDP�F�t�'��KmS��#�U��E�4[[MN����!�˚�)wjs���F;�
����m�-Ѵ��FĺW�ڰaC�w��F7��Z��2:24�(��`3 ��X�οg�]�]�\�/-���	�?��|�m߾=ڴiSԒ��{�Tn�-���k��;����:X���ɩ�9�p�L �&�$y�a:y��g�ڳb�*���j��?���br\��E�7���Q�98p09w |ϛ7/��:;�E�r��@�0eeæأ��#��c�^�j��74qrEchT�6�I�S�l��Ć���3�e#�m�L��.r�p�gϞ�>�ђc.\��-�ܒ�ҹMɳ.�hs�	ւ{�����F+�|�ƍ		3a���??:�����lt��uE䚋4|弓�'�FбU�pM��oܮ��I���������p���r���[+K+ֽ9�	�	�1ePI�L&)�����ZD�C6��n��p���`�ög:ۭ9��A2"?����8������@�;�ޓd-/�P'3Qi����ɕ$j�D�Wk)���ǵ����2W������5b���vVvFW\qEB�k׮�����&Ľu��d��m޼9�I�^E���:�m�:�K˲FIZ+�p.�x`],6�_���!�E���
Ǆ���2(Щ����Z��6R1����Lc�"Hk��ټ�t��{k���[��Ҍ��R�"ʝ;��6oz(!E��k��@��B��<<4T-�ƫ�M��S�k��J��w9|k[bf����ٰ-6u��m���g�쬕�-U�����5k�SN9%1�k�2�QN����Na���հ	<[��D�C�l�|C@h��-7��xn�g�5p���qpBwL)��R��t��mo�t��݆	��������Ϧ|1N�d���Q�"%��L�s>mZ͗�6���|��d�w�}�L��@���Goß�����f��>g֬�������с��}�l~������&��Y�x�h��^���><84���o�@_������B�mm���~��.l�I��3��V#^�d����y睗����m��1d�z��B�=QT���[㑊�3J���0��8�Bk�a�g�g�_�#��cʐoe�?�#��f����n}�h�i�a;�Zۻ��+̻--�1�x
���ҥ��H��;w�*=����{�����l���Wn|�����������w�����)=��C���f�<X=x���uk$Swu֬Y�ٳg�k׮��^���,�y��8iv����������?�q׺�Oݰ�������uU�\W�~!��F�2�Xڷ��_��W�s�9':���;�9�mTp����F�4_@��0m5!�����k�f���{0n�poE't�����2��L����l�y���ln}���G��c�t}�������n�`���l�˜^����>�h����y�9���կؼb�i��-[&5^�s��J� ��@����o���n���7�|ó�l�za�R^U(�-kmm/�f���T=�����E[�lI��0�h۶m�f��t<lS���s��L,�R��k�T6H_Z>�n�m�Xα��� R�Ǆ��2�q%S�T�{5.6
�X�L���[s{m�f`�͗�,L@�`�CHh��Q����JfQ\�zz��v�[*�7�\y�o|��}�[.~l���C��J����p �F}Qشiӣ�^������|޺u��ppp��|K��\.�/�F<!�j�������'Asg�qFB�ҔI	�7O�{��66��f%�o�t�\ �F��V�X'�HD���g��V�����#��c���j&���Eߢ^�E��h�H���(S�)"!�ɚ��EB�SZ�@+P�o��@��E$S;��ݖʵr���w����C=x���	�/��u�{�Uo��_�h��dj�Ŋ+T�uW�z������������������z���f���g���X���ך������Yg�utN��FᜰN-��5�+dX?����_h׸8��h�T��ī�)}��Bq5�fv�����e�qq�M�Ǒ�	�1e��q�Z�z�Cu�1���CJ�r&f�B���)� ��i?��x֬YI�ۮ]��O<��@k��'������?�x�ʕ��uyq�Z1�-[n���K���w���<�}�E���ٕr����@4c��Z}�l"s�w&s'�xBr���u���W$�HY�رbP|��@r�m�<�I@H����6[ �G(�f�c|�v
�V�N���	�1e��nkB�Z�-V�9�F�.gܒ��~�`\��D\�ż<44�a�ՠ������}p˖-w��}�����[��=�����.�/?O��6\wݕ�}�3_�����{[��3fL��$��"I ��������>��h��]�����7�15޵Ofs�T��/N�;[_b��u�|)��n3̇�5��;��cʐ���%*z�o�IM��昊U���V�N��az�>Ơ�̿��O�>-�P�L��9��C�{�+_��~���a͚5�o}�GOe��E��������=W^y�ۺ��՜9s����e[ZrQX���s�|����w_�ǐ����Zٯ�6뮠����F�v����ǖ��Z���jx�V��9�(�X�t8��c
�q�	�wm������&�WH���,m���.�T�������?�u�-���O^��K7*�:z�@�z��ۗ-;i�W~c��~v�Ιӹ�Z�sqX��ށ@֣I�;}?��C�i��J|�2��hF���5�ٝ`C\rY�U�khC��@�Y,,���}؛���"C�s8�N�)�Jy&�Ԩ�Ԯ3�CH��vL�������栏	/�Nn"%��BW~x�c[���C��?|�yZ�9��(�={�W�ſ~��M��zL��=?s֌���ۮ{W5�g=�Y� B��F�4��B�n��A+GCO�M���u��R����<�R9.���~r8� ��c� 2/�/t[���5�:�Hҥ`��6�[�d�vڕB.�*��5oޜ�={v_���z�?��?��H�����~�/��_�z���G�K���#�E1�g��tU�y����OH]k��i��am��I�}@@�����N7<j���M%�M��<�P.e������#���2���5�c��\km�A4o���87,��@ �_��h�����������ꗿ�U�����&s���~e�~p��}���۲�?-�2�2�\�Sow�E�+�`�������O�:Y6D�t~�~��,)S�G�4.�oD���|�R��>V��$��¹�pLN�)CK~l'.�N��^��H��Gf`�kَ���g�WQ��V:#�Z$�y�	�����y�yg�3��̆����+_�������/���Z��#[_?w�1���r5�Ǵė^(�E�6=��H:��=�����u�u�;X¤����ڈZ��}�.���/z{2�Ӵ�d3{����VR֒y��[\��5�����2�y%���K�B������f�ʘh��T� ��&H�r������!�Jc���J�2ǯ_�j���޹�h#s���.��?~��O�<�i�[:;����V���&	fS_w+��"H ����Öυ�����	�Ü/��՜E�)r8��cʠv��N
�dKcڕ[K��2Ul���`,ơ�)�Ϙz)��a�K�Rh�N.堩�\�l�e��ԧn>���G��o|�=�i�_���|��|>{fؔ����kMdv����&�T>�ꖀq�м�	yk?��<�N+Z��`�6q�Zʆc���pLN莩C��	�i���-("�H����W��	h�"���CdD��L�h���!��wo8��w���2r���nݺ�ׯ���n��֏�{_��R���'���GQyنKBkE77bpY��E������n{���x��!H��ɹ��p��S��_YȚ�p��b��a�P�D琂FMD��)k��]�/���l~ы^���ۿ�+z�`͚5��~��k�ly�ԭ�n��Bg���RL��J����O�� 6ۢ�6Q�<ҕ���7���9�`E�Ő&���pLN莩B\�TBW �}y[�+��,�Z3�B��99�"s4F�td���1����opp�Ƌ.��G���p���7�뮻�����r���|K�etdt̺�ͪbl�>q��4{���s뎆/p�n�����:��a~������	�1u(���5̨�íV�.bbS�о�&��D,�nǡ"f�z�t���w�駟~�s���Ԟ�r�o����?������;V�u�Z�*ytV�Z�)�*�QX�,2XK���`����q{  @������.^�)��j�p8&'tǔ�XɆ�x.�e[����!�s��h�J}و�e���+BPj������F�VI���`,�4�����;^��+��=�v�ڡ�����=�?�r��|>ۦ�8���H]�g;�!�YS9���اc,�[�L�BZZ3���Cw8� N�)C�0-[��+#��֒�EӦ��&
���y���$�Ҡ]'�v���m��d�ߜ��B �}����xы^�=�q�����n��U߿���s�2�BKR�^-L�N�ے���i"�L���ȧ�Zs��*q:^ϊ�|�񋄵�Z�K����� ���+P����׷���l�4�\r{7>'���GFDĥ�_7��" �h�����jrT�a��c���1|�uK@������?��E��D�`�:�_�����ƛ�|M ߶�`O&�H�S�8�LW�Uʵ�(�^����!��5Zղ׊=N���ͦ+&f�H�z�q>w8&'tǤ��-[Z�����x��7�$�Y+ۧ��D:7��/�={vݹ��K���I�|s8��*"�W �
S/f{��j(l����`k��m>�x����{�I'����w�;}z�� h%��$�D���M�-Zk�s���xYRl�wk~�s�YS��f.��nl�s�cq�X�����Cw8&'tǤb]u]�����=��}�_�t����Yu�
/��?!\�� bK�6���6��ch椵A��̅0�Ȍ3?�䓏�"2��իK��[�l�{Ã�L�5+ؘ���ٜ 8����Y4�)C��t��%��9[P@��3�7Pq��qpBwLT���_�������ӧ�	�]/���{_C�#�	߸��(
�ӈ�vP�X�;���9 s�B*vuu=H���v8(�}ݺ���������{#H-�r5Yd	K�!_�dI�aÆC��7{���l��'�<+������L���\��<���8�������x~6�;��������a�.�϶=MW�yɔ'��V���O[O�B�*E`����۷od��������xs;X��僿�;����k����Y�j%f-�̖.]m޼91��ٍ"�������6[Ғ��в�Z:�qh��-Sq�`����2���pLN�I���۳�7m^>oޜiz9��2W74i�#qK�hw�H�x�[�:/v	�\dM�5�sη��*Ł0�H"z�<������{���o��>+�h���s�FAj�A�E�+���<����d�Y��6@�m��@��ؠ��T,�����k���4��x!��1��]���������vN��)��x�c��E��N�8A�b}HC�p����@H���W�Z���s�{���]�����(,��(]�H@x�s��9X/�iXLp{P@��5O*��T
=��������G����1a8�;&##=�{��5}ƌrՋ^��kt?��c�e�m�i�S�_�����~�^��q�1�<S����~ږ�\���B�5��ڂ@��F�3�E��ڢ�b��<��}a[g��Ck��p��,��_�'PK-�7�?�� {�Ϸ���A*�݇�pLN�I��H���6|��zKwۢ舍p�DҘ�m���,vL{.�s�{�K���ox��7�tS�hb��Օ9���HwXE~��Q���� g�[�9~q�9�˶�E�B����6�^_�_E��2�����4T�����-�6V��c:���'K�闺Mj�[#y��4y�TӼh��1<mڴ�%}�#�ʼY�{������e�g#<��fS	����Sg?]����̯��f����R17:�wBw8&'tǤA���k�\�fp�(v�[�9Ǥ+����Vm�4���ͺ���z���P��g?��}q&:�����K����F�BXR�� ���9ڼ������6J=�3�B��>t�c�pBwL��Gn^S�"��A��Nj��!h[�����[��|"�	�h���Թ����c��E�ӧw�)���J�er'�A5��g]1�g��4��ZcI�ح��
c�S�i�g��\1Wt�� ����j5i�&�*n�p����1��K=]� g�j���5��j��E �R8fdժUN��`��ٕ|>w�VIVv+�Ղ+�4WI���C"����)<��1�C�<W+�M=����pLN�IC o�gΚN	�

r$��Z�,>WE�T!����mYX���u�! �Zc5��.��>J�b5�vQ5�ѬE���VK��[�;5�َK�x�y<;7�s���F��R)z���1A8�;&�L9(��1/��K:J>����C �~�ַ:��~�5MS� �ztu���������i�\&W.Vd6k]m����=�H+�ZK+oomK���cUQ�:Aq�چfO�_�V֖��g2����pLN�ICu4�y���e3II�r��A3�s�hq�QS]��b9�qs&�-K�:w�k�g���F�6���SX@�?xp�����x�}g猤������p?zzª岕r���\�9�ZJ���#�d,yO��2����W��E�z�h�V�;'�
jh��L���9��V]Cw8&'tǤ!����gkq�|�D��b��Q.�<�R#�	�@�$mK�Z���z�4o#�mc�r�(ͱ��}\;�A橋X&P��D���'�Zےҽ��%�[��A'�mߦ�ѬǦ�5}�I퀜�����	�1i�TF3�>3���]�L�vӆ\(e���e�L(]:�)kB�����aX�j%Y\�����E�W���M��e���}���#`�gA�mg6Z�&��٬G�;��c�P�$o"��2�v\#����J=@�Z'בz�r���u^��s��h�V�G�$�8:�j��JBX��a�*��"b2'(.��3�\$Ҫ��!l��$ۈi�%~y�D��']��T�1ua-?22���1A8�;&2���6^�7i�r�EKl�P��Ӂn����`!	��hy�\���)��9����Yi}��
�d�Lbf/W�Q6h�#�#�3�v�0���*}Xl0�C�֒�9�'S�j���������pLN�IC9N�nr�O�0��"��r�$��!u�|P��6k!���&�l��tE:S����֭� e3x.�cb��0�gVȲ�P��"�P���EZ?�4�ё���F�cBpBwL�I��X��k���Q�����kL}v����1l�9��vF��_�jR�7y~�~"He���^mT���[���U�ZB��t,�4��4j�:�ɴ�߿��Q����8&q�+c,�R��h�b��T#��V������z����-�My��4��8L�"��t��-'�<� U�q�8Q�B��V�A˂�5�)<��'Q�"�Y�f�� M�w�ͩg�5���={v�Ңg��霰O�5\�%r8��c�P��窐jbF��_�C�@�L�D�W} m�K]C�䮓ʄF����f鵍_��j�QkkKy```(r����|\)�ac�5�d�A��ϥ{Ͼ�l�믵�F����r��g�֍F�gϞ��!x=랞�hƌ�oA�O���w�޽{�,?r�D��W�	�1i�f
*�Z��em����LcӾ���H]�|����V��u�H����ᣵd��@���/A���7i�%�_����Q���qkͱph������"ܙ3g6��	�(�J�5��\+zN���9s�$������D H*�Չ}ѢEq �{���/����6m����+F"��qX8�;&q%��-�	�TjÔ��7��R:[�T���������v��!}��$+2֋����Ϫ��K#��=u�HE�X�ԍw���Qk[{�'���+�r%Z�`At�F��?�s�v�ڕ^�D�"����F�5J������5��}�"'sA�jL��|�Ϲuǎ/y����~��>�-�?9�q��4��e𕖊�DS�o�U�]�ૉ�vtto��`�z�5o޼�K�����7�it�4G4?��t��l\����ݕ�]vY�k������ᗽ�e��%节�ww�JK�-bݹsgtꩧ&�'.-[Ӂ&v>zu2N��#���i&w���SK�߳gO�� �ә��K.�dq����<ou��1>�����;wu��0cFW�	��^�IC�L.����s��]�
���.U�Kj�O��4A��>�H��I��}��'eI�-?{�`��/��	d�3���$\��^��W���}o l{FG�g2�-Ӧ�׬>+^�vmt��F���w����aB�"f���������g������)�g�g"�J�������X瀎Ӹ�{n�q��F��%�����P1?��̏|�#�G����#'tǤ����%�ͷ'>�
Q赀)j}k{��c�1Z�M5l�v�������1�ڠ9��z[��N�pr �J88���_����/}�p�ǣg0���k�;�Yx�k^�v�EE�6m��:LKȷ��3	j�h�hK"枾���N���l��D�2�s�1��E��m۶d��qxn����[�n��?���^_u�U���?8���cRp�Wf��?�sz{G{R]�X�U(�&/u�*&�L��Z+&���C��Ah������x�]��:Nۃ��0�12A0��Q�>}����}�m�}����k�߻���<s�Y����oƏ<�H�����Hb����S+.�jYF�A'�X��������D����裏&�׋�=ni�"]Sψ
�.�^��߫�t�M~�����7��ȵs��pBwL
���x�����/�x��k%A��k��L\���Uk!�'Nu0MB�%o;vQ\D`���:�@��6w��d��C�P'��}b�F��o��ovoܸ�SN9e zAy罽ݧ���]t�7���-_�<Y'�J��k�Ef�$���hG�g�)=_K��k1��.�@�O@���H\�OV=c��l٢�G������?����e������	�1)8��3�ׯo/�DC��3AK�]�d�4Zdj/}WYd��k�m߉_]M:�s:�hj�!��}-�5�`b��7搛7�ew�}�;���/���L!�w���=�%�ߦ�[���ˌ��FїYs����vB�����r �L#͌���3 ta)���Dp��ko\'|�[�<餓֝{��㋑��8,����@���f��;(x�JT'�=�k��r��~����߶�y��n�{m���Uk��r&����޽;�t�ҵ?���?�Y�n	��h'�p�����J��C�J啗\rI��Yi�*3w���������b��i��Jb���h��ئ-��^�4:��v������p�J8�;&�c:��Ѿ)Xb��;]�ݖ���_��q��m�r�ڥe}M�w���M�ԵҎR�|���O�;�Ӿ.�':J�׼&����������nok{Y ����G˖-�{�h���Q_�@��!Xµ��6�3���H9$�غ��E�g���U�Vy0���$pBwL&��������hhfi{ZK���
�A������F�m��MYR��ځ��G�<������vo۶�@lG]%�u����o�rꩧ�SX������+��r���V`Z6�o���\l+[ 9�l1����c���f��`-4��-A�'t��I���B�d�>�"K���!oH�f2kv�f��j��8]CU)A��:�L���T��eLEk���1��ٓ�����ڵ���(R��h"u����ַ.;k����r�3�g�����!%�x9�mI�ǒyS��D(�Ե��O����m�Դ)��{��p�3�F��1Q8�;&�4���bb싚*b���!�kN��W,!0����q-yq-���7��]D�w��F
B��
�-���z��z׻�7n��SNyڗ����?�p��%��׿��k��6����a
W~��U�C �2^��}�ɷ��h�i��~��H�}�|�]+��=�� ����@����������Əm�o[���2l%1������Б�9]���sT8#]�*�Jǉ�4W�LK<ik���_�r�_~���iӦ�O8�~E�EOS��W��j��}~�ӟz�M7�8������r�����=�����k-%�4{����Xc���=/�kN ������f���<m���*8�;&��F�&BZ�/}H���.c����'=�G����Ơk�4t�y�۵_ک>�*qw�ܹsVM��o�ۧ_r�%W��=O7R׽<��#s_��׾������z����w$��E�5Y/0���%�`��C�]�#�_��W�����ٞs9�#�y�97��������	�	�1)����&���3iP�Y3+/}������5�9�^�`G3' ���t_�$�)�������5ڰ�0vkGG�[�n�������/��c�?M:~)�|�O,�>��w�򕯸ছn�+����P�;N/z"�1�K@�*'酬5����#xk�c�Ml��l�C:�N�]��&w�cpBwLv���Ebl��(�yY7����+}�!s.�lM��Z<�g�6D���Z82ٱ�m�R⁁�| �僃o������?����eݺu?_�f�S:/Zd~�]w���w�󺗽�6l�0��o]��\�(v�����l��M/��[�"8�sl=�%O��io;f���Ω�����18�;&{���L��S�&!�ҍX�����F��,�Eh8�_s������;�,���ծ-�;x�`�Ph���5��w��Uo~����?����<�T����n;����5]]3�r��/�HB��{,և����7��&i�=����*i�SmV���Zs��6�1��(؈z����
����9��cҠ�8^�����\혱)PM�3x�/�5�d%��7�8��}��|�
�K[��9EqS�)��㞞ul[�����O|����O��믿~�_��}�S[�l���7�y�O���m�b�n���9۶m�W�XQog[i��)�kc��i��1� ��t�   X�ipX`l���@�Z=(��p<	�����B��ՊB��tDs�����`��,�[���ٜ�.�PGPfwL�6��x�T����5�����j��_|�'�ݼ��S~��~�׾���q���}�����Nu����w�qǴ�~�Y���7.ر���ٳw����F�;�d�D�E�S�F�wW�NZ�����t5��է��7搪،����|�G��BHyV��*߮������$pBwL
�KW�pY�\���(im9��l5E|�do�{@&��.f����i�i���1��؊�S����788����qBkk�;���{����8���3ϼ�G?����N;�wѢE#��rM�;v��s�;��믿 ��o<u���3�=d�-[ְP�~����N� zK�{�53�t�!kh�^��J������<��X���������1YpBwL��l,b�~o��f��b"Նv)[mO�P _�{.�4)�0���/;���m��KA>W�$��m�Oi�J�
����3ٯ	�O	�~�<���_���A3�oŊ���_����~��w/Y�dh����@�#�S>̽-�̗}��<����0��ɽ���+�r�t��F��L�Z 5^��"+�R���j���!��/�:Z5Z��t�F���Hw���f���#��	�� �����B���*��[��a�J�Sk�5"�A��B��+�Z��,��t��h��i���tB��4�X�H u�#ō����R)1ǫ�h��6\{v ���mٲe�=�ܳ3��p/ۃ@�D��������+W����Z�|�@ �R���!D�}�e�}��1����7��_xj��={���(�33\3���-�|�W��4ԱQ�a�H����˚i�����c����1��R�J�u���}2��㦣���"�0�r�4.��pL���i�ᥞ988gs��i���<�/$�[[�B(�����r͖��Ja������������99���r�7>�D��k>�L\�87:Rj��Ӿ~L�I�B��/ɤU�J���d��B>�ƙ�5}��p��2�#���o����?�����mG�VOK���������u��c���Y]�ֶ�|�{��@o��];;�����	KyB>�_�dZ ��qˎo%Ȍ�r�m-B=�$�ô��C��toI���X�\�:Ѭ��=HGM 	0�;��G]�(J�����	A�@E�� ���"ݓm�Jx�N�����$t+0�8�j#���lB2"��h���6"ة�nk�7	�4&/��f�Fs���|nkɧ�툾G˴c�d�Ay���mt}&����o	9�ӦO��꬙��ĳf�[�T��K}}��޾��Ol+��l�`FLE���;3gvee	cdR� ���K	�Ep�sЦY+��BA
 q
6��֩���?��6Ү�]'�?��a�	�� ����R�+�y��LE��(Cc
ΐ��*����k�YM��gAK�Ư˵���L��Ѽ9�Z/Z������hӴOp �N���裁r����t0�%N\��	=�V6����h��(���s\��u]z����C��fvi���ri�G��Lm[\�d��Cw8& 'tǤ!��ː6�\��e9�f#��@�휦��&`�Q��\s�ݤ����4��BF6*�NmV�H�C�W�X7�تki���-�Z����X8R�\�\X'4z���O�0t(��p�S<��`4��=mA�B�x>t�K��B�p8�N�IC9QAÏJuA㙄[�;A�L����jCۆ��Z�@��LmS�9���̧��!<\�50y���J����(��0����-�ZK~�tm�%P�c��:�.��ӱ�L���v���d�B�8�=�}�<�s�cbpBwLFGG�c|��f���p�e�9ZJ��4��4��,�� g�
K ����N�0[���f�o���˚ڨ�83Vӵn��[k,dM?V����$���q�&�	IV�8�m�5�[A�
*h�%V�`-4g�CH���B����:[w���!il��˹����	�	�1i���u�t�E���$�@ Q��ђioJ�5��>X��2��y�}m�p4G[uΒ���q�*i���۬v�o�J{Q[)M���O��h�i����TnM�i2��𙯮aׄ3�1l�v����l�w��]?�`�k�ɽ>�j�Us�pLN�IC�<�6S�W��m�RK}�fI@�&����!B���\݌3�а)bB��f�t������x��8�Dm5�k���ǋ�'�;-����I���,��AʘՂ�h}pO��[��>�t���E:���C�t³f|k�?D�c� *W[����p<)��������x�82Z�gk�b�$��٘���|[Z��L0�CTz񋌈>��yA�h?ft�����(��&&g@J�����u����ǌ�� "� i	�&H,m���vL����H�l}z����~��%�M���t�/֕� �A���Yµ�t�7�v�s>�5�[����vK�c� jϷZ)W+-����	�	�1)8��ҢE���oCW��si�A������A�uM�_M����}��ϥ�	ĈVk[�����l-�79�ڦ�f�Ho{M�Xb�/�-mk�𕋐B����,�;�s͟5"�M�)�����1�[�7kI��I)r?X<l�?kg�p.�h�{!�\�
^i?�d�2јk&���%'t�cpBwLN(-^��`xq'>�@{�e]k�Q�e3y�Wqdǐ�%Zr�mu::��'>\��!nϷZ:���w.�\ċF�y�$.�m�NK�}}}�f���>t-}Ϟ=;�޸qc��@l ���h޼yjȒ�c��m��s���OG�[�7dm��bA�z�QMZ�Ќ�h
d�������oc$���>ʮ�;��c��<SA�4ҡ�/�j4��/�F
c��C��hl�6K�fg��cK�B���vo	�c��c귚�MgK�",ҬE�Xئk�[�ڲ�~���֭[����2�$dNОj���̍�����T<�v�p�/����ç���5������(���?�?��w(r8O't�d!7zp�3RUti�E��EJzi��:�d�\~i۠���	�بv�!�Zǣu��f�	�X}�H��2�Sa-}}{]K�6B�����y[d��H;_�re��LZ7c�]�6���D�:�j�5i�j����E�[A'9o�/��:�~��#8�y~6�}���B�Zֿ�8r8O
'tǤ`���������Y�DK��Ҳ���I�7I�I4�`,H*M���m�BU5|��rE��[�1l:�����V���A�f��|ͽ�/��gϞ���o/�>��c��%��4zAsR���W��-Nù��Y-�6J�>�t��=��-�c�h+� ��Z����Z���c���x��qU����xR8�;&���lρ����楦�QXmؚd��D-;��F:����8$�9��	�������mj���!n��Y������v�݈�'� 7��eN߻wor\WWW"�g~��w'�,�NH��2�"x�G��p��m�۴�����ub�[ �Lڠ-�c��D,�#M�V�H:����1������xR8�;&{�gh���9�Ɛ�̿��ٵ��\>�|>k4�(�,���A6�Ȏjn"A�%�W�G��d4CK<h���ui��>��Ct��_c�OvٱE��pK#לI��G�v]o�����"�}��%����N޽�|�'p�����y���m� Z�̄t<�޳.�&v�O7�9�U��5t�cbpBwL
D8�ś/H���t��ى,3�^��Q�/�R�F�$x.h�墢�j�sx�WJ�(��%~�b)�y$�������� 4���B�S�7��=��:m�9�v�o��݈��3m\�9�$`�0�Mk�\��1ݎK@ߺ�c!W��,m\į{�ʛ��o]Ò&�<�6����*u:�5�*.��Z=cb��ؤ�i�-Uk��YS{:�0Y=�-��p'tǤ�\-g�9�RŹ(W�$A]z���EJ�:!ڸ�;�^e���B�ML�^3���upx�Q�E����fM�i��	qCH4KѱҚ�� <r���n��m�X,Ok���a����+b�ٝxG1�SkFD9� �Ls侨��iܖÅ�YW���q��L��b<+	״-fy�D�Ba���g���6%�R)W[Jnrw8&'tǤ@��R���%�ׂ��ftV{zz�:;g
o����3�eɹ&�ܚt-9Px�P3��~�{N:�%_ư�ZV��>����x4nk��%c[r�2���!=�{���xi�n�C�\�o�2��4ϵ	�CP�v��
l�U�O����nQ�ܩ%���7�`s�m���g5z}3���pO�L4�($���8��cR^�q�T0�
�˽����?}z�5��|�}��O��𢞩c� 7�ըR�M�s���VMȮ�lP"���g=��_8]�r��Bl�I7|�&x,0*���g�Ɣk�9�"vی36�5}��ł@w�m{�᎕ a�v�CsO*�.�^�AlA:� �]C�$�J�>�#]�>��V���;��8�;&��s�L)�/�H��DS�3k֏��S���;���o��W��huxu�T�Z�8�j4��|���DZ/�f�Y�x�G�dd5n��v�&���d�GHA�2ą_ئ�!4��sH��P$FQ��5�ĩ��+��l�<�� �3�M��1�',�=M�X1�UoM���x��jf��>�i�<\!��M���\�bE��;��cR0~B�zYW�/������%��Ͽ�U����������v��].��ڒNi�5�l�d<���C������$�hlL��o� @XB���Hҹ��]�� `[�1h���-^c������+9�:_�Ա$��Af|
�P��Ǳ�����5§�o���c��ݪ��X�/OG�ۜ��GHW�҄�Z)�
N������ݛ������F���;G�/]��qˏ��YkW�^Еj�������ϩԩ�����Q�p�����T'^�6OZ �<�Jù#�ౄ�TE>��D'k�N�Z>ިnW}T+I�Rװs��2�d��uʕ�w�4�[K d�F.�9�Ҩ6���7�� c�o�fK�j�#�<�V#�Oǒ瞶,�1�`��G�� `i ��<]9�j��m;T�*7��XW;W!�/oH��$�R�5t�c"pBwL
��-Ҏ�@ �����+�?��3�<��V'`��dx;W��@@9�H��,r�]�3�:�5�6���uSviLd:$�X8~c��Z�d��!K4p[T�c�Ek��[�*F�%+��槏�ӷ���A�'�\��m��<�
� ��Sȟ�G�ڞ�O3�?;&r��jۤ�aA�.c ��Ӿ����̧���O�&w�c�pBwL���r?^⛖,Yr�ν;���o�x������x��W�4h:��sQQ5ޥGͮ[		f3usq�a2F��,�Ӈ�F�t8ȆT/���E�lMt9�%Eit���6��q�W/R����@�4�>�̦�i>�=�cD䐥~�ǆ�!H�S\�i�=w��d�h�
��86�N�(7]��4��p$ �o��:���јj,��n���Ϸ�t�EB�-��e� kf��R���:�;��c��h$���z�9�m��׽���-~B�v{D �-g��>R�i��^:fm>�����r#2\�a������EOs��� ��%2� ��>4j
��
mT�k_7�3&d�1E��͵�W�ӡ󷭧����`��r[�@E���8�Cצ�����y��������گu�1Eole=��ma�זֵet�P lPa� 9�rw8&'tǤ@/�/|�=7��=_(������f��|���:)D����.@���P���5��@����D!�{����m��HS�F��/*�*�����&�i���u c�
��-@�4��5oi�6g_cRAN���S��1�h�O�	:O���>� �d�O���9㤢���ܬ�Ǿ�i��|��Ȅ�\Cw8& 'tǤ���Ǒ�9������IwUi�A�T'�\-X
�x����M�=��[���h�UL�Dl�%�#�M���L�	\$(-U��<kB!C`�=Ō�oi�j���@���u��}	?�s�ώ���A��4t�a�dE���W�w������㟷���&nb�k��b�47����c�����ڊmN�����2�--��R9�/U���|����D�}w[�z�O�oh���Ep�A�>^��e���'M~p��.l�[��
ڈ�		���q�7�Yd� 2��F��?�Ùg��\��'�h�oӘE�KH�<$|��5�-[�D˖-kX(4W�'�}���m/_�<4�����]�yXB���qv= k�>������f������pLN�)D%^����gv��`_�>!hN _7����'��]V딆�m+W�SeN�En�xE�"K�%�������=��Nd�R{�'6��-MY=���F���\�ҸE�*
v��9��,�Ɠ���twwG�W���?���E�w�ƍ�������o�'�@��4�Ơ�]Z���]�M8�ǎ `��a4���y8�;��c���j&��,Ep��[���d[-�jxl��(�ٛB.���R�iX��i|"b�H�]�b�[~jAu�E�v�J��^�;Ae��O>��D(����C5ޞ��g'�	���FG�T��9�@=�!2&-N�Pou]w�ҥ��͛� 7�E�g�4$$h��nݚl_�dI2.���ú? �t�t̃�=��áD~���8�	�	�1e�h�(g2q��2ǧ-X��iN�����m#�I+�ER(��Y�+h���E�"W��Ҩi1Jq���>��&m���j�I'�����kLj׋0/^�#��ι�����?!���;/���i�j���É^�k���vݳ�i���W�Z��%��IPИD�N4'	�Z��F��ǖye)������7��Ng!DN�Ǆ��2��ŸA�2��̫Һ�z��8*���d^l�i�8��q�6���Ym��g�=�����[U��'kFY	E�IB ����x�x��o��[��k{Y��7�k��m�&�"��B9e��4�M��T����s�xj܃�=]]u�Vu��������fl��tՃ(Ar\�}Ԥ��8%W��r4K��Jgp�=���%2i����׻�`.��A��\��r���Y���9��s>�0lٲŵı��}0o.H��q�-[��c���Y���/���QC!̊�@R��j"��2�W��3~�s�-�[��54zM��!������X˟s����2&U)β�A����@@N������V�DA�t���Bk��n�`�b�9����ǂ�
�Ģ�V6��a,c!~�~�ǁ�A��n{,��&��˲;���" ��N�0�=�y �y\�ƍ�m���v��U58��3E^0�ĉ]k��,�S�*�2P��c���XR�빠�<.�k��$��a���F�	]������`�>��³�Co�u�E"ay�����@^ ?���Xf�Zn51�u� #�2ݽ{�{�W�� ���dR���2E�8�g|䌹 �����Yz�����������j�I�t�SI�K���q�x0$@���W^�&�Q����A�,�c�u
�Pڕ׌9�u�$�|7:�OW�N�%�i���F/�	]�`@�U�N�o���w�=U�;_`���j���t��J6��>ȋz�jV6�`\�͙�҃�
���z�R� ��|i�sn؎mX`$�����Ď��X,��I�X$`�n'�x�='���L-5c �G�:�0C�B8���y0�;}�t7V���g�L~̛�q�Q�}�9��C�7�9�m����������$m�����F/�	]�`p ����%G�5��g	�J��]s�Z�o�8�8��21�\X԰V銧;�qpX� >d���놫ċ���;v��ׯ��!�k`�۠�Mj~R�׸��&;H�� �`A���{:΅�>���x�~Qy��LIX�
�@���\��T&1��Na.��9V����u���0�����KhB�((�}�t%j�q=,��r�|��R���Ԙ���:4H�D��;-yc� AƎQv���8'�Ұ/�~X� |X����5�h��x<�qvf�c,.(�l~���ظ>x(��9�ܘ�#�ya;΁�y~���}��,XX�� 8'��S�8]�sH����i�����:���%4�k��6�p�o�Ϗ���=r��$��U�D�լk��)���� �^�Ȱ`;p}Sf0��A��J�~ O��a��U2�#��R4̋z��Y�&g�rn�6;��h��1s�/��;׽b�
q�y�Y�f���j���z)\R��J'�����sp1�.���d�}�f�5jf�=�r~���q���&M���&t���0�u]s?�F�Lg�[�t���)
�ʎ���� v4���@�l�ʅ��N:�}����h�� 1����r� c�\B�{8?H���9��=ͷo��>s1B�Vu�c��g���=���<�ӱ/��M_X��z|�a��4�Ұ���q	v���6x,T�[f�3�Ʉ܆D���M�Q�h8-���D�k?�ʌ�&M���&t�����"��N�+]�t�l����Ϧk��+ (�|A��� � `�sƥiu��`lcq�@�Ź�k��f)���s\샹�e`l�+���z��� s�ǀ�U�������>\,�o��c\6����c�qi�3dA+�^�k^I�����V�a��maߋ��Ɵ�&t���0�0���Y؎ݝ�&����&ȱ�
��� L��cV���@jp�S!�$���iA҅�kZ�x�ʱ�
�f-7Ǧ�
=	�Aθ7�kf�#)�r5��ur�z��u�kĂ1p.P87����� Z��Ӯ�8���7�ٹ�$0��r5>�ʄ�d�w���Ca���wjū���M��s��e_�n�?�,y"٪�.��H.�u�\�I`��V5�A�t���QZ���*��m Vzp,ȑ.oꧫ�.j}6�G��:��l{Z���3���g�9-\���x�h53�M�?u�Ƞ�S���o06t�Sz���cs����1��v���q([��&t�����\�;�����͕�u�fI�̠Vk��?ɋ�yٷ��JE7ČIn$~��A�Lbc�Sʤ2���t�S"Ǩ��p�LRI��u`���"��F�T���C�&p���5�u��{�V`,�Ϟ�׬)���E	�*��T��'�]�����	]��0�k�i��	q|���r(Z�j�NfbӒ�+�V<H�I˚q{��ti�V5�&'ɩ���uҙ���U"#1c���<�(|��ߴ�1���Qםqu���H��|M�U3�yO��x��qq�EI��hT��T������|��U�ejy�2�aBCC�WЄ�Q0�_f��Н�,���^��#oZ��9�`@,$,&��B#a1��$<�G���g$`l�k�MMbd|^��f\Z�|IvpScuN�F��I��U�6^�"�V:�}���s2���8�/�x���c��z��by�Z��F�{��8B�Q��-��r���=4�k��m���t�	��t���~�;���$?�߬��RRc�t)�=�i1��%l��I��뚍_��&����8�ڗ�.&X��=Ak�R�$h�� ��
�0c�������{�E Ɓ[���u�؎9bE�=C���C%m�3V�1�煯� ݜEC�wЄ�Q8d;�EЖ���rw�������# -r�������lt<���k�@���f&��Ç]72��$�9-uzp�*v\�ؘ��C�u����5wa�p��a_��ѺA�\�&���+��Qnׁq�/΃g��q=P�üp-���8p�K��a8���T��X�.�+z)P���qZ��FW<�>r�H��!}�y�� ��a~��K�t��d�k2���%4�k�����B7�{�*�V�����j��wg�L���q^�K(�0�u��|���.�HQ�"9�`i��:ǧ{� �]Â�x 2 	u(�c2^�$�V�СC=J�Ə����x��E��AĘ''�v̙-U1/��!;��؎E ���pe'7�p� ����
����ۗ+K���^\=���MlЌ��Aю��L~��^����:gB����+mS_�����lMC��Є�Q0�)�g"yY�NVP��Aw�1h�;=H�.u�Va:ݕKjS��@2 HX�����ke����1>�gM;��1cƸ$��p�����ٓ�Q��+ȑ�y��7�9��aUC����8/��q�=k��<h���A� d&�$�c���8�o<��u�ܹ3G��#��f̘���c;�_IƘ+�O���!C���H��e� ��Y�G��ȩej���}ާϟP��1t�^B�F��xfw���Q������s��3����wu%suд��a�d`傰A� ��Ah pX� ����i��}�1@bl�r������a����Tǹ�0�5�9���B��|8ƅ��R�x��|�`1���lx�戹�\�3� T�ñԗ�`� ��`�C.�����k\7�ƹ�7]�,��s�vf����'�uz|G�ZtG�7�{�����	]��ȯG�L�G�Tw���?	B���,u;�l��j֛���L�8H��$1��@r<D��e"�]@nT�c����B D��t�)���5H�˕:3���uC_ְ�1o\��9�+����s^?�vW���m����Ǽ��� T�O6�!���~j�:�����M䓽j����:)NC�wЄ�QPdK���\��s�2 ��I�jk��U�Q븹(����]��.g73���@ΰz�G}v6b��c ����`��v���=��m&�aj)��7�2f� �c"��.l\�`a�q�?��1+����u�������׌��b��<�§4-��Y�1�?��I����"��1t�^B�FA"W	=�b����A��TK��b�Ϊf2-}�NUu�钇��1mC�uX� {�ÊQc_�Ǥ5&,�s�=�Mvcv8�wd�#vK�L���`^ |�6���bgB!s(I�m�G�%w�o���y�4i�.`RY z�յ`LZ����nx����#��Ҷ�_t]C��Є�QP�7�n����Z��$85���n	���Ԙ4��"�bb�:5Α�R�Һ䂀�'��A� _�����*g6=�NI�X`?\���f�8noz0O92ױ/c� R��qvcC� �F��Ǳx}��Q7��D��mR1̻��ڽ�� ���ٴiS�;��pOY�sb��G���`|��
&&r��N�I�j��m�q�Z�m���_��54zM���N����ߴ�O��*U��K�ԋ�{��Օ��ȹ/��A����K\�����x:���L<-^�հ\��Rv��-Ǝ��ټy�;��ɦM��{�޽��9���g���ZƼp� L�%�g��ׯ�-�fc��A�8��_�6�c���n�:1nܸ�;�Y���Zyd�c;�@<����̦*�+T��3���'���";�`P􇟛��K�;-l5����Є�Q0B!Gu�S�U�����8k�U�{x$��u@��f. ��[��j��^:�I(t��x �Ќœ�V�\�sU�r�ķbŊ*r�va�2�׃cP3��p���1H���{ pU����*>�$5.�u�ڵ��g� dNbgY5�Eg':��Qaׂ�b!C�>�/p�S���b̝�$��.�W'ɫ�^�Z��ɤ9[�-t�^@�F��q-g��n��<����̼&1t7	�b�$�ѱ/��j����\�bT��t=�;�*�
"$a�(�>����}A���5�5I��w$6���7�hz��Ϛv��� ��K8$P�����0�ۘ�����y����Y�x�"��U�\�[U\F���N8rOl���F/�	]�`H;��8���B��&&���r�~�%�t�;{Z%
�Nu߫�!�`l�.�G�Erg���$-f�3���$>ʨ�:�q ����zn<H�\����b�7ƀs����g4J�rlvS�{�y������q\Ha��!�n�U��������gb����Lr��i8r��<���54zM��a���5�pEO����s�St��%P|�SjSf]sc���@��d,#�r@YS9��Ԙ0��H� Ɍ�T]߬�"�s�B���V4���&- Y��M�gG9zH�Lh㸪�<���w�';H��r���� D����v��k���/�_Š��9�)�jB���4�k|�P��$x���D�k�k6z����e�9I��'jW/���*Hh�N�%��$qZ�U�=\�p�3y�c���E@�C���������Й9Nk���:��F7:= f^k����m�^�P�ĩc���G���A��y��{B�s��M��	]C�Є�Q0�A�~�=�0������i)��H*$/�+G&j	���2��]��U�KU�L��&�=��i}���-�Ο�g&�1c�qj��g�c ���Y��Խ�JH�5��YG�<2��> �a�=�e'6�UB�r�x�%z�/tūYH�8'	���j^]�2\^� �c���&t���23:��n�T9k,�нz���|-�#��U�V�jݫ.wUJV]p<Z���c?��1�αi�r~j6]����&+�Q��(��׌���A� H�1k��o�c��b���B�qz.F�?���c�y<x^΃��K�ͤ:���F=���6"��Jq�B���4�k>�JKr�̙m��gE1�u��H��Y����{�˞�e	���Jj���ؖ�H�/�f�S]�ǣ��"3�X�u�b���Eb��L��j2���s�%��m���,c�������P�b��s���}A�!�9���x~^����.ǡ�׃}Yi�E����Nu� t���	]C�WЄ�Q0�xI��cے0Ifi�f�27��>�/���b�*A��ҭ�ݍR�Х&�tq��y�ĉ98�W�-h���sj�Cq�IvtK����5��1_�vk�X؏er�_���ѝO�Z/�?��}��'2�O��g�L!=���t����dМs�8P�C�;Iwذa�e��	2gm;/؇MZ��ΰΏ�>��)�útn��,�֟�V��Z��54z	M�C*�6�tZ�rC���e����*�=yW�Gܚ��2,&��5�
��	2I�(�MI�x2ɒ,��F�2����P*�j�*�4A|x9W�%�B�':��>�5� ��1wZ�j�=��P5ܹ��yPR����D96r�RȜ�L�[��8���1w��{�=���<jS6�aF;��" �#������-���:GݜEC��Є�Q0��\8�<w�m�{���nZu;I[�hϷUK��m \�>$KA| c���4I��_��a}��������e�ǆ*���:��D4J�b_U�c�U���Iv,�Sɞ ��1�M��1y�d�^`���������<2�X�P���:sH�bH��Zp�#Gr5�P��q�z �4���5D�F�[r��y�/��~?�tb��F/�	]�`0}�m�,H˸QQץjZoKfS���qy%e����t_��e�D��/Z��X�Z�eIbT-I�L#Ӝ�X�(!�Jmt���:�m��8�����x�M�>��R�F)jͶ����ZI�p�3&O�:�$���� ��iH.x<ؖX�,�c̜*q�ze�ǦgD�P��s���l���Ɵ�&t���x�g5�\�QW���}����kf�3�L-c	�6���;���4Ue7,,V��:�$���no�����St����oz �RW_�`\�J�c���2�~��A�&L�5�@�S�N{��q�aҜ*	�{�R?7+#F����������.F���w ���]M��}_\�WM���&t��1�L:#YBZ�;�����Y��eP��ʛH$A&lq�	,qf�s;��h�2>"'�P[�hK
"�u
�<\��	"2d�K�p��< r���E�dϘ7�Y�
W��|��QEqT�g<,���G,P��X��y��:�!?��3C��������1{*�Q,����,,����;_�����F��	]�`0ip	�
���Fh�y��+�wʗ�d���V:���$3�&��`�.pǡ���E�����ܱcG�R3�wc<�;��� �����������jeb��,��?s8�S���N����1��
*��}����sE ��G�u\����)E���P���� ����ӑ����/��{r��	]C��Є�Q0>�1-IF�Kܗ-O{�lwU�\-_S[� @�p���t,�f�q��Y��1�)���Y���@"�K�:-R$�!>K�A� k�I��/5߱-o5yLm�L���a�5@B�ypn��a.�h�J����>���ǵ�X� ގ}� ������d�js��x���л�z�ք���KhB�(�>ͤ3N ��D��*�O��U+���ʮ�1eU�V��
GW0�ĳf�1e��<p1�2��
 *:-h��1��`��@��BD��=��qg�<��1��S(s�M���^ U��V;-_�y
=,��3=�{�m�s�"�����a�x`<\��i����ɚ|��&.��OU:5���/��j��J��T��>l����]C��Є�Q08�4�2�9�ha}�zXo�ej�V�jՑ�`v�z�z�3��
R���53�a�RnlǮe =�&��(-T���@r)�tO3+�q|
˨Is��g;�g-9��i��x��{�}"� ����4���*N79Ef0�����}p�,Cc�Eq����֞�z���d���t������E��&t��C�F�`�)��8����=��;i�{&!�?H��n#���;Ub� @ܟ���V�|�&���ؐ�0Ֆ����fګ���� UX̌�3�NA�ks���{����U(�C�7u�E rh�؟���YP�ȹ� ��/A��D#��N�'�e�$�~����4�k~ˏ��,!t�y�IQ��c��Uc����EJ�s�b�F1��MW8ύ1(����yNUz�1q��ty��ʧ�*	�9)6�m*A\��L�-M�k�)�B����q���6�" I��P�X��7��p~�������j ��7�9���7�p���54zM��$����;d]��n2e�ǗfV��De��Ԓ.5���Zr�qiU�ҥ����rf���R�}�j��Y%/�Ge�8�GW�Z&G+���o�!�uO�H�#�ҋ��)�4�����@����`�l<��8���p�8',uVp��AL$����8���.\���s�K����Fo�	]�`0,d�w[\�8i�B;]�9�BM�R�q��&�*���վ�t�SV͠?]�:�g\xa�[%r5��V,K�Tw=��[uI3�sac6K� s��~&�a���}N�v,H�>���9q��|��3V��q���A�\ C%h���p��Weyi����t��ۖch-w�^B�F�`�9K�1|~�߹�o�c�ݪb��K�2��E�&_�}������ )>=����j�G�T]ƪ�:�Ը>��yA|x	���aM<��u�m�Z�1Ԋ��z��:���ZqX�$h�>�鰨��̮����9�j�B	ʺ�9=�P{����i��'���|�^�1���c���&t���N!)�6��RS�E7!痰��Zpj�Z>i�8h!S�	eTQS]و3����N��LUdc�HQm[�sR�ǪIi�Cs�f��]�}�ϖ�8���t�����{ֵ3i�Ӣ�� u�7���o�<��A�<7�b�T��3\������0/����ꂅ�����!c�%���F��	]�`pLӐ?�	�1���6�*Ǐ?�E.˚�$d��I�*90S�,)��.h�Cw4�SZ� j��H�Zmъ�Qg�s�be�7� �u&�a���e�]��W�a����,}㢆�1��+\M8�1 a̙���\�� �?�� �t��Ѫf��!���ȯ9W�q���΅��}��0̌�Iq��&t�B��Y�����x��b���������� "��IHL��/�bL���AJ�ĉ�@b TƉ� G�i� Q��}�?�����$<��9Jʸ �1p]s1�c@�la
ƻqX�8/c޼O�gb��9YS�x:��hb�!����I��xc $`V`�8��N뛟Ct��^���F���g�F��hB���%4�k�a�E��rwe܍�;�24ƎI> �q��,,����Mbm8�BL����b$N��jiPS���7�}�v���M�掉 ΋� ^̃V��ѣ]yU��1�Z�?�wZ�����O"'i�\1g�GW:	��q���`\��zL��������A���|X\`��Mƾ1����}P]��5�@~��Z��_���c��y�w�&t�����Җϗq��7�=�;Z~M2]�tūB1����w������ 8X��f�;��
�R!�ReR��c(��ة"�f��9�HA�8�$�9�DO/c�8?΁�1g?�湘�90W��e��U�㢇��kSe��r�8��o.�(H�qp/p���s��~F����M��/=�a��0M����5
�02~��v��i�_�?�*�w���qqU�$G��d	�֢*KJ�S�	T�7|�p79}�i9c��<��o۶�%WX�h�W��Ç��a�cLh���W$��pPc��Wel��f��c R��	�	rl�Jg���9?+\���؆q��V7��"�!�{�ӱn��tU�O����ze���kyNM���&t�������dT�+.Y���iv[qj�5?+�V"�ٴ^A�x��� O������
i���Ɍo�2�O�81�	�<c�K�,q�����.qc<�e]7�� ��0�&�q���L}U��q{.dX�N��b<f��}�7��q1���{�9ằ�^U/���jR�;�g�zKT��Ӊʨ��h-w�� M���FL4�NW�L���2�UyU��Il$K*�Q8���{j��0�8>��A	�]Ԑ���/,
����Sw�*r�XU��j�c.���{����5p����񙉮6��˛�u�?kױ�5���u3���=5����\(!�Z��an���X\x0��N�D��B�m�i]C��Є�Q0����)9��s��k�{�wg�za�bdƸZ[̈́-֠��$��@�p�c;ڦ�0�Q�o��}A؈�8p�=7��c�+V�h~��9,\�%K�ذǳ]�de���2$\;�QEef�R���\�P�ݽ�����j�R&r��<9-sz?0����x��{~�>��3�υ@o�*���Z}&�����ޠ	]�`H���i������=~��U���κp�b�]u�����c�1߷o���B ��:��H\�~��q7��sQPf���9"d�U���j��nm�s1��V3���L+��w�H��,��)ê�pĄ7��R=.��k��9O�?�Å=8'9,��ܘ(�㩰GW���_Mp�������O�-���F�	]�`0L�j]�.	(1t@m��Y��\yk���̞�UJ�.3��Fb� �)S��D�Zk�%S� ؈�hX �Z�[��c�S��I�Tkù0?$Eb�f2��G�η���q?���[��=�0v�Ni j�������w��996��SY._����W��]-"]����[hB�(,�s9��'cɧˊ���6�6��iE2NKw5�M֝�z�$+j��N9�ǲ֚�4]�p�#k��h�0jX�N�:γ{�n�XvHS�љ1N���-s���i�03�1o�=�u��0��&��1p1��Ό{4�	P2��f����,�!��2`�����&s�� M��m�֖�#�����nU�!9���	bd]6��Y7��iy��@� #�9���=	�.|*Ǳ��06\��դ;6B�18~���9W9@˙$Ͳ8&őPi��
����^ �#fOmvj��~0��.wzg�6�K�⹸`�6�ƨ]�p��F533֯���i�t�j�_m�kh�hB�(L�pTK�2L��wÂ|<�9�C��d�X--]�XQ���8/K�Tw����8�`h��܌IcLʤ�VD�x;��x�2�����"��j�SuMULSC	\��X�����q^<# R��l���!խN���]��P �1X���|�|k��U���	^-gSA�:�?M��-���D㼽��
��	W���$lhhT� ���$-N����K�Xj�8��@�lnºsX���ܰ�1��p,�v.h�b̋V3�����$<�ک�봬�&�r���)�uЫ��1�t����Rh�s~>T�c��#��abEl�L�,w�?u��S�;��:ā�\�ń���P�	]�`�|�p�k%A��F�~��]% 6!	��I� 1vb�[�����Q����~UU��P��P���X�B&�b;�B#9bƯY�F2d����WqM8c��z��ǐ�ڝL�I��Vg��U>�,�8�z^����3,d�P�9��`6;��9.-t�2 ��U7{~����v��]C�@�F��X����ֶ�А�~����֩J`��E�W��uc�r��y��Ǽ��2���""E�޴RI��F��ʦ�:�SZ� �� S���8G���5��*i�Ms>t��X�x����p ۴ғ@w;�Kbgi[&��x���j�Y��zrz�`�9^+-o���W���1�pFu��ܯ�b��u���0L+?�^A�F�Em��-���jV(Lw�r&��򾖩,Ů���G�^2����ϳ^CO�%�L��TZ�kF�w[���)ZO��`X�bA���s[s�f�3���i�Ϧ�֫� ��u�S��ڳ�=B/**κ��r��upr$
�űt��X\��P��b�>�%���Z�$j�νLv���r�H6��r�h����{����[��$���x�{_��m ��[��"3�d<yor�vr������;v.Ӟaw�"���{��)�I��>o�bfDVl��̻sL����审�{hB�(������#��.��`w!..,�5:�˪��k	'S�*_���`	O�D�"'�������CAtz�H�%C����,{ƨ�uN��-cǴ�i�2��Fz�ë�� �VY.��0��>j�3T�c U
۱�`t���(��n@���w��t"���y_2٩�X4ǧk���Ԉ��|�ѽ�������v��?;��tw�˯p�y�	]C��Є�Q0D������j��z�;_{.c_.~�$��D�۰<p��
�O9�&�d-	�K����⺒�D�I��۩��w��PɊ�b���|&\R����T�+��9�G�]����%Iw�73���n�5/�If19?�L�qPӞt�s��򦻭�+)(��{Ȝ�+������lxiq����ܖ��Ϥ;���]�@ҪZ�q��1\k<+p�J�����z���D.	�gݶY��.��P�H��F/�	]�`��lRZ]�\�,4�r�ƪ��J��5����X�Fw'3W�d��,o�X"mg�IY:�I+4/�K�ȑvg�#W�͸8k�)wJ�`>�زZ�֑�5��F�8� :;.)B�h��3��q� w/�=������4(��'���fw׈{aV|��ʅI��D����\{T�eiL�C������[ �t0��&�-F�n{�ke�g�tf��F/�	]�`�đ��Ι���Zj�2�$J�u�gEL<R�C�#���#��)N�Uo$a�7��)iP��� �D���$)I��D�uOâ���l7�~ ^,M_D�}�r��ߖ�sOM�vp��(��q��R6A���"ؒt�;-�����%G�N�5��q��2r�t�#ޔ��/+�2ǂ��g,=�b �J��]�Óo�{���d-{!�\׿7�2�}&Do������e�{�,p���x6,ѕ������9n��~��j]���o���s���?>JC���Z�]C��Є�Q0D��N���vcͰf���\=�*8�d���-r��Z���tV��'��P�|D+��r}��%pK~ ��Ju�p'ǈ�j�a�R�E��=���׋�[�����%_p��(�nd�ڝ���GꘈD���VO>VuK�<YZ���~�����dx�v���B���1�Tڋ�������'��/2�X=tH�,g�@�j���ַ�*��U���Y�ֽ�8�N��e44zM�C(�?��1�pUP�sE��K���=ݵ&����:dy���g@gҚMJ�Ii	�}����J{��$EyZ��$jd�I����l�<ޢ��%6����OeI�p��J)]����	{t9�UMw>�foqb�VIޡp@N�]$��.sL���]C�'�r3��zO��9�������ae=f�[����Ϭ�t��%��vO���I�Vt8*�ZZs����Igs���6K�xnR]!;K����{4��z�ߝ���Y�B�z�4���}�Q�t��SBCC�WЄ�Q0�Beq���@�N�`%ò���s��xi�z$���t�`dr���621�q�'oq,ILȒ;& ��֟�=l���c1�n�f��6YϭƁ)9��qgz��9@��ea�w}I�ˇ�L�s��ȕ���@��)���sY� A�������O��rLJ��
P��Ǹ%��{L)Z��  vd�c>�`q���x9�+�Z��,]S��9X���a�I9�!���'���F��	]�`=zt��!CV����v�2I@���H�A���l�t&��-���f>+�r�"`ܲ4$g����@$,��n�?����.��%㍹D9�s{<G6*a{��YU���컉�+_�tc���|)�&�*x|N'�r��i#'ĒN�E����1�T���niۻ����)��ML�H>��{[kK��fw�yOl&�Zͨm�{��G�t�^�Iw_U0��ݱH /#�������]P�z��=7���k���:�����E��YG�¢Ehhh�
��5
����Ĝ9��=��C����.mmm�x.h�-��zn�J�����U{��5�G��FDc[�ky�$iw��}Ғu�n�޵��1k˳Pͬ��p��7���8I��
�X�x�	�x.z�:N��}@~�0.N��L�\�nV9<�p�'D��u����m+Bj����B	=����Ζ��cv?+�����j��W���.�@����,��E��|}�9���`��<�\��ñcǚ���y����BCC�WЄ�Q0^���G����e�6���]��/	�C�`0dJ"0�W4�ơH�ZƦ��d{�qi����J�D��SnR�_�{KK��B�Ҍ�@M�-k�I�H:h����dkׅp��8|FZ���>Caa�'���n6
�@�x6���������H&��b���4F����q����w��=��\7��f	�u�;.���Z�݋�a�ŐaC�O��.I�vZX��Չ��d8TP�= @.�:R	̊�x�:n};B-��,��.�����(�sکT�!Vy����,�={�v�kh���5

��noذ���״r����\���0.ѕ(���֙� �_���w�;�ɕ<�T���1^IK)z=��( c�/R�󝭻N F�X.���N&��$x�M�OK��X�O>JӒ�����.b'�M�^�FO&W�s[�oH����@+�]���b���+���l�����R@��e��s�g���{� ��"��{���a�U�s`���,r��l�����Bw�Ö�	;�m�������X,&WQFsKk��3f\��k����P�	�
M��������.\������L&^���6���q�c���7Tf��~��=/s�LL�\ �a��w��3^�[2��XU^���
��--�B��$��t�nI&��L*��9�{G�<V��V�	��ts㩎��וJ�2����)0dZZ���q<���w��Js�q��iO�� an��kٚ.�ʅBgg�%AD��> O�+ ����#md�4�wY��ُ�;8�팓�����l�h������������{y�X����I��>���mK�gSN�rE܄�x�튯;r=d��Z~�_qq���~/3r�`Z���η�_mG��3�L�2���K^�!o����N�x��f��|>�3��ҩڲ��÷|�G���o� yRh|�����0�qF�	]�#Â�NţU��?"���������;wn,9z�X�����vRQ�8�$>�d#�l˴�+���5�>��%�
F]Wp{[<�E�oU�o��E}��>�LdS��!��LYYq�z��e-�H8�!�J���YV:�	;)W�#-MCR�/��<�v]�Ҿ���w->��m��
�3)wf�e�e��v����ؖ<�+�e�}9'I�A;$��fж}��y�t��<��;6�)�K��L��Fʴ��r��m�������=�aD˓8����{�KN=�H����V2�4������6���O���\�gϞ��D"��7��k3�``祗\��#F�H�T�ݙNY+ct9�NёN&}�pI����#i��N�.�^^n��&�%��L���L�v~�3���w�����u�����@�(%��Ѥ~f�	]�@ֵ�J��G�|4��8X�_��p�9>�_0��n�t��ӟIf����������?�K.̖�=����N����,�;����k�Mi��C�c��맞j�ut��ۑ�WYY�:u�n�׾q��[n���s�/�O���8q�ĸ={v|������n����(4�4�k|�2��7�fצ�֌�7��;D�Z>�;Z_?���լ�g��?r䤸�x_X�x�u�6\��&#��w@��7�Mhh�euu'n2t�������ǋ�&�3
M�{\|�읯�����?$���DƱLi��+_�¿|��{�}�V#G&��{��/�<�����ZZZDGG'J���ƺY�f�4hP���P {��j\0�z��P0��Y]=�Nh�QhB���c⌛g_��S'�o�٧�xLcK�Y
	#��]V2n�S�����ġC��6L��{��}���ͻyN(��:d���jWWWҲ����}:.������c�w���W�G�>g���&L���|K��;�Є��$�t�K/-��7�/*�E��W��|�^�Ϩkk�f��uO���t�|t�굃g���N������BZ�!��go�ž�s��\�m��&44���c��?���)�g�Y������}�ڢ~g��5>�w���?��CO��EC��;!�E55FiQ�Q+��"��|���j�~�ؿ�������CS>-4��v�*y��E***�B!��(Y�F�H\�q�5׬n����,���?����䍑H��������=
�jſ@��'����<���_mY��Ё����8�H_{�Q%�PqU�o>R����u�[;�,�����~����r�'�xzJMͱ�C�	C��j���߿���W�p�G�եA�����]�P_7�o��o*/^���N��.W+4�k|b��w��������7,z�uTeټdM]I�
!aɴ8�1��4�n{�����Ƴ/���\5���:�F�7*��g�����t�i�2��j��b醆�]��~��ӧO��L���۶m�p�k���_�r�˯�|x�ԩ�4h�Z �pЄ��BV/~KW��';^X1�����MU%���.146�|"Z.�)Gkk���{�;��{v���>7e�]���ǋ�������#G�^?lذ($\��ʯ�`�E����n�m���
����h��_�<y�M�6�VV�y��i3����t�J�	]��ߺ�l{��o�q��O��+��O�B ��)��������p*y]ݺ��x��k�<�ԟ�,yf��+���1R�S��k�~䑇��~���۶��9����_�x<���[o}jڴi��\Å�����+.�ٴLߞ�o>����կC��SB��Є��D�R?<�܉�Y��������]c*��?u�6Ȥ���2��0"�����7��-y�＾rƌ����i�ҍ��g�~�T�P?|�w�L��3+*���N��e��*�C�y�_��V�����/ھc�g��/��]���o�����F��	]��,��:6<��O~�e۲Wo�./�!j8�O�jD}�Q�D8�1�����M$���w�\�qي�ο⪗�/]�F�ٳ�?�.Y�d�/�p���$Fmm��-���<u�رM��s�s�&i�=����~��_��կ�ݘ���-]p�TW��l�
����5>�0�OO9����~3����}��5������$Se��V#%���8F��2��=����y��5�>�Ƅ�����s��u�M����A������;'�10�V����v"��;v����;��o}Khh ����������w�����z|�؉+����A�Ƨ�1C͎������^�nA}͉k����J%c�	�)}BQёL��T������9�9���+.����ˆN����'zc��_l�$Z ˖-�t��[�V����:O�Sޗx}��7$�?=n�8m�k�ޜL��=y�5W_[q���%�Ϟ�XIQ��j��	]�S���$����O=��/<�p�u��D.(+
�Htv��[[̐i�J��m�����S�߸y�O7m�t��X����n���N|R���ѣ�;��@�?����"2(U�D"v{{�[]t�cw�}w��'� ��������3f^8�0�C�/��ᾱ��B�#�&t�O��tJ�k�~���<���m��}vP�xFQY� 3m���im呈�:�՘L�Ă��U��95�7\���VV�v<������Ǚ�am��'?�q���:�8�N�u���U�-�?�=�,׉p \�<�������%i�����ٗ^�T/�>zhB���"KPu�ҥ/�ݳe��g��zd�7KF�T&�E!3���d��!�7]�mF:;�Ŗ?ܕ��msʏ���]~��m�<�}���8���߿�����h4ZmItuu�ֹ�3�J%�Κ5��s�6�O=$�[ZZ�K2���{�\�b�9s.{����Yh|�Є��1Ǎ�v��Gw��ؚ��?s�ɝ��hK%/-	G�ӊ���)lGD̀gRf:c��C�1�Ȑ���N��׿������u��_�x��k?.;���}�{�n�z͸q�S������f����4Hr�3��?�-���ʕ+��m�v^mm��'O�|iQQI��s�.1b�a�9;�	]C#�X �:!-���ٳ��%�M:�}�M�T��`���0"vg��[F4m�F(��Q��Nm�8�w�7^5�чmY���I��;ۉ�������!C�Ge2���9�d����us�����;ݧǏ��r�-y�ĉ{����924t�Н_��W�˷��YM�y�Z�'%�/�ľu��%S�ڸ��t���HhH���XZ�V,Ŗ-"�0��PI(8�*`T�[�rڃ{��2�e�N�]������NS�u��c�9rͰa�b�mh�k+7���E�������\h|z���c�=6�СC����WTT�%�����t�M��c�g	4�kh�r��,|y�/�_��O��8�{��@��X 2:�N��VQ `�A�=�4��TdR�xDcGW�7�z��m������[�g�1x�Ye��:���έ���v(���;�;��k_��ks����v�|��k2��9��/))o���#�+��+&4�hB���3Ⱥ�$�i|�z�+n�qY�J]��3N����e�S�F��7�ә��X��c55�<��]��,:��3��b^�8K���?0��ɓW�7������uw{ �:�z�3t��X�zu�U�V�<xp�����h�k˅_S,;+�O�VhB���%�e9��ؗn{��uk�<�䑍k��u&���Ǆ}�����όw�)�~�U���b��m����q��_��/��u�vc̘���ɾ}���������S9FZ�n�G�D"���5�w-��y(4>ŀ�������ikk�h���~I⢶��IH444����6m�$4�hB��x��{mZ���o�-����uE<i�J$����hy(dt�5��X�0����eO
�����A���Yxj���>��:~������9y���ES���njr�����5�\s\h|�9��^{m���C%%%F4����v���x��W�i)���54�'��:��_���7,}��gOx��ή[R�}�b�Ύ�Qd�"��`���Ԓج�kV�����wІG�ȴ���W�0�Οx��*++'X�e�����+**:��[��y�/�9R�qk�={�T�ܹ�D�����(��%��ܼ�nx]Z�:��,�&t�������n������|n��;�we2�V��*#��L!"K��m�	�e���j�⯾����k�gi�+dy�����^9jԨHgg��k�b�)..~eƌ���<6�7��ͩ���JⶤE�G�<�H$ޘ7oމ����g4�kh|H�&��Kb����}c�o6���,^�����ut��%�+����F�;K�����'�]�x�Q�9I��+���jI܃3�����]�b1ȼv54ԯ�ַ�񪎝k uuu��{n���H��d�tuu�����+���#��x;4�kh|������O=���߷k��;G�gg�}��q���Dt�5�c+������W��t4���l�m��(�?������p�vvv�ej�ڲC�p��qc_�ꪫtf����˗W9rd��ѣ}���F%D����$��P�C9�|��N|�	]C��l����/.�8��W��=���ܾűsN6�FT���t��b�?���N�`��l���DS��.��Ji�OB���F�T-�$��[�]w�]+Ǐ��z��/}i���R]]����<yґ���$�5s��=y�}����N��nêI�e'���߅�n�hB��8�0,���������}��5G���~�ґ'ZCQ�O�D��U�×-~�ᦡ�j��g�"y��ǫv�څ�b$7���Ñ�^WTT��7�P���BCCZ�m۶]YUU�ӧ���v���~ƌ&N�xFE����>�ɧ����O��e����Eߗ�u�ş�&t�3���}���Տ>rｩ����#�T'����N{�1�$V*�������W������9X\��r��/0-+�=z�p؞��;v�q��k�\�X�r%''�;6�4�V:�;gΜ��L���9����{�|�D�g/��B�sF<է��&��g�	]C�@<cF��r�S?��?��8��r��oF�!a$�V�eVv
������r��{��Kǖ-[V������o@,������F��y�n:�/��/BC:_�җƧR�a�:w�+ t۶[����O�<��Zʇ�9 V��Ϋ�:xp�w���Y%�|�B��Fa\|q��t����}��G��r_KL]�fX���?���CC�m����m�?�;>,��SO=7����@ ����&���3�G���ٗ����Ķm�"6l�P\\\
e��w���|GǍ�q���g̓��ymCM�[n�L٪�+Z&N���cB�WЄ��Q`s�t5-}j������'�Q���j�EDkөаhx�?t{����!w���F���9������#��s���v�Ċ+��}�׿��4<<x����v�9��2t���$q�ԩ-w�qǞ3�n��Ձ�y�͍���9������B�WЄ��� �G_}���ﯟ���#]%��5�O�>F0�*�k:5o���"�w�U�{h��>�W><��������zb�ĉ+�ϟ�"44�k!�����\��VVV�3M�j�n����y���{�g��֣�>py[{�5Gd�M��je���B��Є���a�e7���]�x�7�WN��sU�!�om:)|e�V�px�[[�߾����%w=�~ϱo߾�����***�766����p�v����WZzV��śo�޲e˜P(�߿���=�e��J�+�v�����g��kV}q֬Y��E�˦_p!b�:��	]C�#���ѣ��X�t��퓊¡���$�1��Eẖ��<��TI��߯�sÆ;w�l萡�---��k'4I쵻����$���1j�����R��� w{2�o���j^x�3r^�,Z􇫪���F������^�W���xOЄ����<���g���W�63\Z���l��;S"��aU��o\���['wmx?�/z��}��E]]]~$7�R)QYY�nmm�3o޼5������`Ŋ�K�|ҠA��d2)���Eggg�\���={�����y��g>w�uו�=�y���/��g��I�&t��U��=5z��/ԭ^=��8'ٞ�@RDD2Mdf�y��}�ҥKC_��q�P���j�:o�Ѫ�s���~ 44 ��Κ5kRqqqeyy�@K]i�ے���5j�i�Έ�?��6o~㼉'�+���!��8���{}�Є������־���+��/�ņ���?��)|���8�q˥GW�ޅ:�ގ��o|��::����P&�F�ɤ�^z�/_p��BC#�իW��ݻwvEE�_.�*"R�TW<�:gΜ�g�`[ZZJ7n|�V��/[�����>�3��4�kh���`h�ЩS��7n�"u*R�Z�H�e�/�֩Ɖo���X��kB߹s�����_
�`����e8˲:����/~��\C����{�,�'#����C�ySS�#	�M~o6���gD�
�kW-��ɤ.�,#s�%3�9|�&��	]C�,�a�L\�p���7o+	/1-ӗ��?x_�N�߹y�x�[]o�[�|y���3��V�%	tۓ�䉑#G.���u�����ƍ��ߓ`UU���_CC����vx�����TK���_��C��۩�M-����z�����Z��}B���Y�a�&���.Q�x~ 䋥�&w��O$4hώ� ��[��s���F#�5��=.������?��lԥj*�m�V�iӦ��;8p z��=�žgҤIo���k�9�6��C�\|�y�Mlio骨�x]��c�Q�c����54���1hܘ�+�/�F9���SIa��a&ǜx��������^�:|�[g����*7��l��cYVS$Y)�--���k֬���2z�����:�v���8q��|��xc󪱣F��n��塡Ç����[�1���l� Є��q� V�G��q`�ں�hxd��Sn�Eб|�����7�D/}��'j�=jT4��� %�ũ�������yܸq�TM#��m��6���@v; �7Nkkksee�����3�no)ݾi�M�e�}}��m_�9�)!�w�M�g��;��3hN�<�B&�0�Qê>�o_��[�nnwHw��4~R��}�I�< �v�C���V^y啺H#��۷���^4`� �����l�=�=z��;~�D�e�_5lؐ��[������O�;��EB�љ���54�"��VwE�*�e����L��E-h��?�?vd�ظq���-�x���o];��ᕨ#�,d+�?�/�x�ZJS��,YR$	|ڐ!C,�[�:u
	�ɮ��]�f�:���h�^��/=y�'����&����-so����z����	]C�lBuu���5G�A��b0�;����m��h�Ļ��O>Y/J�S!�ygg���b]���ϛ7o�����?�я�Ʌ�4c�t<C�<!�7[/��W������?�p�%^8��؉䅗N]��Ե��<���C�&t���R^��}'ww�~���O[f�vD@�0v*U�pL�P� �	e�;�kJQQ��t*m��.aKb?YQQ��\�'7i|��[�|����K���o���@�ő���A��?~����u��)�ֆU��|a�Ҋ�H�.���G��6��@���Y���~�]�q$��k����#L����%'����q/��rYG<~eqqQ,
������4y�d��[n���ӧ�d8�8q����#%���*5K�P��;vl��+>�9��K}/��ê�b���_L���+�nKξ�Z9xK�a���чM�g��i����L8�,C$;;E8��m���ڈܥ1�$�M�2e��gM��j�[�ٜ�����w�}��?����P!��A��N�3vL��~B��hnlJw�w�袋���W��@�#f���~u��g������E��D�?���6��'�����C�&t��vii�����^�p���F��$���Ɩ����C��8v켊>}��e@�;�����)S���ֹ��k׮��tr\yy���=H��$�UZVvh	�t��U�"^{��i^2�_EE݉��Y"hZ����?Ͽ��*�(���4�kh�e'��`[&�I�O�e�"#�!n8�����[n�eR2��tg��h�*	=��Լz���^}�U�������nf$�!���S�T|��ۦM�����H�{���86l��VXfi�d���qѯ��]���.��3")�i�&t��ɤc��.;���e��D(��5����u�b��n����x���M4b��|���[��R�0kH�mضm[h��C����D���&,�D2�6u�Խ��A�?|xYp�U+C�sDk���E{�]�	�"�O��|������[h|8Є��q���4�N�H�>�H��3���d2���,��o}�[#Z�[.������~�si������_q��k��]�t8r�H���~�9�㗄.jkk�}J�S����{��pxٖ~Cʊ�J�ǎ1a����(�[�:�չ���o\�A=�	]C�lC:�|���Jf,�_�Cؒ�}�i��iKݵ��&���'��B���/���������c�Wϝ;��������P���w����x|`�>}���@v{"�HE�b�g̘�4Ց�������������"��*ʫ�:{��N��0��W�xD�����54�6$�/�d�'h��T�Bw���4�]�,Y2d��}׌8gDT��6�e:j'M��a����0��'��k׎�D�!��?��|�O�>m�a�>���a��U�;v^[љl���Ũ�-v:Q��+o��������ˇM�g!L��A)�pg��HZw�\�.4�o���I%%%c|>���9H]Z��#Gk�����r����Ç��{�����*r��vt�:ۮ�<~�[/�����vk~�o��tƸsC�t�͞O��d2yl��3�tC�v�k���54�B���Z.A���me�
�����}^}���6�+.*..++s�,tV���QQ^���ˮ=v��Ohh�c۶m%�d������'O���P(�քsG�@�o�^�b��WL�?�"��i�}>EE��J58�uso�y�a�ѱ�3 M�g!P���wIi%b��w�x1�{����SM��D&<����e744�L?���ӦM��v��b�֭U�"�t�C�\"��5������9��O����/VZ)N'DS�)�.�9�B4TO9�O�������&t���T�',tXP�dRt$��t	�ĉ�ŋ�4���*))1�2žr?i�8��^�n��XKj"�JԬ���OX�t�ՖH�����K��ӴDX�I;˴��`:Zh�)��ɈX�%%1hPJgR�6l(�ߝs (�ɔr!�y�������ן�����_��4�U[Nc��L�E�g���-_���7���xghB��8���o�?{��y�������l�EZ�����
0�`�m�1�%��K��vbǉc�qM�8�%�%�L3 0BHB���Zi��Ζٙ;���{�).�g~ϣGh��������/B�7�aK�uj<��l\������ݞ'S*����B���6�}��ٳ��,`�iǑ#�#��hT1��g�w�4�8�^XgN�hc*1&�Q��e�(�P�p.� �5B8��d8M`��D\�ʕA�J��r�;W^��Y�AK^�_�k
�*s� �VQ9!�g���A.Y��Ƌ9?T��hT�\�e��'***�Fi��;o~��B_oעJ�Y��i�B 3�7N�4%%�����w�(�""�6�A$
��	$ArÑ���n�q*/���{��.?��9Ǽ���C��t��.�ux�a��٩yw��,z`(������X1�N�%��QR����R�ep�aJ�!%�H
o��0I�d�B���8��e)�Ls�H��fRG���X'���DQ�DJ�R�ڠP۲�����-[���E�����<���8�ƧX�V�w� �	���\�;nl�7��9~\��uS,8>Ƣ��	�"���qG���^P6��οCDA���@#("T|�p���t<a1Z��cӱ�e��+H��{<#��x��e�����&��q�؋S������e?|�/J�^_-�L�5f���*����T�)�R��$�c�lg�,|�Y������r�#�Yn��� 7��C1Ǣj�\	&�E�x%�f2��d��?���;4D�o��ܴ�??\XU�o-�����|
�����nk��!���^���Sv���oo>z���zb��%�$���pݾ!�i�����w"��u�]"
���(�n$�\��\��%,�7�;��Wz<�bKa�Dx]x/fBu�pYUŶ9s�Da���H�o�H��/V�h�?�q�$�k��m�:�T���HT29B����fSI`���Xb�$�OU����4��r8���:Bz�ȕ�e_�y����A�@	�)��� RJ
���%"�aX.�b8_(\8��=��딯���}r���x������\G�0/�1~{� ��-]�t,��~@���g$>�$�-Y�ӧO�F��v�z���6�<�@��T��t�
%K#�E�|!���Q�EDF�$�f�4oBY� �Ng���/ U��g�'�[�y/�X,�H� �KAO�:���_>�A`\K�u�f��m��xiu��_g��Z��Ve�H
S�`,��I�&���@<ʟK�̈�������Eq	���ay&�9�+,��$M#�,��>��"�*���\X����Y�0��B�>�� 
�BL��&	2c�"#lF�x�<�i��|�r�'�hr�jf�޼��G��p(�j�I��#-��Ҽ�͘���Z��ev����R�X��,�P���!��ɓ�����󭷬m{��?7;+G���d�s� �te���M�}Jt��=�����B���0A�2#u�I�I!5�8�.tf���g��92�ID#y�{�՝�`8�a�l��G,O߹����1�L�uy$�]RR$7ʕ�RB"l"t0 C� ��K�(G�<�I�@H���#�d"��'R(�J�L�ט����:y<�U����z��i^�y�qL��t'%��@�/ըe��7��!u�F�=�H� (�ʑ�z\J�j[6�e͸72z�A]���س�/n7[��.��3�{�������V��()dg�x
�{_y啾���P^^^�f��F��߶m�<�fY�V� ����?⢉x��i�N~�2��B<���yJEmI*��[!��j�3Iw.��pTV�U�DAm$�O�°��q:�A"�D�Q�*�N#6�����)Pi��j��m�㴦0�ٹA�wæ����sadhp�Cs��:M�9�0�)@��#a� �]/o��1�1,�'�,ǿ
�H��O%�,�;H���`)�jmF�֔W�d16JʡF���"�}Y����^Gb�S���0J��DtاbS�.�������]�D�Qn%��%phs�A-�
S�������\&3��
?̐9=Y�ۓ�?)/Ə)�Z�}�/�[8OO� ��ؔ��P6�Jǥ2�����9?����O?l)S~����� g<Pq���ٙLf��aM�����4�z��ҤI��d��6���ϝm�6*0u�����" mA�Ƃ�5�g{
�ق(�""�� ��a��d�=���y�-�uZp�|��6Mq	���-[�������|���ׯ�����ދ�~w���֔��l5��$H�q�>�E�@g.�f8��	�� �q�!N�7�\{ܖ��>��̝k���'ONBw7+Wr�F�*�םN"60�j����W^*q��0[t:4�w�f�^��x$���x<h0��(yQ�2gA��
Z�	|~hki�(`U%Œʹ����?G�����\ɤ�G�M�N4W74���~�%��y��oٲe����F�1v&�����Y����dTA��$��qH<ǖsL_S���D��r�*�Ԫx˟�' �4�l���'N���X>'"������B$�.��R�q,`j5�y)��ASZq�w�?��:���UW��>}���4N���.Z5�}���z���1KvQ�</ˆR��#��@���h��GP�Tz�I��L;��3���_Ք]U(_�������u������U<|�tώ�����p�b�B�8�~84���j��f�S��Jx'�}�a����Y6�J�P�e���R�p�B{w'DX�J �H@{��,&0de!q)���j����qx�S���//�:fϞ�}�En���m�����S�w��)���MQ2^{	$͋9�r�@0:���=��gw�>{[�h8�t��^��҈7 J�/&�)�e��eub?��Q�EDF!(�g8��2���������j9�y�.D&#��dx���/<�]=8G޹i��ͫ��~j���P|�x�&'נ��[�(��C/p-�!Hs�N�)aနy���nۛ]6��'�:�e���[��'�����tbϑ#�z,���U-��8����Z�m5+�L�,&#��R�I��E=��S� t�}q0�$�UZ��l�p��R�h�rp|��/��m�"��2<� t�z�P�{q!���S@�� ���l0�E����"XTL����_n(޼g�����|������^~��D˳����<���L4�5k��SO=���'�#�y��c�Iz�� (*��`2�Fu�I���uWm����8N��#
���(���$�d���`����a �� �w$�z`���s�N�2e�t��v��{����)�>Y�����4�ʲi�ш`l��}��q8��!SD^� ���9�e����p�n�8�e�������Mz��q域~:˖MK�=V����
������6Y��+�Q��_/8��=w����k��@���HI��P���O��u���"��N��$����A��<����C��H[8����
(M&a����q�2J9PFd��b���$'?O���3�PCØ��ٸx���������.��A�e�WO��U"��PA�[�������b:PVV������(��ؽ����]�rX<L.���/��_L\���Xv��Et�цT� �D��,��α��>HS8��V` �d:r��q���+/��������K����A�?�PU���&���s0IVUy�"G�A(����N��	��dT&������.�Eus>�\��he�� R[{ZӸa�z�e���ba}}}U����G��"@��\{�|��ZL�TMm��Ns�8�_�p0�xT(M#��eq͠ri��S!`XW�C�)��Km�u��A���5��y�w�ۺ�4�c��IEӘH2%o��Ĳ|A(�����R(�M@�c 4��z�,h���'�!�IB[��v4��f�-'�N����)��Ȅ��;s�v��W��_Ͻ�{�n�ߗ�p����[d2�H�?�r����Y������?>#��p�8#������e������s^�홱l�'0nFD�WDA�dPL��0H�_R�
:��A�w�v�:���p@��I�^spɅ�{O��y��Ws>{�����V�Ke�&��弐�2	
�` :���E S������S���q�Em�����<�SȂ�9rDu��wVlظaawO�`٪<{�������������k���P4<��&D�+�2VBI8:�xQ	�a���N�_Q�\Z0f�>vl\hL������yW�ݽbϞ�ˏo�z�6���m+��dіV$�b���*+���7��Pȋ�u�,�~�����N'a(��s̹��_:�:e�ӡ��]K��c��|��>�2���;ݭ�����ഢ�BRp�n����A��@e��֯��ݻWѰm��s-��d2�$��*��L&��ygͲ�G����Q�EDF!1��H��Z5�b�
E k�8^�3材F��<nߢ�m�>���	�б�V�+��0���-�����uBnfU��@�'�{!G9&HH�L�9��l��tͦ9�V����;r|�΍�U�.�ڵ�E�`�&"���\Y\P��Z4I���tBOOψxc#�r1��I��p)�L�f��V�9��tWٸ���q5�	&�y����e��/��=��|1s��m��~��pS�E&�^�R���	�/��r�0� �r)��vO�yU`�����c(���h����BMu�k�H)�̾��޵�]�����~_�7R�'�[�jU6�r�R����hkk��Kk:�̙3{���޸��1f]b&��&�"��X����ӽ3g~*�����Q�EDF!j��quvq���o�~H��
5�#q���`rd��%�:��@_z����_����[\ �啚��Xk"�:;a��4E�~�u��T��Oj,�0�������1��cp:"��yg�fŲeU�Z���TuΤ�ɲ�q�аfx�'ZZ!����A&���t���H���DV�uM��&^��UUUy&O�L�jn_:N7l�;_z�Ğ���i>vE��:b	����G�����t�c�S-֑��P�9�C�w�=�9p��ß6u2��iuG�]zӭ7g�<u�1~?[�}~�,��{eG�6�U(J������ ��X��	;����VZYh�g��#��%��	:����hZN휲��#����At��F9o�x��KY�B��2k��~'�(�#�=�~h���߸�+?x���uk߶�Z�UO��R�۲��D<n7�t� �N�iJJ���÷�_yɺ��\s�NM|�|ú���_���r,7�b��fL�Ne�sx1
 ǎ6���0y!G��d�r9Ͳl0�5�5��E�l�5wn�����6�-y:���wr���߿�����j%��lVK���W�D��	���`%)8����XT�.��{w�����-):�T����F=2}�,�8�(��Z�NN}��?އ����o[�������}u�e�^��[P�Ιd2隷`ޡ�3��>>����)�kq��������L\���Vv�����}� ;�Ӄ(�""��r.���6מ>��q�\^�C�Tt*�?��\{�;���o���_�f�����*"��&A�*m6�<;�-�̆a^0Y�<�G�=Q�W4}ګW��f�j���w�F�i�&å_Z]�c�j�c&���TTTF���"t��	��w��[	y����L:�H���2���kk�V,>�~ҬY�����w]v��c��n���4���;Z�/��̍��zg�M��`/)��r�>�}}�d2�o�������?���s0��T�7Cʹ�`Ш�	�UH{{G��|���plH����k}���.��Q2I�(A#��W��{�f�����nR6�Wj���J4���A��hF��5�%��ȟA�� 
����#MzG:C�]�ʲ �Pk��KC	�A�k���O|���(���������sPc�˵%�y�I����a�wB*ò�Znu�[��ޙ���O+�\7�9��ب��'�MY����c�����<˘1c���\D�$�����iZ(S��Z������[�Y�h�\��L�}߁X_^� �m}�W������"\�J'��Gb)�m�@r���ɓ�xg8<~d�K���Y���i����x��5'{�V(zs��xՔI�������~̓y�a&�<�o��o�T��mss�,�Ng�0"�$q�����VWWG��F�A���V��̭(�U'�A$��Ӳ]�XO��SL[ ���ADA}p�ee����^�CAv�H+Q�����qݎ�������������bz��[��8ڸ��l���TeA� �'OB�NqI\����s����Y�.�ɯK�eןޓ�Z�x�����z]W��.�(�h|U5����J0N��Ak�	�xi�%D� �h�N �m��9;�.����5�=Ep������9�����嗝M�k�T�L�aՁ'������]oF�8v���_�t��ˮx�Ňy�^�oٵ�T!/p���C�0�N�*�@)R6�矻I.����o�:��;����t<6Oe2
����ȱ&���~��mڤ=�����9�"�B��zܐ�	�L:����_t
����=[]Dd���T
-M�D����� G���i���%K�|��g��9���S������Q�w���Rj�`�,6p�αoxH�cC ��X��}�u˯Z���K���:��m�����/v�Z���͙-+(�Gө�9��50^�0'%�� ~��X~Q��_q�橳g������!�e0j��:y����lYw�y����d�	������J	�&Ta]��_{㾒E��}�W�����<�ܝ��x*%�'M�rBF�#��g�z�N�Z� ����z<G���m�t.?0�FP��,B@M�����m���ί�-!���_5^'%����R��������~��=G�;?È�."2�@��V�ӫ.//������� �S�Ək�5���n��� ߹�����x�f��3F�WUX�P�Jm��#CR_�q�d�E�\���oF�j� kN�I	����U~�m�U�����Qzaaaa֔ډ�B�B�����r	S�\&�Ii����i˳�?X���XS���ZS����_��w^��s{�xc�cѵ9Y���'�Is����a�قJ0�dg��7;{{��ߴ�9�=����?��T��4�!L��3�O'�nݺ���z����.���+�̴���'��:�L!�d2)�9��Cs��vUVV~�b2����m۹�����,�M���K:7�0	Fk�s�9˚���3�(�""��@  ���O��eJ�^g�t��� �7-���z���+�qG�O����m�m��8��,G-��B:�żI������%�]�ӵ��.�_?pZ�IH�{�Wz�+�[�W����gϕ[MFd`` �Z�@X/Zy�,3�����O.Y}�����3��_���/����{���	�����t3�|!�M�`2ja�=[BX��M��}���5w��'D*��}O?�(���;�\��X�sf�6o�t��7��Z�S�i���/��Y��ɕ�@� )ÐNg%v/����μp--�S?���"�bn�N�f1$�32i�+�~΅�99㈂."2�8r�@A�ɮ��E"%���
�A�I�ޤ�䘳����V)�y�4=��g��[�/���5&��K�mY�ݕ���1Q��ݗ�?�]���s/�� R[��J��;W~��I�7�0��w߽���)S�L���\�
���)�Rτ�����f4�^]sٚ}k���)*Z|��ǿ9�.���{6���_m�Z3c����pD�;e�Š�bA(Q4t��|��hϽe��~���^��D��9x �9`��yu�6l�p탷<��_׃��lذA�~��<�R����0�@2�2u�.[���U�a���Vo{�9�F�ͪ�"W?x�!�D��۷�͜�!���DAE�j�-7�4����/*F#�(BAPHe�&`��T:F��m m�]���O\�p8��h�6��X��N�z9D&Mz1�
Q�kk���;EkָN�T���_}��1�>��*^�W��z{MM�T�Ղ�烡�!�y��T*�&S�.^��[�l���/>�dɒ�}�=?����߱�W���}��G�Z�x"���r����P�eD.Wmm8��G�ȿ�Ƶ]�U'�{]��e�����e+@i�ûr
'�bߕ��w�����?ڟ�p�5�T��M&$$�x�c6ӳ��s닊��R�#�� ��m7-��i�egS(ˁ?��L�:á���S����AdT 
���(���]�g��s�-.�(�I{xW�J*��@GRdp`PB���҅Ԣ��_,x��'�ʃ��j�"��1Y����I���H�{��<�����}�H!��N_t�0��B�[o�u�o�v�L�������l6Tsa����p8��e�	�[k'U�s��7^�|y�� ���ץ1+����7>LX3��,!��^4�L��l�e3g����+?{����V_B��ɛ�v@����/����f 3'OW�,,|��玾�s����h�����;v,W�`9�I�!�
�;�Uk�-]���Uf=����w��{�ΛW[�7kը�9 �X�`��e�d�����W��с(�""�a������q8���I�I��yU�(`Ba(�X@�;�xЯ�ߎ���Ƿ<��O_|��4{q�֤��ّ4���C��Q)8�z����3.8��e�]ބ�L�֥E��9l?����}�^�gϞ�L&S��j%���F~�x�A8'�0��:λ�u�����n�����������׿>�������8��	�%ǂ)��9�XsW�r��o���J؏������}
��9PV1�}��?���}�������[fUXj�붻&�����A�!�LFHy�b�X���ؖ�����U��v�|��r���L��f�/��O&�`�]u�z�<�+籋|���."2Jp�[�e��38�5+U*H&iH&�V� �!_��x0L��>5�ݡ�7B$�ۿ������o�R.-���c���G���LH��<��w��׾>��[��)�'���䧞|��p0�$''�h��%F�q�T+��9�W���~���3g<����u|2/
g�:�ץ�ꫝ7����o���h��4��R��DB���;uE�����68��6o?��7kv�3F�?�*;�p�?��S�����w��	�ǟ}z�R���	�bG:��4cHf�ʕ�O<����1r\���'k�HhIEy�ΪQB���7H����ުXpA��};]Dd���E{VSSS�R�!P�T2	��t6�RFO4.���k������(�^�k�篾q[�J�،"���^�|~�ҌA��3�����/�/�������5W\1�����\�P��\UĻr�eGڙ�A�P�>�ߡ��_��g?}��?���?����75���_��\?�+d��A�4��!/;���P�����\X���!'�?���[��-+�y|�Y����)S�_�fG����`x�BNQi�QKI��>33�hѢ�kjj�R4��Wg�ܱ{�D���*%q��v;0�&���y�؎�r�"���������������L��rQ�H�qPI��	��0'�XL�r^�b����\?�ʣ�O���G?)�i�Hqy��8RL萖R�b�`QX��/�}��Y��Y�E8���,[vmKK�*�Ŝ_TT����@HG�xw�!	I0�WY���߱���.x�m���d���ױq���}��n麱�d�1���!R`͂�c�BC�I�4h Q�����0�����3).)�z\=��M�}�����o����(�[X�P�?� �?J�C�/�䒦������H���rټ1f�ҤP ]�}�KD3��lϛ2�o��UU}DF]Dd��l����x�&Q�T�P�<�L�q@eX(���A�I$�!�����ёZ��oj�|��-cdҺb�\�?�a��q�?�ӽ�X������n��GȴӾ^����k%�����n��%y����\Lp�������%�/eX63���������_uYRQ���A��$����o?��d���\��s9}r.�Q�K
���jujZ5����{@g0�����.;x��%�~���d�w�tL��Ţ$S?�sq,��:i��y����hta�V�ȯ��}+r�r��j-�J$��u�V��z묕E����Q�EDFmmm��Sݓtz#�?T��d@�i�p�u:0�8pL�T5 �B���M�}d:���חȩiyj��T��=�h�:��w��G.��7����oՂ��@����Yz�/?��Ț��|Ey�ؑ@=!���`�ju���UUUo\z��^q��b����Ms��;��^�wi�qz���~9b7��4O�B]A�H7�t���[(�٬��~��_}Y�f2*��M�Q-DΫԀKP���]q��C_ŝ��m5ly��K'feO���&�=�G��J�~`��ϛ��:g��u�"
���FpE���c���U�8F@�N����$���|������H�1��Un|㝛z���0�4'�e�l��}�=8i��n��\}��ˮ��/�u�sh�I��n:���?�E��T��٥��084 �CN�U�����s�<��{n=ZZ:#r�W��?f�\lC���O��R��ú
�~rwW?&�uYT��C����+ ��(t��
9�YY�pa�����E�B�Q2R��\B %�B4���_�|�n��_��9|��e��DrN�U�ɳX���nf����ټh�em�l�"
��ș��ŮI
�܌"��6�	�K#��a �h�T?�	8�D�n�x�Y	Nh�Hav����z���LAG,�s]��#Hq�i�����Z��k�<tC^n�ђ�-�ɵ��r���a	����d�����a��~vO�( _���o���N��㾧T��;�¥���s�@*�e�5��c�>~F3L���]N|����P)��Dc�O����������&���}�����U��X,��~'�Ub ޱ��5�#ߠß���(�""g�#G�(����3����@,I �J�Y����r��� ��#̬��$���0��b�FO��_,���f^|���,������n��ƛ�����Jǘ
�
1RFB/,�`P�-O&�����]��Ɋ+�bZ��C�s���❿��	G~�MHK۝.�X)���J��� ɡ�p�X��~
���.,���15 ��rB�!����"{��>��B2������۹z�,���5j8|���n�u���K������ 2�]D��m׶�p0Te5Z�Y1�hJ ��5��L:å��x�%焜�8H��e�C�?���hL�?ٺ����y�=��<}��O�>���V��;~	���yA�������(+������_L�����O<q�XLi�� S������z���1t8�s= 9
o���PY\
GO��\��1F����6��/�19v�8u
�} ($�IN�R5�Xq����&~�kh���ͯf���u�e�M�A��J%97Ɔ1��?��A�{:�]D�"���W��)���PH�NU��f�+%��:2V� !��Q�!�Iǻ�N� %�h<�}����2sժ��-�O>��̇y�T:=��d����
�~/�:�@�fXO�;���U��؟�i;���OE9g�o�o�~��'K���*��oB�(b�Z���O��x�:�;�dS���������A�ւ��%B����+�w>�����~F*�=��bok��*�nl�F��Lz�z �r�/�:r�k>����T�Y�(�""g��M�<y�
�$�d:���\��k4���}��ﾄa�R�H"���Db���0��C� b~�\�|����wQ�S�ɇ�p��?�;�e��UWKKJ��w���B��t<�t����w�s�Kk��1,�����"��ȯ�����$)%/c��*���&�=�
���|�{�,@�رp�� �-���+v�7�_
�g�F��W�\Y��̶JI�Y�D�n�%in�e�ƜS�Zѹ��ف(�""g���b�5�+��p`��i�d��Ƞ3z��i[fL����ʋ�-���H2��\���H(����yZj���[~ArN��S����z�/�S2j\Y�X<'7:;O�kh�tP�X,�-�R����߿�z��aq���3�����a����U�[���G*$�P�oOk � %r	xN�I������z�����!���/�55ɟ���E�,�W =���;.FP��Z�y�5�~V�i�_ ��!
������c�x4nͶKRr�h:�"L�wJEUO���v�J���#��fPT�w��p4�=����֬�t/��s��CCC�[o�u�+����Z���"A���tI�B����g{EEş����|P[{N��K/���Ԧ�������7{�{�'3�v��  vQIDAT0�B

�!�b_G')dp��ΣG�6y*X,&d�����[�����E������i���|JV��THBA/x�!��\f(��y���jf���Q�ED� ��mٙ4cHgR���J��X'n��">잕o0g�=�P� G�p,Ҳrɲ/��گ�=� �c_�v�E���mr��VZZ*��l���N�Sh��D"GgΜ�̽�޷���6"�)B��h�g?���3��_o�k���<��N�)�p�����o˂��=��>���+/���������p䅿�7m��JFUe�W�����˺2�����8~���z������!�����
�L#D�#o����9Ԣ��:����F"%�v���ӀK��S$$�y�A���y���TW\��>��cǎ���c�F��
E���1eʤ?�}��֞Ɓ�ȿF>g��y�7����2i��2�����)+�bK.���]&'�P�p>t���C�M�_Y�n��������h?�s�d��j�^M�H(�P:Ð	Jr?��U�0f�w�!
��șqv�Y0��)H� �@:�(�̑&SYJ2�ET$,t*R��+(4	���S:~;���@8�%��{��ɧw�$ỸY�֑i���!N�T�yg��������ol��\�d��Ҹ����c��sȮT�z�Hn��CCg������>�"(�+�n����>X���u���pd&Eh���m?�,/5��<y:�HP�!I�L �>_����a�L�8�~�!
�������T(̦d22Ť�f�RP �P�E)�JǙ���hP���B�k�wU���z�h������� w�����__�U*�UVVb999B}yp�\#b
��/���?��q�1ǙA������B�ϧ���lY0Jh�a�d��6��IB�0u�wT.;ZMiS[���o�������W���:zU�BS��$Y�������OU_r��cg.m���Dt�3DWS�<�NXtY�(��ӱ$����g�4�Q*C�@ ��p��C ��`RD� �ζ�R�kٍ ߬���f.�����wgee��B�p����Cxh���u�]�ԃ>*�/�a�����\��G<�@c�68]P*�@��
�^��`������`����/���K�ҧ����{Y>�/P�ӊ�,#��1��b��i��������>���ً(�""gg�I �Z�i������@��V�cP�k�Ngh:ɥS4�I SK)ɠ (*������?X���k�PT��;��w߾��J^̉��8u� '�����]7�x���{�IQ�G�<�����D̀%sA(\��J%`�A���ft��֓'�>�ĳ���.�QB�1�De������ȺyZ����m����6=�A�Et�3Dww�$�0:X'���4 )�.4��i�wJ\$�N�� ��*R����^fÐ=��XGc���\���[H[�㣿���C��d2O4�L��nGZZZF���ry$�||���b~B��5`o~���E�4j���!p��`�CiQ!��+IBߩN(�����,�9�S��k/�3�d¦�bY2�"�th�"�Mӻ\~ݳ�.�X"g/�����!�^�D���)�A��h(p�vxAe�CޔT.�#��&͚�hj��M��(���	P$�#&GkS/��_5�H���k�U>��'��h'i�Z�����8����9p��;�z���n�|��S��5W�]������P��!��&=��N�!G�w'��!YF���)@3�AH%�`$ ����E:��׽Z���v1E��Gt�3�0�}�
\JR
���Aނ3��I0��{u6�K<�h������ի�]7\1{�NWH��V(B#�=N:�V�q:�򛥿�~���׏}������s�l6rҤI����dR蘖t���Kǋ��f>�ptuɺ�-t"&9��	�H��n� �LF�Y-0�����.g/����U#�},�78mELe �Js)���0�K6���?DA93`L<�C%I�4)h�
@�4�2.�dR�L���w/}�yZpɯ\�����w�^��'x���es����֦�#�B���={l��w��a����|iAq����\x��̩s�Y���w���(棏.�KM1VPPh�ʻP�*5��(���`�i�<�t�&���ZH�hpF� $r����͋/^�Q7y��Z����."rp8h8�"Bt�ɌtY�$($QX�,��7�z��5�]>kF�����:3���b@��8�W�77������>���5����k��{.+�ϗ��yH*�t�e�T*�RUU��O<�yVV�X4f�!�^{�iC��I:5�*(8��U� )F@_�����b�s $NG��=�nr�Co:�Ɍڄ�ۧ.]��k���T~8��."r IM'V�E%�����" r�6��|�=5?�?����*Ƿ�r�q�$UL&��	��iT#���ZZ�u��#����7յ���6�&a�\((����T��F��UU�_x�ɧ7�b>z��w)3, �X)	�� X�pCan6�z�hT���x�N��f�S]}�" ���sv�+u�_�&����]D���8ƻb%�b��0�I �J@�)%N�����7�r����1�~��r"��V-�]�f5!U�tv�;��[��KX���=wMZ�q���9?��@B����)��gb�x��j}��{�]W�eE1�Q	�?4��d2��CA��P^�P,U�f���^�f��Q�Uj���	�5����=��QN�b�5{�t�Q�ED� �D��iIb� EQ�fX�0	H&�o��m�������՚�3����;*�A�E�Z�t�����:Zsx���A��������7�)r\n�]��k���c�������>��3g��Ȩ&	�px:���3i
��1��@�ր����<�i� #��MJG!��Z��v�ER
Eh�̉��Q�ED� �M��L,dVH	�ˤ!�a� ���yc�[�g-���ӣ=����[��͞N��C ǀI%�M�T��۪KW�9ɿ����۷���c�*�H�)+ǖ������������ӿΛ7oDF=�u�rR��X,?L���P��8}�CP\Y R%d���U,E48���v:%2~s	�A!
������B<���,Ze^$����s�e��5ƥM A�X���F��[��-��`dZ�c�t:	Z���AcGcC-;���v���^}폖�}�Ɣ�U���"m�-0��p��Slf����+���W�:;�H�$�@������sl�1��#a������{��� M��A�*fσ�6�hk[���m�ڪ�����."�=���Q��u��P��(�F^GQT��eR���TT��v����7��	\����-9����h1�o
��7�pØ��\�����WX�F"p�@�Qe=Ζ��.|�;�h���5p:�.$��X�a� HHs,�C7��aބIл~�	��8�f۠���LB���h�����S��؛�FZĠ�����|�p�k��]?�f�d�|�8� ʛc�@���?_,�+���7�a�I�'7����V������J�D����?���|��u���ZQc�2��T�z{ �H�����q������_���'�A=��)��d8.��8��dǁfh��SV͟|	�w��a�h���7A�v����uv�I�F��6�xC�����z~�b������|�xN���kZ<���$˰����@8!2�4��O�hX�v�����xڽ`\X�m9�19�)�R)X$R�H����S{�~��[Ͼp��e:�Fa��C\�>�z������������J1��,BXy뭷|L2���J"8�.��gh����^C�h8�g�h��� �L�� �WWB���<��1���W����]D�{����L�fj�X�����i 5Z@���w�	�iK$���Fjj�Ғ���{�:�����Ro.Uv����ӽ��r��T�*�����t�tP#pIRI�7������2e�D�:L&S�$�a��Ҽ'�T�j5d��m8ssr!�B"��D�R�8$�$$2>0�ɤ�L{���b��Q�ED�'�`�Ǯ��\�®1��L
0�׈K�8�-�{���v�uφ���ٶkwG(��V'��EB@�V�bɼ8��*�#*�W�a�:;;�aӌA�{�'gU���^����e7��$$�Z�"ԋ�pņȕ�\6T��(!@B$@		ɦ��n6�������>���y��K�	r�����}޼�����dN��|����w��K/_��/~���o��Ǽy󤦦����`H������P����P�f3�K��SPUYN�ƣH�SI���`�[0�Ĺw��Y��l�Sl���<tA��9M�:�"�˝�ɂFc��,�CVE㩖��ƀ�H:��x�Ѩ�;U[KV]�h���� ,�{6������`�T)G6�|P�����.J0Ma���;��;ф@/�1C�x<�ٳ[����"(��� +d
`�@�i�r�D���}�CQ`fY`iȥ`����9[0<U500p�X���.�::�-��Ϸ~��-��NCZr8$r�V�	��P��G*E[�;V���=erk�T��:��AN���(�4���~-�$�B��pƒ,K{���m�Ӻ�l���v���s�?{�n�;ŢD
�yA��E���xLF3L���P���@�	��f �N_���M:v��� L}�w�����頣�	��,7a��'0L-� /����,� ̃ 8���,c?���lt�k�qRA������ͽ�G
,��D�yͭE��M
�
C]�`dhe$����_��e�]6:3��.�niny��o`	 n�9��$!�*�����`�P�P�9�Lv;��I�q��$XI4��K����cZ��(�肮�s�uM�.�᭼�x�(@1�-;�\&rO锖��"A�*#����Yp����k�f���X�C�n7% r��b��Y��n����v����|�%ū�������WZ��Ey��MBN(@��C�L<!I��$��hZ����ALe��U����av�����NUU���3]�utNcG��s%q��c���x:	%��Y�3�C�TЖ���e���Xmoo���X�mɒ\E����U���B�4������`q�l�ؾ����۟�z�9�9#�Vg�������7�fS��4�	
�_i�r^��cSS�������j�+(��#Q�;�`��h�����5+�ΌGt�iFmo�~���l��G��*O%�����h�U1
'�
l���cX"����>�-����]�q���O��w�e3�h͉%��8��)8>֧Z+=S7]��?_���^�9�hll�~��_�ַ��j6UK���<O@8���)�Ї�IX^Y�� �R�%2ʧS`��e�t:�P,5��@t��&��C#sj8��eL�e(�UV�Beuu�ol�����c�hE7�
i�9�<R�~�|�����RThF)(
$�yЖ^M&8�Vel"8��;�܍�pgZ�:�yӦ����o�1�Lf����Th�	���Y�@��ȝkI�4��n����=���3 ]�ut����K�6���|� ��HN����'�~�@�˴ԯڲ��(Ǳ�;�A-=�I[-�����(����ah��*����rR*M�61}����d2�Ϛ�0V�h2��t@ v��!��0	ApB���
 �N@4R��s8�X:���$��xtA�љF4���=wVq$�#T�µ#Fh��)������]�׳sg�v��N�������''�>|� ��������:��Ơ��B	ұLj�����&�|m;wλr��Џ&�q������]�����@,�����;x<��(faz�ܪ
(4`H���$Ԑ0<�)�bw�~:�O�f>����L'����[�f��x
+�x��Ĭg�Y{��4�X��k��>j�9<,Kb�\
�l��'�v��]���?������WD�b�`8DW�}`� ��xSI�wz���#L����������#7�!rP��B��q`�F�;R4L����aPE	8� F�"'�E�β�����:g����L'�4�I�j\4n&	�b��浈�������כۼy�<4l���c�R��U��8޿�m3�����}``�~}�����HX����dR)'83̭�g^_0�}����g�4�d�0��Ñ'@�HE��v�a���0@��C��� ���(��4�EI��l6k-��?�1���.�::�Hj$��IG���jg���,H��*��nm-'z�7oޤ���],�[,R�t�X��^���o`���߶�c������j���8"BjL<��H��ry��s8�B�{�"GH�}}f�Պ�2fCR�RP	J� �T��F����@&��` ,��&+(�r� h�����;��3��]Gg���b�a�XqMГBrbI�"�s�E���RX�hq��]�R6�����dV�Hdv|<����^�Σ�Uе���|䆚T.��7��8���z���
�Lp���
���׾o��>�ǹ��"��ऋ AV	�Y�A�!�@_o,�;��4ÑtF�q)R�@R����@�,�����M�t/�ΌFt�i$�4s@�i�1�"A!Ű��6Q�w���5��ms��!�}4Mc�>;t�l6��jk�F">��>���8{�ȡ���;M6'^*�`�$CD�
��t.�l
\6+�&&پ������6�z�ә�K
� 	J�%�ĜPA�1������&��ad` D2IEB����8E�t�-˲v�M��.�::�H"��iת����"CI�d�ב�z�\�J����q��ԍ~^ʞ8,LQn4mݝG!u N��7o�'��:�1� ��"0�B��B���qhjl;E>��Ѷ��%-7-=����m�ȒD�Ph2�E�;*!��ڄ�w.W���.8`ޢ��� �����AE���H-3!��ܚ�dt-8пD�i$�ti�H1�$P�d\4�q(9���=gΜԜ�9��{��1�LL&�Ǵ4�ȥ��������e�ڵ{��i�1l.���b�d���E1�*j���cI4_(����"������K3�CZ��)K���,LF� RrN�E�&d�QT���93yP8��&!4 o]�5͂��A�$EIV���	��1tf<����L���|���:IQ"Y��R�9���@m,��ڿKA�\��/~|�`Gǀ��G�qB3�V����b��x�y�qm����e�r56�J��DX��j�+�V���Bg���\�G�4��������T�r�hw-�~���,�09u �4~�ȕ 9 ���#�`t��_Q��c�'!O���E�NkɌ�l6��ΌGt��b���3E��fI��Q�\���A��}� �Ciԕ+���܋��}��>:��DuwO��@`�믿NǓ�������B�P �b 4�����C-���~�S��օ�D
��|�[0{4�tp���z�������c,��%Y�hX�A���~N�
Fc�hl� ��>|�^}D�"�q� �a���.��EQ����@t�i"�JbQ0�8��,E��c9D!iuے�(�˗/�775� `��8� f����^X����E~%i2� 01�]#�������}��y)WӬ�X�	��$��j�J��668�<�c�3�.�tf�(R4����@��"X)�Ȱ�dl�p(��8��[C�QC���W�w���dS�3 ]�ut�	jb�(f2V��q�a� �IE�K1����ʙj��y䗻��_s�<��H�����f'�ј��矿�a�,��>��@�$�xL�$���z-h^0s�[�]����qs�a*�@�[�m4�����;��.�g4-ͦ�O�	�4Ә�t,�B	\ډ��X�D�@?��p)���B4Gb�c@�!���uA?�]Gg�Hf2�"�����Ҧ�������i��!�잫�>'����M ηX,�T*H��(�LǏ�\�t9%�ލf��&	�B��TmC�N���y-b>�n�ѽϮ?V _,��]N;؍F�iཽ{����c�ҥ"��l�,Ql�����HF!1��f!�π���LP )�SQ�F���A>��`p\.��~�%�`�Y�#}�At�i"��a$�S,E〜RQ�$k;�X�@�����/���׵�����n7&��r6��$In�y�����@b���ѫrx�c�1�^w]����Cc#�����X,b6���9lG��W��z����3�Q���FGw���iF��tm���R/��醣C#P����`b2 �u���dpp���𝲪:3]�ut�	� �y@æ(� ʒ������H�T�]{�zv�����\��9U*��R���f˕�4we4!
A�X@-+���5W�1��]_;�fw�@=ϟ�����s��h0`���7h��uA��h���O3$Q����C!����H�h�`���� �	r��D�X,- N�S�V+��|tA�љ&TQ$%EaeI�5�ȝ�$N�h:�2�%+����ܹ�9ٓ�dYĵ6�@�%K��]s[�X�v[����-?oE��u�L*�8�Np��X���4�ۻPݾ�(�f�:3��5k_*Y:ߌ��l�  ����c`
*93�ASi�6жqL�*|^��К�}z�3 ]�ut�	/��в"a���@�J� ��)���VX�r��-�7�`��m�\�d2�t:!��]:��9w4K�{��a����f��zN��ܼ=���x>ﵣA�±�M�F�/��lF��@gF�?�`�W��b�n��9���O����f�d�J�HR�(� ���^��hю=�Z�;� �Aqg ����L��G��!0��Ρ#C,)@�R�)�v�m��M��{n�l44s�r��9C�0���B!�Q�TcӬ���ֿ[����6��;v�+�%뫭�7�؁��ܮ��#�і�AgƢ������c]{"F�o�0r,�MV��sP�΢S$xD�1`��Yb�(~<�v��3::�o��肮�3M���+��A�#�������x������_��;�w/�2�x��!N��n�X�{�ڑ# \L�S�Yͳ��L�/����������l��A���B4�W9���]xU۫Z�u�N�g����y����E��;���$$����PRD d�H�#1$�f�v�P�����,˿�⋵���kG'AgƢ���4���`(�;���&�>���?=rx������Q��y�y��CCC��x��]��:�Iˢb+W~s��;��&c1��j���l��_����Ft�~Й�4V�IY��h(�4��ɨ��lV0���#�j<��&��B$���r�"��1����ݻ����m�T��.�::�D�X�]^~hb�[�0Sd4��?U�󮾰o�k�H�4��8^�c�\�����8���������r��L��]r�O{��������O�x���x��j����:3��V�eŪ=��9X�=�b	��WA"U *��T M�\T��D�&�I�af�?ii�<x����Ft�i�D��[�˛����,�*��SA�S9's�%��zꩧ�����:;;���Xn+�/�&�JC]ݰ��>��Z�tu셺�������D���1�ՊErY�P(�j�С�A���h����ׇ����X�Tl���L}mp�������"��fD�	��+A���$����]�vՀ^�gF����4Aд���JF��h�� ��8��Z�������>����R�m6�i-��n��W�p��K����KK�,9�C����?�������v?�Z�	���
�72����/�B������ƴhQ��P�1��u�� �l>[>gγ�e�զ3���"q�0,�LL&H�T9<<\�.9:3]�ut�	�X�����p$I I�8rF��{,WY[[�]�b�[;v�<�����X���Tܐ�q���R�W_{N�����%�:�˗ո�V������G/�nٲ]��Kmmi��%����҂��"�8VWYڹt����)		����-�3�Z�
�H̵>e��b��۷�k��3]�ut�	�!%�p�xۡk��	���8#^(�'Aw�\��Ͽ�c���0���Ea�`P��V��8�y�@�	ti�Tm`uk�O��ѭ��q^4�m��`���a��G"+��jkA.=�N�X����ݍ>�pR!�|	xp*��WUT@(��`C&6��C*#N h���RQ�?��Uk__�5���.�::�G�WeQU-�&C�Zp���ϖ"�Iеs����I�r����9l�g��B���~��?�A��4�V8U;+?x���m�'3�Ns��W{�]�j�P}t�k.�w�tYtf,]�{��յ�02Vv��|�p3Y\&38yDP�E��qU~۝k���h[@�N�G�}�����4a�y4J�,˪��IR(���8a,���G���v-�v)U[9[���Ι���r�����p��o�k�N�F��e!ל9�rG�/DbNoԁU�\X$R��ө�o�e4��]��D��c�L��ł~�p
�#0�u�-F�9��ڡ�`��@D�B>�.����E];����z���.�::ӄ�a�"K����3Z~
�L�P�y���i6�/2,[ ��\s��FH����x�鿜��e�T.]�;��[���~�����bk���2�d�������W����~�]��d�����;'Y�1@.<�BF[(��l����I
b�����y�X �cAVd-���ypp�u��g ����L�ɤR]^�,W��p`�)�THNd���8O�H�ir�\�(�&��|h��|����[>����:�|�T�,Z�p��
�˙tfv2���Db�s� V�::��������:t�>���іo�Fb��d��D�"�y�B*v�<&3Lf3�� O��@�-�k�>�v�#�$I.�L�;::�� ]�g ����Lv��i�I(���e���YWD���g�Wm)��F�J9�T*iId�X,0�Zլ����L��.�ˆ�/E����t�K��[�o��8��R���8�b�p�x��fk���,���>�]��b`�>��eV���L&R���\A(a*8	T8�0�8�%xA�a ���D��Qt9��;��(N�e�{JC�)tA�љ.�f�h6F�\ZQ%4��qF��I�= ��)0N�Ӝ��|�H|������yވ�U����箼ꆲK;U[�]���g��1�,��{j*���6�.�5��d�3��D�>ݥ�;�,�@`y��a����΁�r���H��'ʓ?����
ѷ�i*��<(�0��)��1�1�0���PtA�љ.jkE��.����ME`6���p�#��$�RIۂWm���ܮ	��l�H4��U��JM�B+�|���x/��-�����G�y����$#����r�-�Z���2vly�#���;Z��Aۖ��8�����&��Pc
�ʇ$�,�&#8x#��;�[�Л� MP���$Qt�$q�3O����:��肮�3Mh�E�?vC<-	bQA�E Q#MS���b��$���K���XF��m1p9]v�&�&��u��W}�~�ť_w���7����Z�|�Nk���	���ȱ�����sh�?���i�={�o�~�z����rx)�Ĝ ��&~9Y Vf��e�d6���C6�;� Q����׋��W�^�ф\EF���.�::ӈ�ޗL�r�|֩Y�rP�@��6-���?k�X�H�JkgеL_������f5A*�I��d��
�e?��ϯA���]�"�����/��ՏW89�1>4��.��b���\M^|����Ot�8��ˢ����7+ ������6l"0
�l(-�k!&�	ȥ˥�h�HH%����˒�P��k.]�r���	3���љF8�3[�ɔ�Jf�x��,��b2l��P�9��,I��s�ڲ��i��t�>��j�(w��\��/lB���ͳ�|&�z��/z{���͎ĢDuuTڬ�H)�l�=��ҽ���Jw7ձu��^�o�r�i����@�I_(���I�C�P �$�FޛE����
%�" �(j�9Z�����3c�]Gg���H`>Q��Œ<ˁ��05��%�����?kǉ��*I�����-�grYp��eA�����$300��G�����C~���+ �L:��?�������#	Wo �q�|P�X�M�Ǻz?���ߏD}@���d�]�����+�~��y.��D&2MA*��;W��Y����4�� g�\��e��E�*�2^�S�lIr{\QI�Կ��.�::ӈ��*��d(W�D*	�~30	�$X�c�����I�"ʥ|>�j�&�����?C�	q`$ �`M�8q��7lxi���ڝ���%[^~a�H{����uh|��3{4�<�$��>���W_�{Џ��ˡ�������<7M��5��C�� ���Ψ2т )Q9t9������U�\&�8P8Q>A�C�ؚ�P]���Ϡ�TtA�љFL~>ϘM�h\Hg�$A��q�6���/m(
�F\UTE��h.=<T�ż811Q���fy���X�VЅ��������UUU����9ouݺί�o�ϰ��H�m�ǚ�^,�9���O=��4�o�����x�ϕ8~������RU��� ��A9��H�$%
�
,�l-����a$8�𨝤� A�E]�PY���&�jk3]�ut��0-9|!a*�TYC�b��γ���Q���Ni	_ޭ	�RD�Ų ���e��q\�T����[�h�5H�&p�J&���}��z̓�CW=�УZ���S-�c�_/<��ܴ~c��899i�M0��Cb0{�޶�y��vx�t:�͝��ڟ,w`��z��s��NA�T����n>/�3)�όP h(��t�|<����kY	4Y��x�&�2(j���>�o��\tA�љN�,�+�k�{;f����f2`�9pLt`*T�d����*��E�b1���˸ H�n��3$�l�}�>?E�T�8F�������;o�P3S�j���-�w����9k%f-Z ����SW����K������s��ӷ��'��u��������R	�&' �� �vA9����JJ*�%	�,]�d���I@�=g`�r�5����N��ng_KK��`����4�-U������$M��6�J�N�9t��B�Ʃ�cFtY���0�"AR�P�Ш��a�w&��+�PH��'?�����|k��L�b1����j2�ϗ�w��"g�ԩ"�1�zypݺ���}��+���g,�Uy�X�$��=�?���FQ��Q��/��0��/}n�]�ϭ0�<����JE�I�do�����3a�W�`��aH
 �H��r�4��k� �K��G�E,���;.\���.�::�L��ɗf8����B��JVR�JZ�����	e�ݖ9�f��q���j.��0�Md,���7�tS�>��'���?��Ͷ��L� �Y���n������7}��?nC�3x��i���Ժ[o�K��ךZ�K���س/���H��-o�x�3m��ۃ������?:��Km���ڥw���p4����$�DA)�����c;v\�nh`)�����%H�(D��Imm/� .�N��/�2|&��8�Ot��V�?��肮�3�X]�����hlr�YbdP�l2��0O��@GG'�˲;r�����$�Z�6��S�	�Z�И]�wl߾��l2�5�$��ts8�v�8Y��<���O�wފ_�梧z�뮿���{��3l�Z��:��C̪�C���0uyۺg?��U�]::��k���|��:�|��1�~���� �/�1"�}�c��a盕�Ɉ[}^�`yEcp��� �
t	,ȕ����k�k���G�(��ū��tf2����L3�ܹ?y����`.�����X�,gkIz	�EБx�E��R^�e��y��e��X�2x|�hW__���Ͻ���߽��q^�ĹX,N�sح��ё�����Enl�)���YS<��c۞��{�]T[����)��dČ&��[,cGWlx��ux�-'<�6��F<���Αák\v���W�%��D!�*2UQ�3�чvwu�6VT�5MxxlBKJ�\�2�y�h���(��h ^� [�g�>眷�Z��.�::����ف���
�]�d��q`3�9|<���СjtIש�u�\��ĕ2鄜��@D0�&�&I��������#h�:��+�?�m�j��97V�MK8�g2����Go���{�O�<?����|&����D׫[����kz���������ͳ+�<>����a$��~�X�����/}n�˻���#�D0ǆ!��#���.���?���<�͝��D�]^h۹��bI ��
��\>���ZX$R)���X ��Ə|p�&z:3]�utN��y�b����8�N����cV��?���zxA��|��劏��)ڀ��.��������*�@��`�booG;�M��>������V�b�܇}�usf� 5;p���ዟﻯ��ɞXl�,��5IP-��J&�*����ƛ���'&��iF;������9U4�̂c���
l`d�
@��/XZ[^x�x[��[,^������$��G���@gXP%mH�g!^,�l�7� O��|��'/�r�$��xtA��9�朕48}�h4M&�U��f�X�pw�Yj`�V�je��+�c�T*
�b�b	6;��"�H����5ew���}������{�SGy]�X4��`---� K�D:�������+����K/�4t2Aֶ&7m���{���!��0�q�Z[f�ܪj>Rȭٺ�IwM�w���>}��_|�׾8+�3��~Os�͍�1��I�d6#�i����?�ܯ�~�F,��k0R��u�B���l�$ �N�E�x98�1�jI��n�g㭷����-g����jk��K���߲%.ɪ9�\��aK:KK�X���GL�S	�\]QҪVk���<�ɢf�S�hձcA�o/�馛B{�ݰi�j���Al"8��aյU棝�W����u/YR��<s�7�_}u~�C�ش�g�h�V4|*�J��&B�k�����``�3���w����K����]�=Vq����/t8���]�pAGg$K
D
���+.�K�(1[������jl���H��@h\�3g��0
I��wx�Bټ�Lgz?����[�r�^U�At�Ӏv�k���ۿq�XN�*B�USU��0�"�t�hEn,v�s��s?��Q����R�!�2N OL)����1+���j�?~|�������X�V_<�N��\O���T�kk���_�~��3�*�z��Ltz�gg{��c��d� 2��.,]������=���������@���q�n��FI|��l�DBS �R)���^9���t�_���L.%��l�8�B�#��p�[,@
%P@E�:E�| ����~�ꀞ[��At��D�E�R�#��lnQ�P��b|#>�N�F\mm{�.���1�ތ�Ȋ��8�3�s���!����Syb���ssss�{���+7�|�2��vm.��ì�&�h����{v��Ϲ���ѽm'��&!jW��O���D�d�6�n_<�H�*���
Q
�}��o���GzUu�V[��a�_B��g���א�����UQ����D9sQI��ص����'_߲�@����/5���c������;���S,`� �A�� �3E�������װS��י�肮�s���ȟ��Mۂol��H1-�\�8�x�d$���7=p�3޳*g�m6[O._jF�H��]>���8���ۊ.ك���ck׮��_������ʑ����_{LDC��]x��~�6��{H��O�:0w�z������A,��#�2�$MF�6
pf��[���Kd�T�������o�����W��-��a�F>p��,Y����[���_�p�����44�6����T8>\;I�]��\A� �V��|l��+wA�8�Q肮�sY�|ٱ'_}�;-�-�T
������S����η��ю��,Ȭ���XQ]�w��Qe*��"e7���4��o����r���cG���'�FF���ojihhh���'''��п~  ��{�����8��{��,��K��}�/=��_��v���D�r|�9@�\VV��x��/��GAm�՗p����7?��#��n��o-�aY����Y���B���g�c��%KS���?xm�XhيVuM� 4>�� 1Y��C�V�/����@`�H�C�,�׿�3]�utN#usO�*��c�ĥ�b��*��T��r�}G��߲�-8I�q�X��_��ȁ�CŜ p�R�,6+3��[���킓�i�i";�?r�K/���:���>44n�����Y�һ��F�2PZ�񓴡M0����;������چO�J���HV3���ZM�T����>K[���;��!jW=��_�6=��-U����h0ͫ�c�xF&�pO�!La��i�߻{WKeC�����%�p�� (�,p�<�Ƭ4,E��(8"�C�$E[ue��S�3]�utN'g�]��z�����Gܬd�'b���7�C����x��D����җ.X<���?�sł-�L@U�hN;��׶��i�>t���Χ#����,���x��d����T�`6��!9��u�7b�ׯ��5�\s��l���DS�Y�ٳ�]u���X�a�u�,�e>9y�?�u���?���&�v����͌<�d4e2��H8�sDIHb�tZE9�� �=(b<N$�Ǎ?��?�r�����EU>���&��Bpr�1��&&�q��7:���1z��%��d����!�J�A� O��nB�.��x
M �?�^�ld��%�`	�A�g ����F4���������%��)�*��"0n����ͷξrd���忝�?����j,�M�t���*�[���l�8���ʁS�hkkk|t��c�|��P8�	���ɥ3��%�3r����
a�[����u�����#'��ڒz����C��ꪫ����$���*��ǋ^{�w���xbbr�-�j������D�x<n��;\щ�-�:���5�-�I4�%^VeJ$J�J\VEE��cD���T%�-[:�����7�R->�pY,@0�p2y�B!�Q_LƉ�:��M���f���	�"чLj�,�"��8�|d�AS.�����s�[�`���r����i���g��>�-�ݽ
	zu>�#���.e*r~��on�����ج�Y=G�3y^���x����C+v�ر	ޥkM��Ķm���7�T�S��f0p���q���Jk��-�JS?}Ƿ�?��c�|��C�(�eQoo���}?������Օu��dU����Y(�K��e����R�$~�g���p�xww7���g:��k�9��X�remxjj>rޕ*A�U�� ��q-�>������p�X	��(�y�b,C�V�V�H\8k�Yꇗ/3��
V�B�σ�����q�)H�)��a���Æ7w��0V.]%$�}�G�,A-�C}���6Y;C����h��Z���Ƴ��i�Г��肮�s����?����c�G��T���lu�����iq�+�/P�o����10��U�m�{��Ёϊ�"���1�ǉ$����]]]ڲ��ֳ�����ַ{���dS鏘�f���f�P��@X�VO����u�Wj��4G�����ҥ���������{��nYy|`�U�"̯�í���gd���-���8��������N������H�������P�MZ�Y��� �$I�;�J2�`�;K� ���E=EH���H " �E�H�ePsY(�K0�3�W͟�!1W�h
���`>�9I$�Y��b�W�S_o9Z>K�<�*�x��� �b`�q �i�e(���q4�H��I4�`��;��L����j��T�3]�ut�οi��W6�]e6m|I 3���\�242����6w!!�['���c����g����1�r�6�E� G��=�/���*tO����Ĳ��?���nY��A��3�620 U�5���9���������L�����ZᎿ���B��ͻ���?�34��En�ꑱ O�"T�T��˦F×n��j1�����SV�{?A�Mcj߾}�-[�4�r�-s��+�0}fE3&��ɉ�LI��)P��
%���3I QUʵ�1Y�6>����0�s`tY!�J � q�%��QX쯆�/[�E��;H�<享=��p,g��͢n�<�I0�+�d<��?f�4��}m01�^�����f�PA����d"�QB�����PZ|���7.�3]�ut��3��?����~��A����vz0+A�$�������?�"�`F�o�;���b5���65�D2�$K��V��w;~|aGG�����O'D}��������5�-E��|:#c0w�\��v�_���?�&&C����+�}��N�W���oo��Wn�mo"�h6[�F�h�A�Ξ��72+�K�=�����@��_-����0����6n|������|~9A�ȁ)�@K��k5�eY�g���P� !�$���H�e4��<��a�}k+�*hhŐ?��}GA&3C�N�ʩ�V��ų�`�����Rв����@��xh
��Fe��VW��(>�Nci4Ih�7fϙ��	�+C�����$��Po��E�����dZ-�TF�Z�\��O������.�::�K.�b��駟��o3d�3cԎa^���&�׵��T�C���tf�.Z������b�&��c~���\_o��W_}�]v����	Qz�����#7�L&g.û���&��y�a�ڴ���O�l~�W��]�k�d{�m���?$��_�m1��� ���J�SI�@8v�+�y�&$3!Qײ���	MП�{���v����;���|>We�ٜ���d2�(��S��`H���C.\Q%���IRQeI�Y!qy|L�TU�$����+�$J%Q.��B U�)�O��l�0�6X|W��Y�g�x	Z�͆�Y-0��G���\�TQHf�~�u�Kۋ/]���TT¼���&o�~8Lu+!�&MVؑ�{L<�cH�ד,]�(��՟����A�Ft��	l�����|뵽z���f��L� V#F��z�e���߸��/����Ӯ"!j{n���t��S(PH@�b���Vmܸ~NWW�1��im�5�C?��O~����/!܄�#�N�}���SQ���j�q�j�9���O��g�w�yǟNl�u��j��������VH��W�a��� ��%�So�F�J�K�?��F3IV��~km}_D}vfÆ�W^y�e���Kk��mV�Ĩ�x�y(���PȂK��2��$.��(���(���7��R9��=�d�$�5$�S�l2��n�Kf,�0���.�s`5;�U��h^�4��y#8�ȝ{�a�x@��^ձ�Ə��׿�-��p�%��?��_xpR��N4�`�Eh���E���L�c�U�mV!ϑ틯��s/���N�9��]G�}d�G/�ط}��x$YOK��K�SfRE�S?��T�����R�U�&.\�����g��qs��ļ^/��|�x�x]z/��m�����ů%���~��dl��2���(d�%p�<����~������o�|���������;n��7g�7o~�߻��d�_�1�B1�2�Ǳ��&lYs#�ON.>����
���%�m[k��������ڿ�m��v��-[>�޷�`6�r a�TTY�GB.@F���\AȉGr�t�,��3h�[��.w���~���*T57
.�E4��k�A��S~��W66>�u�[M�8���-��a�o F!�m�78�4^zq|���n��w��V{s}S#v�ŗ ���^}e3�XJ+m�Sp W^c5�A� /�yr���&q��W\�Ѕ��mVW�/��@t����U�U�_����w�2�xI&-x6GU�݁��v��=H�����^YYY\�r����}_H���D"A��ց��d''��]�v1����Ib���KS�����ɽ���$Y�K562,r~4͢9E�����ys��;���Us�|��8���,�ڞ��M{������y���h�,���e6̫�")��������|M��߫j{?�-��`94ѱ��w�[��|:���|�\.G%�I�F�% T��QM���NUE)��D�8̶�-�{�^tv��fe��WKK�,��'Ǿ���·���7��T��Z*}�ܪJ4��x���M�M�`A������9o���YЊ�^�8���6mU*�� ���i|L�"4ج�@3HH%�DS�kho=o�~������tA��yy{/��رo>?x��!*>2[z��u!k�b������g�j��]>p�u�K�z�{��-�L�&$�F����&�������>��t����4/]���u�=�%Q��11��مy<>00,f2�e+�7����o޵p�Ν�۷���˗Ǵ6�:����{�}�{��\��x�M[���`��0���p:�5G�o��7�nX����#Ǐ��ln��o��֖��gk��W�z͋/��	��^SQQ�����޸�`�\*U�i��0�HF���b�8��_�r�/�N���q�\
D"*��A��֩p�u��U��NN��ttpO|��Vl�q�l���:����P�s<G��l^ ����<`�>���;(9�;_�+WW�4��4Qa�PB�Ȁ k�^aK lc�1���}^X��{�lc�m�1z&� �@	%@HBa43�h�&OO�T�]�ޭF>����ƻb��9���P]Up���[��/Lm �s�O��{{<-H�ˁ�I�Ӧ��B�3�`�j�6�WN���� E��TDopgc��ʢ����o>D̚uV�,��}�B�`��!�YJf�+�~��yaF��2d�uQ*��S�������;1b��J���W,ϝ����/m�ty�N��^?����tΖH$V<��3��������Y]]]I}G�������X������|���갺����wU���m۶-�gϞe߿��ׯ]�=gΜ�u}�ܵ��ɇx<���I\Y(���}T3J����Ej�㢽/>��<�z��[� ?�.xK��B��裏.��/�mY����	:ic����8)�xV2G�(2�������?s��uRI�MY&Y�)�,%�]bh���sO���@���������
i��K�߮��G��G�Wΰ��έkp��U��\uuCF*�F9�d��0,����#��F7�̈́E���(����w��U��}�X�P�F�@�@c(�L�R����v�/~{݆�- �������O,t�,�s�U#Kyt�O�ls�g��l{!�̐6[�.�n~���㩭[��/�<o%��6o��ƶ��zQ�$�)6����Ձ�{���߾k{�t�Gݗ���޹s�������u��L��T~`�d�,E�`Su�eS���~��G/~q㦗o�四{S����5o]&x���~��Ρ�0m���i�Ύ����B[�T"�t�YJ��y����;o�x��O���,�q�����J�-<p�M���_mF=�:gu��Z��8�u��<K�������I�)�x:Iۊ���o`(�`9�Fwe��ZWI�d����`�J�*�蚮�A3�Kh�0��X`�</4���)��<��P�K`"!+���F���]0P����Aմ&�h�%004��*h�x�tn+�����P��S��r�"Gdv4����u_�V���|0�A��1�� +������;�>����X�
����2]/S����ǇF����X�BZ��/L\z٪�_~m�D&�Ē	����*d���y��/w'���^���E]>�t���Gy�{ӫ�^W*�.p
vO<6A�&�0����4�3�M�{���]����w_������C������k����w��J��F���� IdGW'�w;`is]�q�O������������_Y��>	���LyVfl�/8:0�۱��O���נsq���u$bqJG�dY8�ֹ�a�@�$xXЉ7J�~��*�/zl��~+oCi��榬/����g�f umìt��X�i�S�\>�I�H�B���CN;�
�--`��9z� Dq��.�;h.7�7<�F �ڟ�]�y��6���G������n Q���u�i��6�%� ܁�pxەW]}d�7gO�
��?�`�c0g	���⛯>��X��gt�&�ӞE�|`Dn�?�tG��~jtى�"���K￰c�Q	��:z�i_�
�E���@Owߚ�l؃����^=#����e�����~�tOߗ}����l��1"�L@���[[�-WxNX�mf�}�=W=��ow�z�7��v�ꞅ.z�Ww�3ᠴ��T���cm�r�R�%T&<5.HM�uF��~�C��m���yW��b�z���"�� ?�?4��	Y1�{wÆGO�*�Բ����㫛g�s9oss31� ��U�f�_�	l	A�H%�d���<.�V3��t�!)�H�$:|k��Q���@�GgP�d�#��!�JA� �@ �~/J�21� �&����������c18��2:�D��9]�����p� i�ZV��� �っG�B��A���@Z9I�Pt �Bdʠ�x<�����}m�w��[�HW�[���8X��Y�������b�z���n����5�T.��F���9���}?�ݿ����ƍ[�/9b�%m{y�볼�����>�#(-��X*=��O��[���Jk.{��ݧJ�iO;�_<��#���W�O
�}�`Y+3c�D*�0XCm����b�ꎶY���y�ÿ���ǋ/~��oݴ���[E����2E�-��1�L|��P_� s��Y���cC�����=�_�����K��f�9prPIgm'�O�����������cc���/�L�eǛ{��ŒHz��y�k렐΂,)�#i��.tMp�t�Xpy�4p�&��hUYG�iUo5M�0L��L
='�E�6���X,��n��n�5|r�,�J	�~?4Oo�֚]5���1H's ���)��qE���N�I��Z@����ASs+t�8	�G� ��Ǡo׊E�+8��Ǌ��E�m}�����͞�wќ�#�5kʕ1���`,��1���3�^:W��n{�q�P�YYf�(YzH�(���phQ��p�� &���5�o��C�4E�>x�a",)�����{r��h�?�[H9��sh;o�w������׫�?|�j�����6�@)�*�G�P����fr�5����r�tϔ{���9���y���5��Ҫ�\�sҥx��I��#0�P$B���ӵ5!o�\\,�0{lۛ���|_,�rk�9��(>�����-X��|���|w?Hh�[�e	��4h%	<<�n� �\NU/ϫ�MI��bV��J2�뺪J�Uδq���J�h�N����׸h�	��oM#�D�V���hjj����C�pzh�iln�H�����1����/BC-�9wh$��;ЮH�vz@-Ɋ��&x���i�9mm�-�f��ϜY^�`��YZg���B�`�2,񚝝�d��w���x��b��R��b��W�L��[FF���K?�k��}u�U�gdG�ʅ<��f�L���e������}�8�@�g����ݰq�{y걯���ˋJi����*Q###D�T�a���L4�6�с>�h��+^����Z���n�,�&���48I�<>�L���*�OĨR����3s�Rg�;�DZSI��K��"��ܰ��7�}d	��S� �2�+�*�D�:���ɓ,�L��%�idY�&J��,	��瀫�f���f�-'8����6݂���b�1N�x^h�X����ЭuQEŪ�g���U!���G	�#�;��|�(�S>/�'�u���8���3k�,pE��tz�{�4�Y^O \��袅������K���^���9!f�R���=��R�>��������D����H��Ir��j�qW���B������xsh�r͗���:�MR����o���yތ8�t�'�g�Ý�չ�?=����7mY�O�/��|��h�\t��SF:+6��(3���./���C#��r��Q��:sfͬ��Ҵ�Kp����Kg��R���^p���G�0^�����k�SV�WWmm�!�-��xHښ�f4�*&e�B᪭m-�C~O���)�3���2W�U���fe�݁����c�����ӭ�x|�K��ڮ���*\5�0�B(��{c0::
�Q�P��Qc�A��Co&��y�����j��X.��tC��'J�:�r�<����_���V��n�a0,t�,��DJ����\^$O��y[]�zyFR9[Q�j�H���%Q��E1A���3�$�X_?��<��/j����_����1�+f�� ?��K�<��K�?�c����R�<ʹ�#��po/���|cUsQ�4��m%�%�\v���M��C�e��rBC$$ŀNP�s6+!�� �8p���i�f@��i���!�F�%k`��Aj(<Vʾ�5��m�
��+��O���d�ʺ �z0��9��晈��x���%+�c��L�ή����
�?
�S�!�(Qk Kp��QH%3���:M��ɴ�P*' ����]�2`k��tyaBW`|p�^}t�t��/�eq���wW���篹yݱ�V�q"�|��1����Q2GF��B�_�7�`��p�-�����3(�
�N�rY� .Ӏ �a
� G3`��.��d�۾��/������m�$�1=#k��c�^|k�w���>��q��������T"����p�����&x�A�z�(�:��U�UTU��X��n���8�I��̡��0������8s&T�7���0L����N��V:�d�i�u�{�i�C\��΄8K�"��������MB�(��]p�9���f�UA�o�*�\��ô�s�>�Cc�P@�t��P��L@�� �y�K�?������j��HFFG�����9�8�T�1��w,]�t�ڵ��Y�&��U�39�B�`�r,��4�/��o��}��F6���M���ʴ(�qH+$���i�-@�"�k"u�M�ji�G�b���w>��ú����P�89S�Ś�MA4J���iEIs��	�ľ#�u�b�sU��MU=T��(1�h��^��"nkU3	���E.C^,@,��\!_Y&�$�@��H�v���#��J�ᶙ0w���K�y�J�5�T�:��.��y�'!��k�5''F9���`�SVM�}���!��/^�����FK��ԡ�ˁ��C&�L
��24t
L��,��W��E�A1'G�a}������@��ޏ����1�~�7�L���,���ϝ��k���[�.�9� ��pf����P�g���7��:;ֶ�Ff9t����.����4J�N$�J��|��(�CA�I�h�D��sg���;���oڒsۥ};��*��T�gup�t�=$��h	�H����B�O%D>�N����'�D*�R9�4:��l"���:i��=Ba�\,�8�,��n�!�Z����@&��l6��	�ZeHr�G����G�,&h.'�����Aщ2~u5̚5����+B	�� �����3��_*A��@ x���A��@�OT6A�t�0�J�t���jXA-�!��D5
�"н�h�Z�])�hby �N`�w�Q#*��6�b��(����νj��� �Ӧu=�e��J�%y��n��k���5}�V��̯���k��$�B�`>%���4fvv>v���oپ���^jj��NE�)���%v|�j��Ƴ��xȜ�d�)�Ʋv�ꙷ�����#�"i���<��%��$�0tS5�ilY,:4U���%L���ۣx�$y�$�*���:���H�=�p�p�L��r*�aAZ�V�e�|�%�����D (J(��H�"r٪���BFR�'�q��e�X���/9�FGb�s��RI���U�6PIP�����
��XD%j����e<σ�΢du}[�eL]U��MU�I6���P:�uV�:`�V�s�@�Xȡ@%�Q�A�j��3o	�3���d��c�ft�����%m{W��b�̙3�.T{�i�`>i��1�O���Y=w�={_x������~�imhnv3�<Q��	US@V5`i�n�U(�(!˲�ʧ�y�Y���P��)��ɪI��iu�[�Qz%H�F�N;�7G�x���F�豵�(r<U�>G �]U!�J�$*BL#�j�	e�/"�sYGm�XLI�����BN3��U�l���rz�	�(��IM5,��J��@i���8D� �$p�](y`g(0Y ��H�4j�V�u����j�ǖ��::���k6�r�n%p�T���9T�B� "�6;�)��&$F�1�R��Q4H��nJ�i�o�T�((�x�{J��H$T�qѪU=�-�.X�@���1o��1�O!g�0h��>5zt��w6n����W�B[˔z�Q.�$�t
�V��r
�<�O�Z
4���)�!+��	$)ֺ�L1`$0(�S��6 �b+�<�X׵�<�E$�|I��JTEQ*����V4�@NeL�0�2�)$�fuS�ɥ�ɲQ������Uk��_6u�O۷�x��gv��Rֶ�Y��]�ª�
Vu6k��L:Wi(���̓T.@�h@�:�� n� ^V�A%��"��nU�C�G"Aڶ�������Z	]�Z��@E����M�X2i�ʒ�74M�i]���3咪�%�`t��v�V�S���>�����74��׋۶�:�)�hm�QZ����~ӿ��[����h�ɓ+E[Tm|�@�UbX���b�Xڀm4�����,IV�E�H��Q:�U���������,�Z����2�Q���Is,((իH�I!�1fFҐ�R�\��7Xn�r:{��jO/��26}��Xc󌔣ѯ�&Ҟ6�:��x��zZ�+�,��sP@���p�x'R�i�\N���%�]�S�13>2FU{�PL���S�O�Ai���L+m��(J"��<)��e%�?i�aʚ��e]Td]�tM!(U2M��\P!O�Dl�j�D��}���������3���dKK���РYE���,t�S�_L���~��?mZ0���&E������E�,�;8)f?���I(�"��(�Z�� �s%`	��&*R��ȭ�$n��L��M$uC�U�BW�e�hz�4�(�FAH���Ԍ��N9]��<����v���8�]�Ю>	�D�sÆ���Gn�K^\
��.\D]t�e(I�`������UI�^A0�Hf��w[[��M%�bjk(� �%S�� lw"Fj�a�p���*�)U��F&׀`����ut�(��As�3<�P6^!Y^������ٚ�ڼ�:X�z��UU:�ب�B���c����m`�c0��3�H�;��owfp���C��:�/8|��*�	3CU��N�,����Յγ��h�����%��d� 	�bE6�b� ��E�"�4�&I�� �}���N�X$�O,nmI7�̈3�ZYV���?O�2o����>|8����+W~�Ҿ��/��y��Mk�A566�x4
ｿ�FG�n��!�W����TG"/�~Ǐ6-^|~KKΰ�;|�I|x���a �w��V����	g:]yMABϋ"!��D�Q4)*b�4m���l���O��7�A�rUƂ�3��h��OX��$��5v�6l�̑��'v����}�}{$��B���J���c5aȗ�`��mw9Ql� �NC�2��Y�����iS��q}#��>��q�/���lrp�<ZZ���<jK�'N�p>���U���iٞ�{����%EյNm���H��]i@��y3���A����k�ht|�e�_��[��O{.\��W�B�`>�)Ns��j�C���O��8������\.�XK��Q�fM���Y���ӕ�:�i��=3.X��2�&!��E�k��-yR�"O��<��;�\��k��}���ѱ�sLjB���m�4�*TE��CCC���Q��S�5�p8�b��Q?�~�m߽e���K�	b�ߴ�3��B�`>#X��H��ԇ��_w�K����k�Hd!иB.KX��m�2��X.[��� H~���՛���#e�}U�x��.���t����l�P��$��MQ4��oh��4��Ekc�X8�I�q4����)S8��MZk���n����Ctb�2@�m�d/�9Z��o�[���uk�?�dɒ�����w�B�`>C��O���s?��G�����9�~UU��F�e:�I�f���k�!�iF =�n��Ɯ����wP�Ϫ��0(٣�R$ARCّ��$y���sf�!�F�9�`(�ҭ?24����nU��xƈ'&П� Ő{�3��o|�殫��:��ac0�q��1�� Q�?�l�����cǾZ]]=���A(�˄�zXt"���vY�	0L�(8''�nB`&d"�Z��5$gkD�S�U��JA70�U%�q�-k4�nh�[��Q"7(��R�Ը����6������M7ݔ����H`�c0�QΤ�񁁁�_�x��?��.�������>��*H����7�P+s���=�Jt&Yk,8P,���	Ph�|� ��1����iM��G	^)�
֤��Ͷ��l���]����kצ�}�����|t��1��8������������ƫo�ٳ璡���,�@bG�E#Pr�����+VYTdu��*���(�[ϗ�b�P)H����v�a�=�W�؋�|>j���p��瞷�}�W�xz��5�"%��u� ��||��1̟����mW{{����<���}SO��6��bk�Xn"����t Iګ��J�B��"�FH�n"�i� oh`I��8�5Ls4�L�{܁�e�_4z�o��ւ��7���`0�X���a�ܹVչ"J��݃��KJp��<]=�с_6��Dɮ��]�EsFg)J�XV�8:�PL���x��xC�����ӵ��^���}�ƍp�m���d�B�`0��(N#��U�e�ϯ�ڵ������C��9/�u����;�ߏ�}��_�`��`�c0��̊+�(t�,��`0�I :��`0� ,t��`&X���L��1��`�c03	�B�`0f����`0�$ ��`0�I :��`0� ,t��`&X���L��1��`�c03	�B�`0f����`0�$ ��`0�I :��`0� ,t��`&X���L��1��`�c03	�B�`0f����`0�$��n�F��0�    IEND�B`�PK
     mdZ�З�"  �"  /   images/2fc28fee-789f-4880-bf44-0d05ccb6f4b5.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  "�IDATx��]|պ���lͦl
!BBE� ��("�WPD���>���l���TiA@��R�C�	%$`H����f����;g6�\�}�B$����~�ɔ3;��|�����>�'����c�YB,�����m��ȑ#�q4n�


��������t:�^�z0a���ȀѣGAP[�3������1c 55�;ݻw�e��p�(����������֭A��(��Ά_��j5�Z�
z��{��ٳgôiӠ6��	0` lݺF�)i����&���d�$�k4�H�D�
p���3���u��)��h���%�}N�Pd�ܹ�vӦM!--ڶmV��L����*�:j��ÇK$`�hҤ	ܼy�2m����޽{�" 	��y��Ci�Je7�!�'FI+Y�5�e� �E�D0����E�������.��kҜ9s`РA��O?�/��5j���|�2���<&22r��H,\��-��MZ�$qD��bA�6Yؤa�s�b@Z����q��rmF�}��+>s�\�t	���WQ#�`��{�n$`�i�9�1X�� $L�	�=����D��-���K�121x�ID턫T�q�XKd��m��|5B����!>>	����$�B�,Py�Ɛ�yx���9��
"*5o#S�-S�i��4|5BH۶mP�ʡ�1D6I������2�c����I��)���ʚ��Â�Fq:퐙y�Lj�0��J�������&L|�<C� o"��X�A(wѡ���èB�X!22�B>@��)��!�=�c�<�	�́7q�%�+�0��
�:�N�ͣ/�Fa(~Jp�}�y�~��=f�<m�N��<���Uަ�����?x�c�d?"��
Ë �D�B+���2�(�f�^.;cL^�������Z�1O�8&%����K��#	R�$<�IĀd�P��V�o�5E�jF�DWN�&G��%m�i
pg����&S�v�Ӿ�n��AG](|m6KT��x0M2=BC� J*%M��B�KE{�Tt�|��U3��$����� ��W���K�H	�eW�e%o:����h I��w�˝?��Q�x�n�W�%,&�^e���	!�Hc��ӨBH�C(-{�
��B�WUjuo�Z�Q7
�=�6��^�3�[�RS����C�����;
n�FGG�'Y������0�?1YUѦ][ i����%%5�YɊ�_�<���6G^II)4�(u`20.\,�CC��̙,t��^�{��ܲ���*���ˣ-�صP��x�Ha'�eڴ}�9sYY8��r��ԝ8z��={�������_/z`[;w��􂒒"8��������;&�;�����;��E<vBX�E>Ѝe]����,<�^NNN���,�����ui��#�넅v�(E�8��%ة�
��.�&a��d�8��sy��߱ ����1��q�b�
(+3fx����(D�H
�Gq"�(�\��U<~�.�ȩ�
%ج{L�����A"a�������;���_��9P���"o�g��BRXu�_�.7}��<�7o�,$��$x�@˓��O9�s����P$�����m��<���J�$�G*2uyL�.ڦq~3y�d�U<VB�z=8+�\�i�\.��c�a`�BQD�ٕaau\+W����|������^���&�G$���	���x<9��]�f��/^8���JHqq1"Í�o������l�F+!Ţ>U����/,,�����l���6?�>]�����-��eJc�e�"�%��&�-CpP �g����JNڐ{�EC�{i&��Z�m?"�sN΍//]�0*9�	4o�III�q�Fi:Ў;৴���aΜ�0z���駍�����v����bM��x�!JNՋ��_�c%$,��1%��x�h�;;�\�J/
�G"2ILz�Cכ:����6o	��޳l�rxe��W�-[�]II	�)��$%%��)��p���<m�WkZ��́DIP��h[I����g- Maa�!g���_��{��
�	mӂ(4lѼ�_������|���3���&��E��/�1"H&)	H��
�t�!'����s	��"��A��A��Avt>M�%��EW�k��{�� O����V3@c�!&�w��
�	be���0�g�Q���_�UU��:�=Ǝ��?Q�7�X	�Sj=�K8��;���8���XD䔱	�f"��8�5��8��c���*����xM2+n�
�qr�w�
���ѡp$�q*r�U�wK��[���%g�G
��Ǚ)��O�
� ���!�_w-,8pȕ�k��H��<�%?���*�k���`B���[�UI��4�O�#T�0�<m]�~Ƕ5�	�k���.H��M$'���v��Zm��]1�����6eXs�~l��,ަK2}��{�x���2���`4��ĉ�(Q�*�'�BxH���؁cAc"<��ʬ[7���>Lއ��9äȕdobP�̋���JD���۫30�n`w�t�%a���$�b��"�L�M^�>|�<%UFUm@��aa��D���PRo���X���ݻw+���M��MF�Q2]r���z����� ��uc�!�a����i�oD�۰ �~����y��`ӅL�[s�?���y�6j�,ѳ�8�+6`��R)"��#O����`1)�o|L���Xs�_i�2a���)����By��I��ʽ�!�-�;�ł�I��ʚ�}�z�~b� <�M�fpU�3fX!#Y�r��a�͖����oə��3���,﷫*���u�1B��h)-=ø�+z;w1�`q."�xL�\�~-�/O#���	��r��I�S�QY�EH%r��,CY�����y�\����ZP�o�ʃ[r��ۇx���IԔ���-�	i����8��䜣jrW�N%���2Yr�=�+9|��?xFg�0~?@ʜ�y�ޯ"`3����c����ϓ�x^db�����tOL����&��/yʽ;r��3Rd����|oT���_��"@<).>H�z��k�8���%�K"��{#2!{�o�����QHt��=��!�R(����#	��$HV�����;Q9^1s����=�"x���f�x���L�i@� �L��	���'�<覞����_@�$�n�.'"ʺ)BE��Su��J�X��:\9�[qT��	)��16��w�r�HI��9��Ξ=��GQ9��}����f��������j�f�r�yJp:�Z�ȵm\�M�ɠ X��Jك���d��D_��O %3�;R��
�e³I:�Z��cnF��*�2;$48�d����W��DFFCR�d]��\����f����i�)-h�"�fw,,).�x����;��rκ�Rn�ȹ_v�i��
</t҄]KI�L���a������_0��a?F��k.3��CäTl�Q�b���V��N2����{����n�Qz�vk��ٳ�K�'�A��O������(��#��TE9��?:��� �9�޺Y��N���P������Z��/��_QQ1����&"�Ę�z[���LG

�6����0t�[���/_��~=�Qzشe���~w:���z�k�{Ymڴ�ܞ׽h_~�-[��au2Cl�O�L֓��5N��J�戼����������[[~���G����K!..6,?��d�B1���lkA�mD��j��C��^q������<���!�����v��L��#�YG7,).�q�1�o��51����NՖ����`���խ~''4>��	&<(]��,v�~2_y6lZ�曣�k�.�����0~�x�����8�E��F�ɒS��k�?L��w�3�`L>tΟ	�4,��4����Hλ�q.!���s�lx���2�vb��K6�}�Xܿ�U��O<!�Q\l�����A�I���U���7����R�aÆ�ss�-[�����K�~#�H���W�)B0:M�-��2N/ʆc[��v��!y����G�.��K�'���Ú{�`��x��tٍ�ܜ�O=�RR�����V��kݺ5����eYvk�.]\����sf �s�dF�!>��}�#D�������:�y���|ѡD��,v�C-Z��cL��g�%^�o�������Ñ��0&�>������G��7��^�z��P�^��q�<$0j��Хk'��� ����+)Az�,!2�]"������=!b��������SB��fş��Ӵz���c�u��|�٧��[�w�]��;v,�Q�F�*�!�M%8��R���-&K��C���	�1��X��2J(i�r�p��뽉t���"��UM��|9ˊ��{���?�7�9�-8u�$�郖�(�[��������hJ�om��S. �Z�����Qk��q!l��Ns�,*�R,�����n7ߘQ*ǣDSzs7==�O���=`,-UEEG� S�#���%�+Sg��	oL�6�;j-*���40p�+u�ZE�_t+X٣�Q����F��:R1 E6g�v[^��Pؾ}{e�i۵��m6$�k�.��R*\l�P�� ��`���t8��gh���yo�ό{�-6��,�7��^�P�)��zt�d��]���D������0�>�3�*B0���� (.��c(�84CO�Q�<�����zo&���=�(���#/g��=�t�����ǧ�q]�������~1�AH���~�jH۔�_\yߡC^���up4���G��9w�����o��S'Ҥ�>��﷕�ALL�C?_�#D*0
<(	0� 	���t:`DR��/5� ����|�&����JU�]͛4jP�B��b(�]�Rf9׸q0ʳ�Z�'�R\�Ǳ��k~��>�|�����)o�	 -z��p���;�P�y�c�N0�w���۵	pXR�5~�Ȉ:@��x��u����S$U��"���2�̻�NmaoJ���WF�o�ٞ��Z��>'���M�p�5AQ&7?�1���U�6
�1P�2�Qt����W)�f���m�����?}\����6C���L�V��p<7�ͺ�����~݄�3�|��+s^�W��CҶ=���:BX�:k�Z?E����j-�S@ӖMa���>�M�q�ǲ��L����;�s!G�G���o�n����n��h=4R���BA�yA�mw4�l.�c�	*�j|���><�%g8h�(��v���XO������ץ@����H|�) ����u�X�E�~�t�Ȧ��C�����Z���Hɤ�t׸\ɻ�2�5bX1�{�?q6LC���H��:"��尽���!�a���j��;]��Iq�S*՗��ڮߗZ�o�4F��m����E�8]�S��~�� \%�i-f���~��A���Q��Ϗ��ZE��=�ьY��k��;N6�Ϗ���Xp+�/7��E"O�ګ����n�u���[����C�f�t�4��:��Pv�&���s�B`�X:c*��85�Y��GB?�n0<��b1_��?X���:��fa���5���������^wI�l����% �>�7�k!=�������9{��GJ�$r�x�g6��[f]�T��G�
T@E�pa��걬����ҔR[6������_C�杤v_ښ�6�����v.�; (�F����Bȉ�?/���l5E�{tݱ��5��w�7��k��]�N�C;uH����X�8�yؓ�a����"�/-���2BC	��v�o��.d��ѵG��:�͝@��Edk�!Ҩ�a���5i�d��`:�~�>V(5г���MZ�ө>]g.}�v;\�������a��qW4�K�
����w�U�3�*Bnd_��VM�KJLIQ*ꔒ㛗���jM�]�F��?,�Z�,��j������(�ܻڶ�]��A�>}�i��YZ����Q�0�J}��R�Gd���u��96���_=��1�L¤�fgq��K�
'��j��W�A>��p�芨�2q$e�`�ZI��e�A���C��A&jǱ�h�"`7�Y�����xy�^Xߩ=�U��G�3���~](1�H��)�Kz�zW�S~�> i_�"�5��X����[�)EH�`�izQ-�
�kn{��nU�5�Qڸ�e�h���/d^��Ȑ���+���a�Wɸ�����pȶ��;�u����|��
��F����j}�ZCH�g_�^�R���8Eɗ�۽����^z|��ݺ�s���[����+}6����}?">�$'Ah�ͥ�]��U�JJ�EԭSO�^۲�~͠:Qk����;`l��C�Z��¯����j�YO��w6�$��rY����N�f�;���EZ杖��,���QbS?�
ǽ	D��%�V�vV�<�>����� /�#���������4����b�oQ�IX��p���j��1Q��m�.cDL��Y̓[A �l�䷿A�ԙ�g�VBŷ� i�.�1�E@�j�Ô2�ʭ��Ú����VTr�'
y� -�.'{��Eh�H#��*�>�:@KP4)�	W
j!'�Y !��2�i@C�$���-Bװ�W�1�� ���H�®]��x�q�aѢ�pe�x����!ڞ@a-��
2X��Kȕ݇�����*��;�	�� ��>�)~ٴ�8�:��(�����yΜj�o߾�as�(P*D�3F;lv��L�U�m�~ҋ�j!����(²(�l���F�����k����.7�M�Ѓ��΢&� ��Vm����&��^�Ɩ��I�4E�1����C�Ν�:Q+ �:�ך+�^ۻϑ��K眮��^����nCo8@�u�3��n7���j��U����yaaYq��R�����N_Gd��Q+�^�	�d�m�Q��������v~�X��x�ϋ���(�Tj�*���՛����'��/f}�*TY�B)BQ�[k����V��k!z�K!�h�p0
&T����`�_'	�;���rXxL���5�_w2����YԨ`�/��{?�g~[��d&�;�(^ �(���(�J�����Q+�i��;wOӅj�n�'r���,�,��s���\���҈�ϼٕVN�3��-ugM�.=|6��4hh��9�;�	�����NpU��	�����P+i��l8�=�
�����z��s����.�]ο��S��=C�{�JEZ���Rأ�E��}`�q�����j�0܂���p�R<�����"P�� �Z� =���֭Y]��Z+)?�w��S8����QJ���Vd��hN���i���B�M��b����#Պ���d��m�:��x;�A�_#(�yNe�����۷�ݦ{/+Y1�X��l�bc+=A�h�jSxh\�v�ڟ�V�o���k	WX��H�)�����´���d\,��r��=s��袷��99�$�v��3leR#H����| �������a�w�Ir2��<1��Y�y� 8�ܢ	D�t	�<�`�����l�bX<'���iS����Ѭ�-��
B0|4�O����u�k�z=�n�//
�M���L��*Z��plJ����Xͽ9������ߌ������ơC��Ր:x80 .�;v���Xm�jZn�'���I0@���<��	��ϕ#~�7�n�R�s���*���#�A�?�����o�~�-
K��;*UK�ә�b�O����q#'�� �f��Q���3M��QZ�Σ��.�Ա��Wvm�.��@��
�y0~�DHm۶MLb�w��䧺J�+��P�H�H��?m��N����%��N� �gʌC�TE_��o�?2lK:,��,H��,Sx�*��_�������}�xM�f͚n?�´���A\��_�����.��&�ز�w-3�����J�`�q�I����
�'�E�n"��T���"CT��N�h*�5<�u���"���9��w�[���k!X �zw����j��~�}���d�,��I�_Sk?9��88�%]�YR�mFi�P�c�Qu�׹"{�5��G��:G-���!��Бv/�4T(N������#ř��zʅ�^x6#bV(���CTh�K��wtݞ�T/����?ڄ��ZCƐ{`u�xhz���Nm�l�����r�_ʵPN��I��OZ���Q�
DruVqQ�?н�R:0�����~�guBd��B@C��"g��:Y*�j���J��4}ԩP/MI��b:w�7� ���w���;a��Lx���CF�"k������܏ �v����!��vX��d���ɾ�:�a�r	4	�36"��qs�+�9���&�X��]�]6�b�{�7W̳�8w�n�u��
r��Gý[w �n��S� ����򌵊���_���a������ 𻖛^|�b����m�K��v�򪉤28�f�JUk%E���� W|o���O�
�1F#�	�"�v�-PB�P��A!`�����³�z�ɯ2a�c"�����3�-;m%��Z8ĭ�N��޳c���/8L掂�ю��"E�4q�����=���0��Ӱ��mp�M�����5ש���[H_�
F���4㫯�<�g����h4x���ѷ��vC⵫6�ͱ��t�Rj �����7�<&�Q�����7R���\X�b�j5!2f��DZoڱ��=��h7s�)�޹+�z�dN����aҤw���A�������._)�1��Q��'�	!>��_�1��H    IEND�B`�PK
     mdZ��Y�kW kW /   images/9bf2961f-aa36-488c-987a-2819190a8ab9.png�PNG

   IHDR  �  �   �ֻ#  0�iCCPICC Profile  x��||eE���6�G��y�]�$�{�R�f�IvC�]�%�lv7��l��.  ]�4\�R��4������I���̝�x����/�}�Mδ3�|Ϲ�^��3��¹��I2o����)����gu�W���o]��z����-]]	~���{,i��G�i����gݙ����a1~���a����_��B��'���u��Dc���!z��G�w<9�����n��oե��w�vI2n���ŋ�d�.�4���`��Ҽ�\ ��3�͜�$�B"��K��>�Ɯ7���9I2����ó�d-���׽G�5{���69�L\Z��~���ӻ��ĮU�2֜�ff����[��?8<4�u�d%Ӵ)KӁ��X���L˅M�M=M��K��n�ٻ{�e�'+��IW��d��5��N�˒f�J���֎�5��׭���`2���P2�l�4�]�3�M�^��ɼ��gI�Ԯ��T'~{\�s	�Y�ѶA{oR,���g����u��e�C��,��@����jM$=	�Bos�8}l���-!���Ƕ3/L�����}l3%�&�ڗǶ�:IV_;Ink���6��+%�%[&�a������S�s�K�k�ے�'�W�ViؼA4�Ұw��g4\��P�k�V���>�Q��zbte����|�3c6�;��1O��t�̱W���8;�q���J�W�����/���W��ʏUX������\叫v�z�j-�ݲ�^��5�X��5�\�{k~���k}����[��u�X�����{e�C����ڠm�?o��F�lt��{n2f�k7����=��1��/&_����/�N?����b`�m�|m�k����[|��m.n�ӼCm��{_�Kzov��� �s�^z��Ӷ��������x���h�lҭ��N��N�l�s[��׏�咎�:ߚ�aW�K�/�y~��sv�f�{N���|��S���덽w8e�s�����<�O��s7�/|zx�E�.����6Xv�A�|�w�<����:��#�?ꜣ's���vܣ'�{⸓.<����O?⌉g���Y�t�%�w^��Oλ���.��+/?�ʽ~�r��k>���q�~9���o�����x�7O�y�]��s�}'>pȃxd�/|��O6=}�3>���S_������.�m�Ƥ�v|[����}������bE�W��h��(�v%&6�6\7j�Q��zc�L��^c^{�u�ݸҬ���/�|s�U�]���[��5N[�µ�^��u\��뽶�����č��x�M�lz�f?����ˍɗ�0�ib�ӷ��ղ����Y�\�ts�ǿ�B�f�o��j=����6n��W���~��w��k[�tj�E��k�s�Ǧ���;_��&�sש��u���v��;~��3v�m��G���=��G��ʷV����V���=u�o���E�����9��p���z������7~2�ʢ�7-�n�.��y�вesЙ_򝛾{�!����Q=R5�{�=�%�������?a��:�ړ~q�\u��]z�O��3�=�̳N=�?:��#�=�����%?^�����h���t��Y��v�˶�|�+��������磯�\�ε�]��/��-7tܸ�M���yѯ��[O����/���_��7w���;����w�q���|p��{���x���=��C�=|�n}��G��叝���8�O�=�詽�����gv�v��6���ϯ�¸G�4��[��^]���4������xs�['���|�w?����o�����}t��ϭ�������5�0j�QG�zg����������m:��f�?W��r�*��z�jǯ~��y�Z7�}�:����zoa��m��F;n��&�mz�f�l~G��/���q6�شŎ[N�j��~��mNn�q��k�|�����9�*[�[5��*v�m�����m��ܡeǩ_�v˂I���<��m����)���|�;�T:���թ��v���e�w��4}̌��M�}�=��o\��_�O�~c�����͜1�?kh��9G�����^?��yO�}a��Û/b�ۖ�t��pܲs���~�;���CW>l���mG�vԜ���Qǜr�y߿��k��儻�ȉO����ϟ�ҩ�����o���3�=��?��}x��~pއ�t��?^q!�xqr�'?}o��.�å7\v��'\q䕇]u�ώ��)W�uͅ�^y������nx��'oz��/���_�}��5�^�c�_o��-�ݹ��������̾w�}s��灹�~���y��?��	����S;��S�8�O�򐧖<=�������.���\�����~a������}������m�^�����ז����K޼�k�y3���w����Z��ZN�����㙟��H~���0�ἆ�G�5���j��c��d���4n�qo�t��+o��߭r��v��g�q����u�ڷ�s��O����W@���ԍnrڦ7m�Lu��l��K�&>��-n��^���m�mڦyRm�������������y��m�w���:;L�Q��e椃[O�|Yۯw�Ӕ���~}�]L�n�˦�h�-]�u���;y���#v�h����ܞ+���䷧������3��b���>1���/�ys�}W�����;,�Zؿ�~Ç-:m��%�\z��>�����>x�w�w�~HߡK;��K����Ǐz��c�=v���q-�w���N�wҒ�:��S�sڡ��ã�8��c�:��ct�9'�{�yg��?��U?����/���?�����K{��.?���<��~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW��U�Y��U�w������s����`����������cW?~����'�{괧�������ß=���z��G��������ۥ�\���{��7�zs˷��g����s軧���_7��������[��W 9,��Y^��$����]�bŎo'�Ӯ<��wW�x}��a��r�I�����I2�KI"�a��g�lq:0Ǫ9.͹�g�G��1���)Ã����&��8p�C'�]2���Z�ޕv�[�$#��j��::��&��F�$�޽�{_3�m��u�:�����W���u/�� ���};0{�^o����+r�����)E�=�?�Ư�8>=����z&^�3�"����F�6�������п?Ϳ�~��W�zF?�W�3&w�o+��9�v2� ���z��3��i/VJ����e�hq�>�[�P�"p,HH%8�����/����\�� �����p�e
�Ҝ.p�j�����n]	��%��o��?I怚���W[25iǘ���|�}��n����&��[S�p,B�2�:�L8�=Ȁ�Au��z�c&8���!O��e���7�} �s�;�5-�:��g��?�?�2�\�M#V���+i��A��"N��pmS@w���$%31����Bf$#:W������S�7i�D�� ����?�!� s?�4�@;��J�:�-��SX����e��|�I|�?o:��0� $�)sd���2���K�E�gC�vs������l�g��A�s�"��m��j�R��������;����2<{�ܹ����C{�/Z0���?<{pqu`N������Y������i��Sڧ���:sh���������޶��ƞ�����eUf���V�m%sՁFL=�����������8�����e��JO��)m}��;�zzۺ�'��uv�M�nۣh� ��;z��;�u�u�uU��L�n���tOi��k����=��mjo�q���Ńա�:K�ۿ�kxAS�u��ÝK��;���|]}�{t�aܝ��zv�6N����Lj�i�k�~��J�(�[OW[kowKGޭcz'�6;���Z'w�j�5�eƤUkk�k��j��Z��e��2uZwgKG��m��z���ї�i�q����ʌ��m��:�����aRwKo���}]�zz�'u�y�ʤ6�TİGGGD��=m'z�Si^Zm�oN�����܊.���D�ڊ�\<8�����9A"���k�fk��?f5?��Ξ*�e5�Xm��a�������K�L����=���Y���H�C��:ZZw��!?:���=nW~3��sw7d���������8��I��3��z �jc3���sڴޝG0u������Ӷ��6K�qZWo{'���	c��iS�4�T�2uz礶�>ld�����=U�E<����o':��JOKgW�S
��n�����I������������#��i��fZ����A?�c��V�2���'[�F�
+a�ҽ�U�jt�W���^U�ƅIU�����~�������8���R-2�YiҊ�����~�f��k�q����O�����2��~�	f��ʚf�[�O0�
Q1Qz��8(���8:���'%�JM��=����&2�9�Ei)h�V)�T���c�e�k<�R��<2Z�Hוl�����AGͳ*�]��(4�M%�2����*�)�s]iMs�Y4�q����u�r+5�`�Iiy5n�E�م�Y-�)�@g�٪�%�#�%�_������Ό��Ԡ<F�J�J��X�05e��T�B�)����U%�%�1rנ�*Nf$3T/�i%C8ľS�v�Y��̬#�J�F�-6bY�܎>K�MX�6�1�HJ�H�U��&�2l�p�4[��M-5�$*���NA�� �Ժ#��e�F���ƪ�fRn����I�2G.�R�H��
<P�C�G%�Lf��5!�$��j�x�י��5��56��@���0�)l�8�z�k��~��R�Sk+p
��Q�:��Ƥ�ր�{� ��)�T�[��^G0��$��e�TY�#f��p0ZV��dXOp�T�9��@H7�R)�F+s�u���I)@�����r�
$�tMH:�z��mKx��ž�K@�p�D�G�%���ʩ�%]C��T�
ǲ�Gs�Q6+SN�����~*���L���p�8w�9iwRA#�5f��	%�AX���K�uRKK�uk3if=�Fa���K��*\U��y��#2���"�'����&�q4�xMl�i���'~D�T���@+G�$ͬ'������ ���B�%�ZU8|,ܣ%ͬ'�/����;�m��>�"���N���a�dA�t����,U�YUX�ι�:�^��#��0�	`��FA�֕�0�j�:~(+L	��CU�q	Q��u�Dq,����p���?CGQ�h������?�>�����=PH�?C�_�?�*L���ʩE��;�:��*J���+58��Iޖ��	�LC�d/n6�FC��� \��_1�?�$U��N)"�(�4����@���#&��I]�)U�6�2�)p
P{سդ�������z��� ��
�C����{*qR�JM1�T�� �42�U�hB�TJ*t��b5,���h;0�\��Z�F���*p�Z�!�:�t�jx		,��a�`�FT`)��| �#$9bFhf���Q�ë�R��%ͬ'$ia9Eq˒$�TFp\W��a�_G�,Q��$�#�Ru怈�HS5�@)���76�R�Zҹ 2�,�R:J����4��pE���$"��(���p�_G���r��>��P����j�PX��zB�n�w��0#�8y���(�؎$�'�0��C
cB�"�R�iA3R�z�0	�o� $CZ�f̠�p�v�u�!p}�5�#݃[� �Z(|���	x�a�����G��j ,*J�d1����%!�B,a9�8�]E钬!Be��'&���2� h�LI�gD`E��Q����.8 9�([����
�Ԡ�O"e*O%� ��d:EG��e:PFX�i�s�a
���X!�F$�.}0�P�9e,��c}G�U!(kd�FƁ�C&������ܭ�#�i��)�%�j���QĎ��8 ��A�=9X�/ WS���wD<Eg9X�?	��=�ȭ�;

� ,���{���P �K��x�@*�@� Dq��<+֋l�>Y�R�g�C���	r�W �b���A`��SN���D૘+��()���@�vd)*�������� ��)���BN<YuT�Рd�Ry��Dq�jd8��)2��(J9��*3*�0#I�p�BW�,�(���)�T�j2�3G�tQ ��W��(�G,U��bV!����?C �A"�/�-wE�k�b��d�qF p�d�>0� 5����%�*V(��F�RR�wK�;�O��g� "wnX4�T��R��1+���[0��+#sQ��+p���W�@(�"ׁsd��Y�G&+��x�(@ #C^N³!X��
�W��3"��yXE�3tP��U��)����������TE���U%�R)�g�	�����
�е��=�T ,�ܣL��(��q��5 aԹGC�F���pl�{,:
�r�F�s:P�I�-�J������Pmi8a8��Sa���f%=�bIU��gR���TH�>����mZ�6��"���'��DO^�[���"�g�[����� ��(q�Q�3
v�%��(��:��eU�b`���� 	E>��C��YVG.z"�d 䒪3���u�3����w�(���Ѯ~(]-����YVK.zr��T�#+�����jmy�񫥴�CH)ὔs͚`z%+-'�@��`(�%���%�	;��e��ؓ���M�@�=m��=Y�(4�� �1�p�䝡�����KL$J�����մ(u^2@��)�T���2r`K���fN�3.d;��\�I:~$=��@�{�~��*�5z��t�S�V��9�jڧ.q�q���s��"�	U6��eSY���}�eS��)�f�)0�iKzFϔR�I �`��J�+S���@ rZ6�D�ŠU~8��L#��� -���/!o�ی��-[Pi�ϴq��2�Ig��D\���j�yY��y ���%=#A���i��Ǩ"CePڧ,�q�������T3��%
�SOU�5�& ����kAu*�Жt���U���dÆd��	dwH�H��Z=�Z�QIy*�Q0�&+���%^3���q�yBR��w*qpNz�KӘ��`S���K2��Pt��A�����OQ�_S�q�z�(iNV�M�$&H	��1
WlDO	� ��L�Qqr�Ty
��H���cJ��D�7��(�J�¸K�0�0�
=Ed�?'���4��\������`t�L%(9�qZ˭��P�3���� �!����U�'�g��g��=�}�f�P���L�H�EO[�f�����J�r���0�(sy�@���Y�t<�aj�9EV�

M��)���r=YfiNF�G�A�c��KI���I����U�HV��q�Tw�u�J'WyOn4��(K�cOzPĀ%H��H�)a��\�,���B֨W��j��J
o���Y���+�g�łzl��i�S�`���p�����e��}Ҝ��g�'��	�h
���.
�V�;r�p�6��fȊ���,3��	�
���~��C����2+�QT��/zR%�S>'Ҹ~H�����V ��* ����J	�J^�o�O���(��;�×t�R��ۢ'E�T@[2*S�(�I�"�0���#f�̸���P>MZ=DOU�3n�����:=Z�甔��2?�Isfy��V���<�8z�{R�R����K�?�ׄ��ZP}Or 1:F��q�TR��cq����A*0��W�e`��SGeR5��%�z䚹�^=�.iĞP�Y�F��SN�9�O�}~ڛ }̃7K]D�H}��J���(!��P�	 ń�"]D"l�dIt��Đg�(Rq�Q\d�V�ʒ�BfX[
���1����)\�t�����vȅQ.H�o�,�Ӕ��� ���'J�����)[�
MȨX.�#(�ڼgF�L�9�x��=�|�t=��BBz�������&�bR���a��F��q��PyM
�i��!�	I��F����pʤ���<O=	�iQr�q�����N(���)�)���Y&�
27�dqѮB7?�����C���
۳����ڭ�O�[��Mb�rÕMVm�o^�y��Ӽ��c�y6�u�yVF���mD�̪��]6���EP� ���!������&z�Dw�4E�j���9-��`�o��yCs��1��%s�-j�6��=�r�VYrIR�\�����$��uH����!��-�G:^�g\DR���ݓWJ:^M7��+i�Ƚ礥��@�x���8�Z�*����ע��b6�K��缔���$2c�tňx��G{�UѩOZ�	��2�-����Ll�HCT�=�����jEh1:��N�|T��2�EhE`t��������9�@��9^ZB��rFO�s[�/�uG��J@�@��Μ��;��?1��N=���%u��RbǫSzt�Zm�]x+��At����n��A� �����,�W�7;���D�I��'qX��E��}+��n
�:W#�V�zU~��x��|H�HԎ�~rAѵM/�@��٬���Đo�n�1�I�9?��x^�$�Z�6�df�r��B�疛�k�I�
z��0������9�L�d<�D��Gb�\�	"o58='��|7�e���,#_$] �����ߦ�3"�d�9��7$��V�$�~�5Г%��*52�Y�u�6�p����,_B� ���U�nЄn��x�Q䭈�~��":Jߍ*z9�SIתa�<�$��|~!��f�i�Pf<)����s��]�kuY�$N%t�����Bb�0y�I-�9�)�r^�?^�V���Ҧ*��X.3�^��`��ZA�����r�_�s��z�Z��yu~������a�s]�ru��_A�xA7a�v�㕩7H�D~�#'�)4]��ym�g��iH�Ck��Y�n2o��o��S(RɜW��H|84�TOB�r��(Z�V#�
$g~�ty]z^�_�r��MV� 	�)��&�F�DM�9'�nN�y�5�\!�N�<
��<	��K* 3HV&��|Λ�f�ji	��6���r�Z%z�@ʠ%�J���7����I
���`o�\+�_�� �K����V1(�w��/�$�c��"ZAx�J2+F��+ϋ�٠.ጵ��S9�k=/9k�j�)�u� (�t�d^��N&2?B�+���
}��a��;F:Mu���v�c�tN�:��PQ&���E� �˱��@������q/�\x���>P+saϓ�z�D��܏�è�U3��PH��IN�]�[\�g��=L��K�)q��0�g�,�"��|	�X�j��_I����\�X�\+�i�z�5{O 2�^�"��­	�2V��~��� �e�_:�˯��7�y�,d�ݵ��D��e�C���r�*@�6tC����C9�*0DAfE�������'����ޠ�{2]|��I�HH��
�L���{��/�� p Y�ܤ�j�N!�d�y��t��n2��0L���u [ɘ�![|΂yO����������0Z"���D��x��0�W��đ����0p�և[�ڛ4'o�<bfl���OhE��yC�@��Z�'��1�GC�8
��{.FW��-0�7�HN�7��Uy_�#��Ⱦ�C:������EuӬ yȬ8��a8D�'��&�V�}��d�0}7�9��1�#	���p~ǰ�=o�a�՟0���1CF��/���{�2{�~܈ahZ�Ρ�2�Z��1��7&�T|���6�WO��er�Y<���_ʲ0��>BrJB��"��xx���ӄ���[`(��a
S!i���+)��H�׳�a���%G���$6ă�D�)Y�D��8A�q#��p�ޭ�L�ԑ���[`��F�{؁��WD�i$�QyI�g�y��g>nR&�]7�����Na96+��n=o�0X:��v�]<� 恷�0Xm�r��y3�yC��T�%|�IY�1t�� �t�6�,b��=�a��>��F�\[�#$��I��ﱧ�BR�UP���h���-0��2��T��c1��[r�S�1kU1�i��R��I���1}އ$��U�5���ɽS �¹�"�z#����,���eIoC"b����Z:pR���E#$���J��] x�*"��y=�T������[`,'�E�	gA7e3�[`,�ER#汧�F�'D �O�;�֟E�0��4��U����ED�� w�n\i)�-0]m�NL�B��)��F��X��_*��AF#�_xCY�&z��-0�>�f�e����GɈa����̼��TH��AF��2���T�j_ޗȈa$2'�}���|��g2b$����&�t����0HWT*�$���1��a\��x�g�"#������0U���x��H�UэPYNbX��2b�n�R�Rg���0�"������K
�y�)�O�%9J����YDC�\�NC7�9D#	q�@j���F��
�xT��XЇ�a��yX$\E8!����1"w�- m�:�ce1��Oɛ@Zx�9��FRu1LL���I�fàՆq�����~܈a�¸D���G����d�0hաbZ�:ݤ�k��R�nP�2�𵷋�a0��A Ï(�㐊FR���`��i�3�[`��S���5ؼJ�x����JB��`��U�0��/sOʀ�1�J��-0ZC�H���С�i=o�a��m`���%�>��������-�'��W�u(�[`�����w�i�k
*bŘ�ABk��MK_�P�(�Wo�
*�}*=��511}ZW�����*b�L�+�����n��T�0���+}���	0��uZ1�E�U�;���>`�y�(�{�!z݁��>�Q�(�[�ިXx����1���?�ʐK��k�y�`AA� |�Qt���Y�0��3�a�*t=bEwȳ� |ȧ:��Q�F�9}(�=F�1�k}~���xo�ȭx�F�3�!X��Ǫ�a�e!��A�@�P�V� �����҆ڕ��ޗ�A�p��V|mEG�+}D媠}p+��a���ح�礦˙��FY�@א��R��ۦ���D�=�?71��k�{���)�C�atV$m��R+��:b
�,�&�&���ǩ:bڭwx��T���WG�黩�s�9i����a�d�^B^�C�<>��h�SAPT��"���k�x���`��l��?�À�{��X�Ky݉F#��O�#���5D�"|2K�T 9=�p��`
�Y<��O�Hn�`
��%@g��@執�a0��nE+���Iz^��FCS���B�J��a�
5��M~M��sވa0E𓚤Zu�Y:bLa}�Hw��,��5DC_�ࡄ�¹�}~�#�q�گ�(N����y7T3<���lz�c"���)'?�:���8d"�A�

Co�2C�R¸�Ak�{����5�bW�G��5T$	�E]��-�뺉�Z�Ã��89o�a���!�׀��͛�a�5���-OZ���Z=ޡ'����%��1�� a�n����/��a{5�C��X@Z_G4��W���W0o"���~oàU�:�!�/H�k�&bËg�=4T������pև(�:i"�!��^ʇ�� �L�0`Pa�z� ^7à5�>�X�¸:�L�0��Z�;��ri��Ɛ����4�<7À�P�pB*?,�[`����-��GHz��kL&b��3���6X<��g&b�{Á��C��x�D�PP!'�q5�k�&b0dv�CӰc��#�1�e� ��]<\��+11��Z!���b#o�a� ���z�J2��[`C�)�Y��z��o�0�M�c f�&�k��+ۈa,}Q^�fC}�����1P�!��.Z��f=o�a�V�<�����]�����{Ɲ3�!7����E1��a�p��`0�c�����Bɹ��l�0"!B
̛��/����0����o����(��2�����xa	��q��_o�0��*�W�����<o�a,U�Āj^�ع�b#���)��R�y%���җn�7@��Oڈa0��
2@*��5R1��uK��wA��<o�a�G%����K�d��-b�3��ᰃ�4�x�-0����n:⃔<&���%�;pt�͇qrPao�XCߐ�I�t֕�r��Xz�x���[��Iϲ��w�Z,]��֥��Rw�$�XRP�Ȟ�   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �    �  ��    x       ASCII   Screenshot7�o  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>946</exif:PixelYDimension>
         <exif:PixelXDimension>1274</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�g.  ��IDATx����%�u��2�-�WuW������0� HP�HQI��l�lю`�#���/���P�G�?9vXV�"E�C�@�$�	�`гO�L�Kum�ꭙi9��{���w+_�2h4���n�\o޼[����4��`�)��ˍ�Q�>��ۣ~3+���3|��5m�LZc�Z��[���~�^�z�HG�^�f�_Y,�`,�/~p�Ho޼.��q�Ʊ/��`"\g�bl�tye�HO�zR��;Eڌ�E�ĉ �q� ���������ﭝ�"�F���)閤�N���ߵ;�I~�=u�H�g狴�`C�_�t��s�rM���w�^ρRnss�E�Lf��ݔ�q��N��H�c�tz=&Qf��ZY����V��R��]�=�����9~�Hy5[�oC~����:+�.��N,יdM�:�t��X�g�(Msau�I~�V��?8�}��ø�~%��p��+/��#�M><��آ=�~�*����?�ѩ?��c��)K���I��=�ⷌ�xT�ic�37��q)�q�=/��J��<���==E�o��I�<�׳��|g��ND��ɯ9n����g�Z3�����,,����y�U��i��b��M���{i~�Hg#�0�)�7�y�^g���Ƿ�xv�����aϻ��}����^>ƚ�`��,X�`��,X�`����ۏ̋�,ߛ �k�ɪ��\W���z\�a9F��۰����ۇD���kN���L�G�&yg2z�#7�[�1��"�|��lG���������ٔ�������ʒ�\3 �b���t�?��X�GJ�����g< �ߣ�����W�n�ڝ;E��������#!�,�e�\�yO����O|B��v333�q2�3�_�R��k������o�i*�?|�p�=~�H�����Ŏ̏��Q^�D�O���9>ɏ,ⷜ/ͥ�F(�q&�Ʋ~����u��;���F�!�+u~�y��H��O��OK~g�~�Yrw.�Y/��F��ے0��z����<��t��_?�y��}�K�YN��w6�����$�9n���+��p�Aݟ��)?��.�8��Z�?��L�o��$�r�r��;B��G;X��H�c���N�6@`�)�:�vK���YM�G�>��+-7�_>�w�%���8>pz�`��Y>�]�cb|i��XnL���|$�>��a��$'s縍\R��$#s2�Q41U�4�
`i��s	&Fw_N�T4���>���3Kg���j�����/���>�|�V���%|��'�Z�>j�ٟM[��<|\F·c?2/��,X�`��,X�`��{��G�E��1�5��/�[L�>y�R6������Q1Aa	�{���ͦ%�u�ɔ�Wב��Y�-��<������&�հ���U�8H6�Z[����y���B
��m�yh�X-kK�+8,��=�8Kn4�p]��hB����|$�vB�]�}�H�LS=�c��ոK��>J�|�|�6���i���kE�8/�~M��DɆ�XH��]��nO҃�BB=*�_DFdA���7��R2f~]�3����1�7���m�/�w{��^#ѷ��N�o�Z�`g��\- �b�m5�䩖�%T��Q�7_{�����?�%�k�_o��C�x�?����>���C�W]�>��Oi��s���>�k����l{SQ5�䅑�C?��A���4x�&	o���Ѿ��k���'���L\m�-�L���E:/�Y)g�x�~��U��������|)���	�3^w�'��ݕ��`0r���4�d�q�O����;��]�q��rY��G�q�♖�_��A��q��o����%盗�&��.���H~� �wvq=�z��t&�]��.�|��t�����K���6�G����~��h؃G���#j?/��,X�`��,X�`��{��G�E��zZ�9�=��H��3�7���X�P1��ÛM^�����a}ضo-�},u�������N{FO;��L'�ǈԐ��#���v����9�ES֯��ֺ� ���EI���|�y3Ѻ��O�4~H�Q�.���(O�` C��١_<�h�o��� #mD�Umx�57�y��}G�����; 
H�5�$�V4pHҭ�"ps]�w:m'm��d@��v�[�Ġ�4�zC�|])?��,��.I?Y�G�*��@E�#�WjM�^k�%KP.�cw�z�El�˃��}S��w�����S�VJ^L<M%?q�����9>y��#�O��\�I�y�|���k�����Q7۞+�e���ɗ�Ԗ�1�Dو�q�;\X���o��,I�(au���J�	�0/�yd�ʊ�[���$�|"�yF�|C05�m8�j���A���,�a��ؒq��-7o#�I���=�cГqj�q���"�×��J�课�*2N�>�#��6�1�9x@H�C�B�//ʗ��+�e�D4���7)�/s�&��-�rb��ۗ�����E����o�v|D�ʌ̟b�0�IN���/���0�z�~.�n_?v�6u�����?���~�_�,X�`��,X�`�����݋�J�+��
�6�Yo�ȍ����K�H�:�����q��\Mj`<�aKN�Ѩ�������QM��1���զ�������-��\��7�_�s�Zߌ�.%���$��9)�q��c�"���V�l���G�p�]!�f�����n�X��?7'��h}����I��\C��q��@��~kD-���y������-c��\w�Mh��(�V����a4`�,1��䳅������[�^���$�p��3d4]x��(����Gr���� ��Q{����S�Z�zQs��^ۣ�n�����x��;>sǳ2�{ك�,9��gg�#�	�i:����7)��r�m����!�S�{p�|��|`>�>b�մ3ݕT���Llh���}��a5}|��郑}#�qQ�H~�tn\�����O�������`�~$���������-�Ԩsɵr��D"ƫ��ڲ��.��M� ߷1_!��Q�C��t�K+�9H2R����U�DSj����sGʵ5�>|���d���
R)G�'������C8�Ը%!�q�'s^vgC���y�F�^�v�ǫ �b�m�G$E:�l�jT��-�@�}X6�U�e\@��MM��-���Y��[�݋�`��,X�`��,X�`��U��E_%�,�HJDHA�`�fC<Q;]�XQ##��0�fV��D=qJxx�G���|�o�5fý���v~�o�y�z<O��SjY�2%��K������W�%��.ן����vT���<��]j�!�聴^�L�����8�����ds�o����qC� �Ξ8V�s���&Lb���G�#=�Ԭ)��y��r�z<!��7�i	4�Eogw��K�q�����Ls���  �5FC�76�=8~䁒 cD�-I����V��x�I����M�;��ݒ(������B(t: �K0[�E]�ש$R�,W���Q��w�O��"C��MF�=��艷�2��Arley���`F�\���%C��|UN��9���	�4�┄���ZԄ�41�W$^9��x����T"�5F�Nq_�	������;5�fe�ю������ �e:n��|P�?�2+Zd�6c�nz~Q�&��	Ħe�C��ޚ��\����'߳���:�X����[^���ZjԸc��n/Et�4s��Q�=.E�2p��_�rj��;S+�Z� �A�@�mfV�v%��ԎE���:�a�2�&��$��|����[ �7�9��Z���6����)��0��~�曇Ơ΃؏G��n�b36��������O�76e����Y���[ETc��JB�|����6�w�ە�l�D܀���r޵�B����|A����yn����w�yh���-h'湏�r��w����(�S%��<���㙖 ���������p��e?4/��,X�`��,X�`���G�E=������c�#��G �n�F�ZO<<�T<g;;]��x��2�$I6�GE=�ƅL�,�˶捴��}�!Q*���z8sj��,��[�:zkЈ�jKT�p3�j�1?<�!���|�jIƌ�H� 1�J�����4qԼ�c�<ߔ��fb�ϴfv�hsqQ�E�I@^����E:@kE����F�("I3j�\P�+�oj`6���E]E�Hi�5�����H�32��b~L�3��� ˚B�N��!���\����0%��$��?
�@�L�$pAV�lRR�\���F�l�� 1QF���q��%�پ�#�Jfa�R[HCm�a�Z��˅�0��^�DId\�d�,	<�k]!26��Ɔh��*v�$5�h$]���fj��M���r'�=&���b�D�I$�VW)I��j3pZ�?��k�����79�vHm��@�ɣ��v{��%�"C�-/.9��m0jdx�ԍ�|_���Ν���8b�P���?R���"Q���6��U�i�q�vx�s���ϼ|���~����db�I����Jr���%��~�z��C~�C2�$.�4�m���I�˯������Zf��f�%�s��o���1�r��"��(�$�H��8�`�x3-�k���!�J�Uvt��󓈴Z������;����ABn^�ۅy!�����2IH�ߒ�J��A@�n�-��uy��n����!4ss��x���/3�$�$![&�����ݮ�?��fd&�H"ٿ��d�ϬV�~A��7J&����-X���&O��w�{�r�s�r��5�zk���s�ܦ�>;�)�o��>��_^�~�#�u�G�˾��,X�`��,X�`��,X�z{�_�����{���ô����| �F�<��y�3�D�cE�%*��s�e^�W�j��*ē9�LI��	�GǨI�Z>��Q�,IA� ��O��{T�V�WX9��#H����T�C�+{���"	)��m��{�
J#K�6I���-���zK�E�����auC�:u�T��)<�ch\e֓��y��&4V��"�D�[����<D�KkNSF�etX��6��a%�G�:��̻^I��|����Q����#��z�zH�>��xI��R��$�pG����.c�OF�"C$�z��	�K4�ɷ=<+Z��}�2pCI,V�`$&�TQMCF)&i���@��� j<�$�h��vf���;��牠Iؖ��FTæ!�I{����Yݘ��w������3�Q�?\�"nc��c��(�Z�����~%n]�/M��� W�m�+d�F��������xW���I��w���P�-\3�Q����Ʉ~Y�<�4�!�l�x��H�q�6�!jU�|H��}m��"=}T4T�^-�X�e{�@���̷<D���gf��PV-��F7�tg�F]�l^"&f4��ە�r�j��*QG�<r�#%_�n��j�q��`�>�G$�AZ52�s �	�q�������;>��g}`��8ib�h��'��l�)�!���߭�o�Vq��I�s��:���f��s�����{�ԭ�<����Gq�咴u�JZB�O��rL�� t���;��y4b��׉qtK��fgdm�[ȿpsm�\�vwd��
)�MA���<�&1�N��8�i���te5�����Rs뛔~�Vq׳�K~޼|Q��`��D�d��e^"0���%����	�ʰM�_��"���xL�~��r�~)Фv�>W���|P���g�˒����MWΕ�O?V�_=�e�*A9y9ǹ��ZM�:s�+~A`G��j��.���L8��0���gv��=�/��,X�`��,X�`��6�}h/�|�}_J���0�6�U�W7$���@<D=x���*�Q�x|�NJK&f��e��F+�o�Z���d͙Y>��iF����ۃ�
	a~� ;�,KG�� �(\�D?5����4o��-:�`��פ[!^{��E�m��B�=.���Ҳ�OA!x���E���"�z�R���Ү>��G��`,�������x��1m�J{�ɠQU	��z���c05W6��(���K��c��s'MG$g{k�c�D
<�J���=Ǩm$"E֍���2��%,S:��4"d���ãN횤��z�pt%�H��D���b>c�w�K"��Z�^�$��$@pS�O��J;̽/$@�F�ν.[q3#9=͖ԑ�F4�Μ�'�(�6ȁ��Ʌ%6�u��=ޖ�lZ�[p~��{��Tȅ���/�D��'�?Q����=WI(ԇ۷E�pڅk7d|���~\������!��v�U�Ĳ5�p��r�j2Rc�	҂�� MlgԎl�����~��iǥR#��1o�]��1�����G����#�qm>�4���G5TA�|�o����#Y�(�؎�'����ZT���vc�83_<��, 	9%���EѯRrgG��^��mfFZ�����{�Ǎuw� �J9"�g��*����+5�Myj����]�h�T�4u�W�{Z��=�3d�w�L��Y�b���;ȲX�!7�v���Y�qO���j��$L�< ��Q��M&�J��D6��nW����8�s~G$�]-kއ�|%e4`�CF�oK�1*1h\OeBG��D$�Ϧ-�;�;$�0j@w4���e�vs��]g:Ώ�����|��F���UIq}��E����,�mt����ܟm���n�xֆ�jI���S���J{��)*�b��=~�\?�D�3Cb�,S��9��~���:��̒�>��$����ͦom�ĪT�ilڿ�����m�q\y��ˁI���m�K���1mu�~�7����f���K���6hn$/���XH��̱�ՙ�'��}h��t��`��,X�`��,X�`�{�/��%{F�om,�ΕM�l�M)� ���,���3싧h�hV��Ѵ����(���G£$����5�4�yC�/�-Kf��2���z�&k4�,��R�f=��ME�oJ�����;ޜ���N��~�>)�S7Dkh��|�JRC̍�����2�K}���U�!%�6����7�r��}��ϣWI�n*����{�������B�S?!�����AxWEt�c'�-�֓/��-!n��_-�g�>W��?�_ޗ���1��yJ��j�����@ҥ��c�5��:�N��&��yԼ��ش_��疄I�vG��f��a~* 2ɂ�|�=&� ��MF�%�Fk�!i0��NT!���	K�f�J��s��Mq�Ԩ�����}a�gyY��l$T$%I�lR��e�Ҋ�!Y4�6��j�\M�3�ƴp{ VlL����)������_����ɔZ%� ;r�]�_���ڎh(}�O��Ho�X��g�HϜ9-�c�]�[b깓�&��I�/�w�Hߏ%���g�,����DS���t�'m�:�D2���O<~���{P����	.ϋ;���\�4[t	l)Z����ϸ���OWru��j���Kϼk>·�c�,��y�7��Փ���Q��G��BBͯ��b�0j����vv���@�ȡ�8?�5c�8��r2iQg>���܂6�Voۻ�V%6�߱�#AA�6E�mm
�����@�{'؏W*�\�>�=D]U��m6h:��!�I�&A�q4V�,��X�H�q�ğՒ8� *�!�G���%�-���Ps�#�_C���0�	�>F��Q�L��K2��/x�؜��J�MIhj}�Z9��8���ȝ�0�:��Y_b�զ_Fhy�(��/,�;�k�e��9��}��F�ο�~/���twG�9�i�D�(�<K	'%�Ўp��2���V��k�{��ED-�iS�V�C��e���iyE��94 i�4$��2�x��$1IN��u�Q�'cJ��6:�~y��I��Y_M~u/�����S�hǙ�$��y'��Yԣ!�,@��=Pø��oM�K�&?�_�WM͚79�2��,�h�U�x�J̀��>��f;c%a��@���؋���Fn?W�`��7�c�2���7��Fsh�����Ӱ��.�������d_ ��,X�`��,X�`��{졿�#T�oG�+;⩸5��ɛ�Q��x��H�7���`?�ld=xz�mw�(����5ӆv��e_D4�yxvRx��������-F}��a��#I�hS1a��R�5��B��K�E�h�Y�f��'T+hi,�M��y�!����"�9ڔ�ӣ��r�5�sjr!z��Q��iE��W1=�V:��a+��c�G/?�B�6[��y�Z������J��w�z�H_{�{E���|�H�8&Z_�ƪs��hה��h֤;�|�)��g>��"��	ٷq�Z�~�s�wv�=��j��H�İ%\�E��'K�1�~D���s������Ők�d�����w�W|�.�F���#�Q���~�<���!��Q��x�3�N�ϖ|U��1q;�H�u�D������斧j>A����Yn�Hk2�m�q���FIJ�CS���X�j�R�-O��h��R����B�Qg��m�gԧ�����̦�A���vy�i���A���E��K/���ٟ)��M���[��j��V,�~�%����(�zM�����7���	��{�y!�c%X@P��S2�m�������i��n�K=�a�G�qV�Lv��|�^�}�@��`�c�ё�0d���J&6
lt�W:�Z�^j}�֏g8�QS.6@��6�����&����+��g^����g��3/�R���{���'�!�!�'��'��4"�Yg�.	�Im���WE��٧�tyi��!'�ɢ��f9K>W�!�+�M��n�#s�ѿvy`c�0�\;#�/i�p�3
�oop�<0�裦-��.	����!�4�� ��K�g�!�y���ko@�m�q5r��Zm�w\����(�u0����[6��J=漅$I�̔�#2�&��4n�O�pp��/T[�%�IR��Wr��Z���H�9r�AR!�����R�[���1jm.v��X�h7��mgy��:ٸ��u��#y���~��ѠU��s��cy����t��2/d�������n~\��rM�Jo`���/�<���?Z���y �c�3}�y%�������?[IGxo�/Zr{��a���t��s������j8����ܾ�kw�5�}�+�F]�~�F+6�ő�Gi���/���yhKϢ���p`Z���_���~��"�6���`��,X�`��,X�`�{�/���/p�b���!��֮���F�:m�c�M�xxN�1<QCIG��:8/�^\�ŁY�(ZF4��9񔶐1�Gq��ͺ�����ݱ���n�3����zg]<+�&h7�x A(�.h��*I-W�`Zφ��:R�D�j��f�Dw���g�i05jm��VC<��x�{��"N9���
r��x��|��j,�V�pP�1$@�$	� �1��?���ڥu���n��e���>v�����]���~SHן��h�-̋'�Zc�z.p��d�G�<d �wwG��S?��"���Q�����"}�c���>��.���O�8��Q̘�ci���,-��UM��}�����ܨ���гN<=�z��U<�9�����yR��O�%y�~����L4�LE�,�GR�Zu$���O�I�E6Jp���w4/���̍^�rL�?�M�ɔht�j���d�]n4�l�`-�ȍ2�fۋ���,I��Ҏ:Mi�J6�6���%�{���~;��{m k���4��ѷ��7��H�?�uY��yg�9n	�O&�JRfr=�F�P6�e���/|�H���׊����E���dP
����H� �_�|A���)��W�.�lm$R&G�~h�Z�J�F��ʌ���?)��$aU���ｸ~�H���rXP:��!�"�!�p�|���k��+�IO@�F�����	����=>�{o��1�h%2�����HϿ&����i���cF!w�5-3���{Ը����\�$ڔ�����\}�M�?ǎ��C2�mBKh����dYo{�$%g"�b$���tw��+CD�!��eR����R�i�Qg ����j���rI.՚�̼��p&ڦ%�b%�3�7�$=	4���7��ƶ�7�	��&M����B�e篞�7��}a�Nj��:�rq��|��BI�k�c�1�.��I��7���q�Z�DN#��,g�[����s~g�a��d����,5ݨ��KM�O��a��$5�����m�^~�}!�o]�~���~'&���i����%'���-ϕ��~���muF�B�U�@�K}f�C�(�Gs��ț�g�x@bYE��X���Ćܯk;B���E�h^�����j�U_�4�ߺ�����mQN-W��3߰��/�*�
�������ۯ�,E���8�LD�\ҭ��W�uyl~�H��N:�ԏN����>*r[��Y�h�?lD_�`��,X�`��,X�`��}�/�H`P��vC<	x�:�pH�5� ��0Y���(?C�a�KzpN<��?[�G�����J	�Ǣ$E`ϧ���tG:Д3�V��> �x���"]��u���6�����
)2����� �C��b�� V"��)t߼�h^�!h��O�"jQ��Uc�Q.�&^_��8}xһ��1ߍ��I��3
������Mh�U�?S�z*�NZ��rV�4�KO��F���B�~��oI�=D�42v7�>�	�ڄ��}�'��Њ��6<��'�Zb�=���'$����$�NWH�0�����v�}�_�R���W~�H��!����g$_�	1<�G���@�u�+���C�����~R��A�������	BC�у\h.A��]=�.ͧ����ѯ�?%�rz�=���-gP����z��=Wx5��ׁ�D$�BzDIX�е1�!c�a�_�$�xP~VK�祕D'��R��d�+�K�F�]�JD!!ѷ ���oo�R���9����q9����ʅ J�Fl�u��"j�4�VWE{�$������I~����=���I��R\i�1j_�'ǙE8탫�><��ʛ�mwW�{�Y�b��[B8�Ԝ�~��񤿅����xV?����N�F�$��7��^�ufp�r��m/I>��Խn�c˃���V�nub�R��d=|)��47��c����_�kgH��yL�'��h�D���ڊk�/5A�u��>u�L�D��1��Wߐ�4T�d�t6:�Ⲍ�W@�^A;����r>h7�.A�(�$�l?3��b'7��/J� Ǔ���/A66d^��K�Y��?�Z����3�d~K�����޻�!����x��De�#��ٓr�Ȓ���y5�8o���D�~/�x���$�Fntb������@VE�+9��Ő]�!xu����.�_�����zQ%᭹���ѐ�ņ��1�k e�����~��{��O�Ԣ�X?Rh��1O����<�"������E�l���a4]>GP����Ȓ�v	#ޏ��d��@��K$*����e�釵7 ǯa�/������x�A9g�O�s^��7ο^�yA�p�g~N��ޱ�|f�c,_ �</ϭ��2�Fx�@4_����< u�?�� ��7�߹����02����UHK�|�f��jHj4mOw��a���j J���o}c�cmF�o��ĸ@R�K�="V�����_Ra�j���,��I�������/�<9�u=�#��/Eq�l P��bq�!2��y ��Q*�mzc�?���Ȍ��/D���w��ڜ<�%��|�aY ��,X�`��,X�`��{������ƚ�E��}C<�#q�7F�L�}�.	��x���9�x�H�:-�ܩ%!��1�/���4w��[ow���u]�y����ϐ����Y����⁦����x��_~�H���E����oڍd�zͫ�����������Lj���ki2J(<|Y�D^?�o�-����g ���|6Z[�U�,�"v��:�z#hՠ"�mzF�75U���Of�/�'�m���xV�y#�zFO	�ސ5Kֿ��hQ��dI�!4��������=��=D�>�Թ"����uAc2m��Z�d��s멒#��+�#��c�^i8�c�t��4rO�D�GK��W��1C�[>i��v�zfT҃$�'�Z���}$MYK�U�a��o�-��v��'�^G
X�=�$4(�*�
cNov�q���E�⥇ބ笞ɓ�?�x�;��5 �<���=h�a��xwrio�M͍}�Fsg�
�C�O��w_�v���'� >�h��.��̭���C�d�xI��׮b��َ��K :�߆�f�F4�ED�B9�~N�����H�c�/?�c�(��!!�^���}��'���#ܙ���?�,���i����d1��K�l������3f	��C;郄f��5��0�%�|����2�����!����V�)w�5LM,_��#���qڋ�<���$%�y����x^|Fң�,5�\����H���8zgm�Y�~�ݑ�8��[YYv.�d����L������"}o[�d^ntg^�k�3v��V�H��9�ڑ|=q��"m��縨H��ۈ6��@�w�L��_㋗&*������K]BS��j?�+q��G��H��0Os��0��������RSn���G�-g����W��F��a�c���Ο�<��-�3SοA$%w=9�A*�1˝�.j��C���f�ER����o4���<���c��x��qˣK+���z_yV����`#!~2ԫ87������7���^���Q!�>�y?���+����N$'P��de��W��;���󻢅{ڠ��v�m����Ͻu��"�6�`9a;*	yw~n�]��M�:�(�l/	�o䤑��Z�����Ԓ|i��ѳ�^σ4w�6sַ
	o҇vM���Փ���?֔�j�ch�dmF ![�~�����¤���z�}|��Ǽe�'�k�I�3�q��%Jh㋢�$]�y�n?�����q{g0�Lw���c��/H�@·�����Z��s��i��}Z ��,X�`��,X�`��{졿裇a�������D����X��R��O۸�7�=�����O��������ބxH4��9����ע��޵Ծ��=m��o��g���!���o�����;R��R��d&��|�Ӆ@�%3�
�義���27�%�D����c��_(Izp���u7�d�f�FOƭ6��09H��u�����"�s��,���E:OO<�C�������dd�)��Z=]��ݮ��k׮a��������>u��"���Wq@�w�bܗ��qBS-S�V+�ʍ�;X�ښ�z�faI� �D*�f$���C�g�hocE��6��H�8�\U�գ�Sz�[�~S{�}�͔�[�(���G�{%e�$�q%h4F�m�\�O�Ԕ�f�F7V"�ѧѷO��Բ�G����h�VG��c#�x�~�>�BIr�x���>�zD���'_�����U����r�|\~��	7#�a�b�zUȿ%h�<(!ITj��c���1�o����wDunvN���#4�hG׮�O&?T�����W�s���Ǳ� ���VxW6���� g�&]'��+��GK���8s7(��� �s���!X�S�L��R��=)�hl����I<�D�tY泌�J"�D��H�v3�ٿ,.97��Nۂ�e2'��O}�H�����H�|	3�P�Խ�:SRRp���0f�Bl����%[}��}��;|���vJ�0Ze�ki�ĳZ�Z��'�}%��/CJ"Ռ#$z��w�	JFn�MI6z�)4����~u�l�O���M��C>�;%Q������wv�c��j�KZj��|�yUO���㉮;�^n�+	36�\>�����;���;��3�'��{�]�2��5�^o���u��@~.,�<���>&�n��-򠹜���GuB�%i2��7,x���_�N��q���O����=sD� 8s��.�}��<���k��3Wf���(�w�W&ڜL��<P	^�<��������o
��$�GM>���โ�����]M���=ZT3!�*���%������y4&�-��.�<��X/���xՄx����_�U�!���Z���y� 鷠����n_R���4gtn�����$�Yq��!�7U~ԓ��@$���Z���~	���gq:Ĝ�L�h��k��,X�`��,X�`���1�����~��x2޸}�H�����7�)H�h$Zc���7�xZ���> Q��-�0j��.�a�����,O��M��)=>�������|�!D�����鷯I��~ i��7����!	�s�W<nt��3L�Z%,��}I �hM��Ѓ���~<�g�J5I��(^n�;�|�Vz&ݜӱؤ����q�Gj������#��.�gνP�fŃ��s2�%+f4�MD�=xh�HI�GnԻ8��lB�͓'����q�݆f���l�)�?�$�+�59��*�O��zs~m]t�Ó֤�Z	�N5fb���6Y�jƔAz�]�/ը��?�g��2�O��#Z��a3v5�|=M^!�����l�1MI"�?c��y���fͷ]�淢���9���~��D".s=�JM�=���Ƚ����r�.����iT)�i�S�Y���Z��Z�c��t��f�����ǟ/�����E�ҵ�(d���Ǌtx[��z���w�+<$����nv�D�������Q�^|A�?���o��_zZ���!���ܿ�ٿ�~D���H~'���=���A�l6&���My[|����q� �@���V�������P��Fe;��~�$�͟%����TS��6�g��a��o�x����(<�� L�����6�8���hk��	�3� i��̸������ot�g��d�A����B^Z���׷eܥ�g��mɑ)o�6S$QH"�5z�$)����E���ߗ�8;z�HOM�H��"W�/���F2��Ж��xBRý��!̦��i�V�<����f��t�^s��{�G��d���H���8I��d5_s�e�Z�`-�3�����]��]O�C-��\�ɿ�Ȓ٘G0��<�|�e�%&������2l�MhP�����<;������l�l2�s0@�����
��h��B-a|�@��>��z2�9����.�q˽o:�ޖ��Z����v��cȹr<a�s��r�钄������p.�o|nyF�>���o��9b������߲�v��[�I�M;OV�sO4D{��^�$��C�>��aI2�Å��n�5� t��"]�9��m M�Ѽ��#!�{ �nu�8����h���g=�H)��IUԷm�g���C�7�nJ;<�X���s��yA:Z�x�_ݫ�/X�`��,X�`��,X�����>�l����j�G���L4Jet�V7�qA���y��!�����L�.�}�}^@	�*"w�Ǿ1���Gf{��0Q�艛̭���������l�ߔb��q!���/���"�r]4����4oa0�]�*���4f�;*�z+���L�#W���H��U�G�U\�N=��d�߈���}�C���)Q���!�-<��>�m���F�<*����Č��aӇ�Б#�9O���@��b���U�OY&��
1��狴�h�Ծi��z���"��������H�Q3����
�Մ�	�1q��o��T��͢�����Q�Yƅ�(c��ƣ���y��������WK��y�<��=�~jj���+�|�Ԩ���3�KT! M���Zb��������ȫƒ�rEf{�e�����x<W�������
`�|Q��Z��Bm��=�����7�i�a�;B����}\vC�m���[����+EJ��<�h�̀�nB�����;[r�g���w�лqC��iLmR����ѧ�}��R;jv�U��\���%�������$!�yH�^��;�X���jr�)3���{��y��̸���H�ƶ]��g��*@}�ŏ	�� Q�a���M�؟9s�s���Q��hVk5�L��M���1���!�l���|���"����EJ�ق�.�k$�m���J�h��Ԭ��픴��tgK�Y{4bw��G���$�l?g�_���-j�aE�z�v� ��&��^W�k5��~"�yB>9��Bƣ]�ۖ����b>2m��O9�2Q���/o8�f:���u��8��M�Z�8�j�5�r�<g��2�.A�yp��?��Sҏ�-}��~cn;��k�֫.�kSj��K�Ò�e��a�GT�L&�����h��bg��d�>���w��e�o����	5;Ͱ��>�8$�쁃��������J��,�<78��:������9��{��-�g�������X?�@{��vK�F_>&ɗ;)���w�"^��7����>�����8P1���a�����:MƳ�Ro�j������}���j�v�Ļgޡ�ҭܺ��S��12��ꌼ'�XR�ή�߷w�D_CJ�F�~1c95.����Cj�����:ڔq�آ�gg����e�jm���*�y��@�,X�`��,X�`�����_�ոl�OWM���t�c]�M�hR�MY���姊���|���t+�`����ܔ�Bݕ��Wo,����S�Z&����SѢ�\���;5"}׍7�������:���&��~�H�Itԯ|�+E:{L�-��y�x�Q��jk��������qd�4��K}���d��M|{_�o	����_����ˬ��a���-���|�e1���x���Qz��H�0Z���nA���,�|$��`TI������1r���2j��y� !�@ۏ�Aޑ���u2��{�Ӗ�
��Kz�"Cdiyh�1���~\j<�����?Ur�
j�h���h��է]�J���6SN~߾v�_ty�	�:4_Z�$Y����}�a�c�������k��]�;8�Wk�E�`H^Z(��g�D]�˪/у�xl{Z��B���k�}�xGm%�s۟����w�N�D��,�@��_���I��.�ι�$*��,���n;�"��!��++EJ���)!�9.�0����E��z�C�m^q����sw1��է���L�^�čϣ�%��kQ�o.�ZGS��*����F3ZO��ڏxr��f�HK���w��b�<Jp�$)�`[H�X�.�v�;2\��	�D~�*5�Ʃ��?/��M���M��lo���"4+#��>�h�-�K��!�-�Y�v�/�Qp5�/H��A����w{��E�C������T����?���~�a���A�����@a>�������XES�ܯ2j�eYX�vF��B#�F�6�Ԏ��{�1�_�m>Iر�t�:}.�KkI}ϼ�F9o�I�vl�����y��|j�t�����˝G�źx�}+ES��*On�f�q��΢�l��9�e�_���S��!��k8���g�h.�8��K�&�&�i �lL��w��|Q���&��h�G@�bgŚ�*jڣj�i�b�{�f|`�Q��<Wi}���-!^����:�e���R�������F�}�O7�0��k-`�-j���s[���b�~��9�=+�}���'e�8��Le:m�J�Vvsw��oA��,�x� ��J=���U��y�d�_�K���_�G���lG�sc$��R&����<��95�����^I>Z ��,X�`��,X�`��{l�}u�WC���sW|/G4 ��xG��D��O}�HOtD ����*��H�T��j�����u�+����h�m����ؒ7�[�βۓ7���F}�o^A�ER���c��"�>yD�"*)�>F�%_E�٧ˑ��4o�3-!�������j����$��"
�TEB�e�#��oZ��F�dG�=G�*�';�@;������~߈{��Qb�81e�Q�U��l���6wԎ���Q-U���@1�V۵��e�!z"l�`Ϳj������(C�Ф�5�5��C�A &��'�QM^��g��ѯ���j��z��Q�����\�G�l�ǡ�S	_K��_�&�Au+s=��zi� �tP���-�����U�2�g�a�7H��Ë�R�2�������'L5۸�"iH]"�B�-�L�r�!ͦ���J;���mԧ'O���ؾ����K6��Yn��j����Ð$������_b}f��ܔ�$q���O����]]Y|$:��u�zGv��^6�\o���n;�D��Բv�ڮ>׶os���簾��㗨��#��̝&�g�6G�#�2c�^Qd��V����KPR��	�=O��_$_�x�Sc�{:��Rc�㮎��;>��Z�z�_�������b+U0�њ����@�x�/�P�z�/T�ێ?f~�d��G�Z%�<���<�
4yܣ�hI�s�2D����q�<�0u�_�Λ���q��]i`8���\֒n{G�d?l��Z�:��vUi���(��ӧ6CTU�>'[���;P��^���H����s�-&)��7�.#TN�&�s�_%`��\ٿ���6��<q�sTn��"�Q����@w�i4J�����.;Ft��(�vG��9��e���әyl�n$�yJmF�y]�K��&�Cmϥ�.Nī�<��i�j�Q;��tH�]n��R{�2�kLg��y�v�)��d�/�;�{Tb#|�h6��z:z}b��O����`�	�O�ܭrw����H湭%!��0��v����My?t�{�HǊ6��'2_N�|��{"Λ���{��Yi�	�U�ҌG�ћe��d�}Z ��,X�`��,X�`��{��E�=:�S�.R��ǫ��@��⡘ŷӟz��"=�Zu26�g�od�j6�2�Pa��[��ڎ|{}}C��n!
�vO�2���KZ|�=�czLd�۽�Ez�D��΅׋���Y2�K��B����p��T"�a<�����f��z��E�o~�Hg��죸��,��j<e��h��f4��	�׽`n^���.<��o�g�b
賧�#�zR��UqDYO�<��p�gF��@�V��H�h\����`�O�U�k�Vs��I����l��#x�����bg�=���[$ެvOù���xC���D�Y��/�;�K��%XLvKK�
�άɟ9-���}�����qJ�Օ�S���!�L �X�<��K�մ����S��C��h�S}nT8�)J�I4�:�vs����X�u5�T�s�6�]����4��U`�w�%�M��������K[��s;�C�\��چ�"4Ѧ���w%����uG�hhz�5���aJ�Փ?S���W�$�4z�!�h$��d+f���Մl�UCZYңB�㸤�p4t����m-Ըj0�7��q��������ߒ��!3д�qI��T}|�r�ɳEz��6�3�Ӝ���g	4|a@�SC���n�;��u<�8�w,/��n�ۯ��[��F��d�W��|��K*����ʘ������rj���d���q6i�(�|Gw� �1;.��<���3��?a���y4�v҄v\�l%n��4�/0����լ�'.j[Q��׏��C��'k�@�X3��>�z%$���Q�u�-�D�TIc������C�*��Q���rO����sYOU��|s|�ѝ�@������:����$�ĸ�8�+Q|Sw^�#e��sW�,����sz���I�U����-I?��+Ezn��"maC�gI+b�X�'g(�lo'��bJ���iCl���N"�K斥�/���-�H����Eʨ�1�Pm��a�ɟ)�z���Ci/m}	�s7z�E��b>�U6�?�L��@�,X�`��,X�`�����E�}���z�=A��ѕ7����'��$_��#�o�V��L��q���u�=߻-с.������|[���4G��Dm��} ��I(O��2ʊl7��Gt�ݞW[[B޾-��FT���엊tyF�\yA�x��A��N�"��O{�H/]�����"�;���!*YTwc�vɫ'X��cE�Ґ}�`�7�c�nq�*������פu���׃���W��q���(=_��I�>�(�{�����i/�z��rZs/�ј���sj�4�|��P�i�G�s��V��G����g�$�.�2U�z<�'�T����苄�TN�̄Y����2`�ii-D��ͿJָi�)��%O�Z�SKO�z\�+i�;�K�*��3ܶ����_��4�g̟��xD�Jg��wd�\��Fu�1OԹj�Q���Hl1�6<��b���ٔ��ɛn�Y=$�t�=�C���u����q؎��n鱣U7�����4w�=0�Ϛ-�)ǭ,��]XM2+�|'*����@X%Tm?�)?K��PW��$��>1�m;mV�c�ӣ+1o	���%U����	&��M��GEc�����)��l����MR{r8�j�܆��b��36��k�h��*Ѻm�pS�D��d9��H)�S��Zz��%���4�j�	0�-\j<b||PD_%ʮ�_ֻ�P����Ch�Z��ѯm�]KtƉK|��+5���V���-��i�\.��%���K�yIĊf�����x���,5�8_���/4�s�=Ac���h���Ψ�F	�p�f|�L��#��%�خ�X�����~>���t�a*f�M�ڑE�,!�J��}��l�>|�X����E���h��=����)�k, ,��/l{���R�����ޮ�3m�7��J���oS���������t��?���ufV�����k�^)C{G$�pj��C��6��.�kl��lEx.K��6�wͣ?(�ʽ��Z ��,X�`��,X�`��{����9����'h8B ە7��~�H�js2b���le CR�f�ꝫEzmS��� ���-����.��7�3xC�"*(�i���@��B��V9��B�t��A��᢬��psS�/���]�g��)����_�7�3�pWc���Zl���s�f�w������V�4^m	k��_�����{h|���� I��=M��yH��G>\b �)���0��=IԂ3� ��R,�z��L��j�F��f�[^c��6?/d��<�-w�ɷ�<���:3��h����(�����bF�5�MC�-����Qb�s=��`�r�h�hT�}v�������Әu�����z�����#Ѱ0/�q5�w��R���E5q7�[N��y%
�d�=�F�ѳi��� �����䶣%Q�nv�u��@8�(e�P�zۢ�`�<�֣�v��,��x<]�3��])i�r��G$ٟ��v�=���lm�\���ñ{%���&G5��Ȏ:��*��;_e���	{�}�J�!�*��~�T��?�<�Q�s�3�EК�ԣ����C|�B��T�)��@Pco�����VC*��׫׮Lu|�QYÎCXo�k��;�/+lPt�vd����/~�nW��f~}u��KT�q�g����� Cĕd��GR�ԺC=5ao�&	Q��g껽��P�-j���E�+����ٓ�(����چh׆�05��<9Fy3�uI�s��yx_\��&����_�DHB�KQ�~y���V9��([�MӚ~���>���'�;�&*�K�4��7|���_����x�0��;� ��}vw��k#j���e�ԫ�������ߪ�?�uv%��K�*ҧ�%�.g]MC�j[�����?5���q��A�}!C�cy��d��9��"�:/t�9fe~�H�f�yb�ig$<� �:m>�_ �gƓ9�;�<���O ?�\ޖ/&I �1�ئ����`�~���i�Y;�rHZr�k��%Ks��E�����/X�`��,X�`��,X����}���#���A�˛חO=[�|��T�$�t��Й��⍋E��#o�o@�om[~����!![8��B�]z�"%����exr:3�fzN�'����QSf���At��B>,/	�spE�߼�V���w��_��!~�s?S� �QW�A��?5j��^M�s���;���`p'7X����0�#�9@�'9�z-a�߰�sf=��GY����i������Q�o�+�=�3z�ՖQ����I&zP��~�J�_6\m>ZR]J�d���Ԕq=�K��ŗ^*�7��[��F��_y�=�Qф�[�O��a��6F�K���TA�-Y��!��'��ڱ㢝D���w�SCi���q�E��)�����ZO!=�v����]���� �������$�OU5��$�ڦ�s��ѻ�R�	�S�z��a=��-_tn��b�k�ӹr�x���\�!IG�h"�i�Kt@�!�����n G��#E��w��d��:,-�ׄ�/5Ce=�� �:��rf��|��b��<�o�yϜ9�^H��ϳ���-�3�U�)i>d��B�=��Z����IAO�ه����{H�r��vR�hd��_��f����<ĸ��x�Ƽo}M4���F� �JK̗ZT�� �����1'ߐ��/���ݗ�5���5c-)�H6Q�2`�M|Ŷ����h�ݫmmI9�:: "K����DR��D�гZv:����+�K�E̎j�����fƣ�n��,o������&���4�ˋŔL&���%�,9h��Ҏ2ΰ��F�0�%I�򾸤e�i_�~���V�Z�j�����0&Y_J��^q����)�j���22)��h6'�y�x\���iFe?s�$�y�ѽ�iTdSO"����_}��{9�ݻ��k���}��f�S�9�1�T�'�~�H�X��2���d����,��t��9�D�&4�?��~�vw��J�+���>��@��&?�a�����𪪃��3My?�8/ϡK����A��.���ٖ����vd������h@:����%�Nx��iY����WÓѯ#�E�H��r=[x^li�$׽��뛓yHD�1�}�Y ��,X�`��,X�`��{���χ*Mi�&oP[�d�#OKt�E� ��+b��Ż�'o6/޸P�]!��7��`����~G\���L~���������@zZ�-4���B���S�)��5j��$ǿ����i��ɛ�c�遃��������s醼��?�r������r~�J%��r_����O=W�W�	�׃vZ��!C*���K�G���u�E=�9'��Q=��E6O�����ե(*[�G�\e9=�3R�vwA��<�~��"���?V��]�Ңh��h,--��L��WwC�%H>�ӆC��[ ^��[X�vu咴�#h�_z�9�z�}'�TGzF�);%p�I�<zVp\�`��A�]n5����Z`���_�?��	�o8)�D����?���~�_)��*f�3]^��i�?f��Ѝ�\W�mTM��������L᱇fa����΂ [�#�̡��Q����?.�3G�cƻs�ԯ����"m�B�#�o�܎A��	���Tc������˒F�>y��w�_�=������^.)�M�h׭�D�(n����D��F� i�&��}Dm_���=h��~R�����_jw-�G�Z�Q�{x:����
���&�:���/K>w�&2N�?���qo���mo ȿ�M��j�f���cG�����xh+H��ɿ��ט�<㕯ZߣQ�qH�G�~䃫Ҿ�}�"�4j���$�~��	�<��2\�S{�4���.콽A�Z�O�?��h�FӤ��ح?���q��j\�a�<�
��>.o�I���C��q�߬����7C1�""4�5����D�u�����i�>	f��F�%٧DY�` �a�q�4���8�_q���%��<3Z�%�j4jT���h�u�#�t���s"S�qJ�5��~#�L;��n�fwE���_��/p&�?��$�00��f�Y�\n&�S�|Sk �ź�J����w�����ߗ��=y��-Bn�|��{��+�>b	_XF���q�𜇱ս{C�� �n�˗�Y.�:�Nm��%<?& �Z ��Ʀ~��y�_R��ޔ�,������;2�w�20~�ُ�y�1�/S�:����d���9&
ˉ�3�=|R�������߳ȸ�����>�x}�[}���e�nO~�f�B\3��X ��,X�`��,X�`��{�|�W�B{JG�n^�6N��s�s�=�03d�_�.o�?�&o��  � �@t���y�lw��w�t�'A����/~�E��'>]�g�R��Q!!Z��j
RcbkC��vw���?�j�^yGH���&}�|S~�؉"�uU�H��J�ܿ��C����#xCl����3�R�?�i������HSzbf�j%xI�)=�4#���x�5�k���?>ͲJ�&|����LI~O�?�7��ㆳ_�D��p?^{��"}��3�7<�*D�����#�FC�Ӑ�U��rԘ�����B\���g���E:F4�p=�d�%��܅���d��F󥶠�nk����-�hl� 3_<��W�L.A�syQ�/kw�(�W�N�(J�@��΋G)�����C�l��'oPFi��^ܨ�>�=�Z�$3��b������'ƃ߆�ƭk����/��"}$5EX�g��qdU<����IDX�,���;���[!�\dj��d�x�E┐ �d��<6@��~$���_���~ZƟA-N�"~ō���q���Q������K=��H����8�k?-������5��RI1Zh�#�t80�����NHܺ-�d�~��,��Ͽ���}������?Ͻ�'&.݇������ݷ��D������gJB4����{�� �o�E�k���$�0��0��sR��@4��?+��v6��A������Q37*���|��\�j�a<"�  ��ޑ�xZG�,�|h�I$KrE���6�bj�a�D	���a5��mҨ⹫���2��O��%���)W��K,�3y~�%�*�@g��l�� !���F~P~$�����F]��֔�l��D�j��Kj�q�46d��NΏ�?�khl�VoL�q<�QL"X�ؔ��$T�:&���w~��6_&�b�&�~����芉���j�~'�~�6�|Ѳ�:���0/���5�}�|�\& �o^�o~`�Şq?��ޔ$߃6}��/�o=���q��`j�K�E�/r��<m����	��������^,�S���d��:.�n�e:���\-��._,���%�{j�'�}v��G+��2��|A���;2�ÇX���Y�:y�3x^�[@�(�o���$܁6��M��x�x���"����� J�a��.i'���{�(���%�#��@��o�0�锺dq���m��pN�7n�\�	�x���@�,X�`��,X�`���ؾ_�M�h�@t����!�:X_y�n^p�2=������֋Gl�����f����x�͋r�����EԾ��k�H��H�����}s������6Ry���O�GE�����o�/��^�"��r:v�x�^�)���P����Hg�E=��S� 6J �ͣg�?]��޺X�C|C��~�W��c5��7~�hDIc�g��Yy�^[�Jus��hp�'y���gԘY]]u���g��+X��/���k��"������oE��׊t�IM��+�������O����\֘�_j4����@�����qO�=+�A>�����"=�x4nnK{?zR��;o�8;/���Mi��O?!�ٸ��1J�)��V���$���̼��~��#�M���n�i_JXh6پI@#�b����U!�Y�iJ���J�{Bʭ�����ĨE��3�G2�gntI��j=��	��Ω}��@j�<��S�efV���
����f_�}�q"�M��C�؋%�/^��"M���Y� $f���f]��^6�Ĺ� �v{2���~�?-��@Sn���Zwޑq.�H0��egI3w��O����E��#�ì���¼_�I;>�h��>%��ʸ���<��$��>��Dɣ�م�ߥ�����e�p�}Q4@�u�;Ez�9�����/����:�쓉�:��f�yV��{�47�d���m�Y�����f�r�=OS$5Z��ی�x��-�3%��F�f;a9�(�T�R<+�yC��W����y��pI�}pI��XF����h�F̀�Z�w�#i�b�������W�N�^����lI�ѯ�ЙE���y!�w�<�&��N�������_���*�����}�s_�u����v���@�9�����WLҞ[_�xAʅ��!'g@��5��B�$Y��6A���.C����zRY`Y�0�G��?*�dD����,o�+@8&��f���eT�4�n�ҽU�;��gL���|�S},�%-��8ʼs����=��ϓ$�va�/��nI;�����f#����Z���^�gQÆ��y��j	��Q��7$?+�����|.��ˍ欔Kr�}P���Q�����y9��}���}\iT�w<��J�o�e�3*���	��
��@��~�/gPN�+�8��~>�h�ym�[����}����U�}���X�4��Z	c��F�ܳ���j/' b�"�wg��<nb���<�4�tE�"��J�#}��E������ҿ��U�8'�j��]h����GM�9�gO>)_�=�/gg���zs뺼y�]���p8�~daQ���Q����wvVƿ�w7��M���Iy�勩64�,��6��$�����䋙w�HytQ������k�3��ƅ>�E�~�ŝ1���7hb�Z�֏@�,X�`��,X�`�����/���7�x�}��F��8'���j���2^����������P��| oj/�#���F�+뗗�������Hϝ;���:,0�*����o�gē�E�S/�H���?*�k�&��qyC������T�\�'�w��*(����#�Ds��&#�8
6��{��iL��T=����ŖT1˧�غĬ�s�xx��ܦ%�%2��#�9rJ���!k:+�1�g�#Zx��?�u�-I(ܯED����{��h&,.�8����tl����S�	�p�����H[G�=���"��J��+-��u!kg੹������C(�1�Hcr�?�YϓOs�Kz w7�4�]B�=�-z���x,��t�z�T��G������8s���N$�����?�rz�</�l5�4֜��$���e�I[��~l��	�Q�,X��g(i�S�r�$ˡ�]Ҡ%��c ��O|�H�r3K \�_jtlo�罪]c͔�!H(��K׎��㋒��ۈ��q\�s��'��22dS��%}�D�zQ�#c���6gp�P=�Y�����"}��J4�G�hK���H2���|$�4���XAF�,����^�]���b��^�#����/�O)���mt�@n-��i�q��^�j~7�zV�tf���E^s������e�=%q�]e��}uۓ�Z��M�j����b�6�F�(�!zn�oCC�i_��?+҅��?{XH��e?���T����_�F�cM&],)Ũ��W���_)Ҿ��d��%��$�we|"j�,�s�����!�y ��eC��L�7�!T���>{.H�vc��M�~��*p����q'�G��t<�>O��9��A�R.$�_|Z�ӿ���$��t��e���I�ǯ���e;L���%7S�ig̫��/THR�S��nf�xQ0�2�7�M��]f(��7d���o���<_����Y����O��R�����-�Μ�3Y����[n6��)I@��&4a9Qd?��	�ss$���<�>��`��_d���85�/�fQ]�6�h߇ڋ�qI��Ĭ��V�Ӟ�q����Gl�/B��6�Ls��_=,_�e;�w��g�g��Z˧[o5(uu�.�;�A��Us�C�_�/-�PLO>�^�Y�5���7K��x�i�R�$���HZηUy��Nhǽ�/)� ɗ"6޿��we�i�t<wB���ҏ�D���7��~�����{�k��5�To���"��������H/_�X��s�g�96��z|銼O��}����k���*�'�yF�M)ד+r�]D~o]��h":6�b���1D;�x���ܒ���|����7��8�/X�`��,X�`��,X����Y�Ͼ���>��v�q[��I�{}}���CD�Z��m���,G
�`kM�I.�'�5Y>ȥݹ#��O��"=p`�9��יh�r��������O��W�����ɛ����7�Y��~��t��
�x6|O~�%o�W�1��n���s��/]���Q�<R��.jm�jhI%�ϣ�7�*�`��M�x�M�d�DO�1 �)vWs��׮��_�D�~�߈羉7�$X��/�6��K[�/���d_��> ��yi���Z1��O45ɒD\�	���wES2^�fY*s�iA=DE�# 5Z���<pH<��#�������r���J�0v獠��q[��!�;iDR��7��i����g�0�o
i�h�1
41Zich�F��0��KR�s�Tj��[^����Sg���7�_��c�)du-���[��]�*�7p+0I�Q�*�TE��U&$�6�ţ��h�z��@�9,d�ր$�w	�EJ�_��`� )+n�/�gJƙ�EbB�D7j�|�l��/#�߰$���!���%����/;�1J��S�?���A��'�y�h{��������d�y_e���������3X	A"D $DP"A9b�Y�pX!9����dXr0d+B^eR6i�A�$�3�0��`�}z�����o_�^����|�͹'뾪��g �����WU�ܼy����������3Nk 4��e�%�רI9GC����Y�T��p����o$5�6ڒ��������D����Z���C�s �تC�9H׽Z�(�'{����}����xg���D�A�%Qx�j85�4�����b1	R �Y���gw�B���S@=�Γ�����h$�Ve>��A��r$�GR�ѺY.���
F9�1��̫�I�0��(���na�x[1V���ز���a��dgd��l¼�Ю�DW���GE�Ƒ���4Q��ϰDۖ㐭aN��i���4�D��Mg���ءy!��|��	���ttcJE�����D������:��mP�֝��&�� �X/����WV2@ޮ�
�]A��Q���V/W�6�8�Q����Z�E��y�����ݓ�JΫ���O3�lȕ
���ay�#��B�z��8���;N+��y�1'����F���Q�5�Ͻ(�N4�����v�u�a�V�����kD���}���9s���Ͱ�ԸfJ�1N�V�h��(D�G���ݟ��}���&����,�H}�+fx�Gr�=�wuEH�7����cE%�u$_q �bᰬ$9{B�W�-�iP���j������Dz*N�~�q����������XIt�3q� ��x]��M�|���ه�Gݶҙ���Gf���ې����0.@���i���=�;X1�(�������*���}޼y��͛7o޼y��͛7o޼}l�}�=t�>�Q�ȥȳ���mcM�ʺh�ժ����6�+;^�$oN�]�/��7���`�7��[qʵ�t��|Z3�&�N3�M�=�t���٣�V��yӼ�hUK+R+kBR�兞���G�=~@�f�.��R��˵��	���?�QK�h!8<��ʕh8kn$=ˊ�ٯf��l�=ьZ�hd�ј��i���B�����q��3�7�����ߎ�_������Ю_�c�@j�ٮyj1a	���m�v�Wωf�b�{����2��֪��.�3�	��4斯�������t���E�����(R�n���#b���v�cپ�_>Ϩd��d=�K�B���$Q	��r�g^��HO~�4�z��u�>>oBs���'oOٻ���D�e�F�8W�3�MH�����0ɘ�D�	i(�y�:��7�d��_�C2R����|�b���h�<�C����eژ������9/��2�+��-���h��#73��l�ǡ�ם��+�+PekS�O�$�ѽ�nH��W���_H�_@=���:���޿��8�Ɨ�l�-H�����K����`h��!�F���}�[qJ���B	�
)�R)#����<Κ�J������h�����=,G���U��홱=14��˯"FO��x�q<��gM>q�|"����AF�NGOU7��7��=u2N��ov������}"N�����i�"�3*4k	�D��L<d;5_2ڨ��`n�;B:]�v'����Q�L��5�]T��/��Gr���B�*�(͝�g��v��WBG�33�aw=~��#{{CD��$�n��t�U�Ql�\�H]o�iv�<eDM劅
�&흨(>S��MC��?4�X��G������L�����a�=��$5y� � ��Kpx��o(�F��ΆlS���Ѿ�	��c�6���A>��|�M���9��u�v�b�ⳋ�ޭ��o^�
�S2��#?<�o����`���P�~asc�u?O��I����B��B����#sS��n����y.�+��5�'��v0���N�N�l�9>�"s���ݻ����߳�曲��
2�l��ڇ��]]w{(�E�e�-�dQ�A�� "{���{��h��K�^�"����^+
��ߧL�ӏJ��3�����N��S��i��}���墐z׮�{$Ӯ��j	�OH�F�|��9�#Mee\���gkM��!���|/�q/G-p��O���������d���f*8��K��/�-<��͛7o޼y��͛7o޼y����G����/T)mQ��3����q�p��,�n�qַ�*dœ�˙�����s������%��]��{�C>2V>�k�o��_��7ؑ��>=�]����4Ney��o���|�o��<�V�C�h�ؤ ?v@��>sY�՘7.h�u}���z��&��h���h i�(��E�N���)h/�x�_�=A�g�v2b�vIF�|F��>.�
��i�,K�ɏF$�͠�E�,>,�_������?�/D��Ձx\~�O�8N�����B�.LA��! �*(�2<.��xf"h�����'q�RO��I�B+��T��<��R�>�Y�<m�{-�������n�q�l�1]�r��#V�i��$�㮻�������"��v�(�&j(��5�s�x��ſ�_p�hd��1D�Hzd*u��0�=�Yxv���똞���e!�
��3�}J��h�9H�T�9���ʗh9����Q�� ��d|8�x1N�������y_�z@��~��qzyU�ɻ���̣���q�!��*H���e�*6c�gŲK�h6��:d�sn"�#������.�ēm{���	R�?�z[-xq��]����D�/������}����3��/6��x��[q��/��G�į|����3x�r�pa�Q��Bx��s?�ӗ��7WOk�����Y��|�+���m���.��0�Y}��(�np���C�E-B�gFk46�h�͚�_y� �،D8��NH��SZ�f\��_�Ճ1Z�k��h��_�n!���A�T[�&�5\�Hƿ?xB�c�xH����3��D";�j0�S ��C>�k�6��������������B��}+�J�����8��8/��1���&/���}S��Vp\7�쏇�ӱ}Q[���{3~��Q�V������d�E��_S�2߼�&���7ì�� Rd��+5�H<S-U7s�,p���e�緈�ۜ��� 4�,�<�¹��/��oo�p|��]��|����d��������"��� I?���*��	Uh�1�J�OpEZ��d�x�m��Kk`E������/�|��}�;q��;���!�<+�+AcMM�F���ȟn�k�����_�vr�C��ZC�=�Y�ũI�[V��hQ8��6�:�Ôf�>��Fo��/nm�Ok����b�k�e<:���j�Y����c����+2_��"����Tѯ��v����i.u��\�r�^A ��Ђ�����_�g������O9�W�_V���k��Cv$?S�e�J��"�V6��*�Nr�V\�`E�fW�/[�<�����?r� ���� ��� 6E�T��1�<��͛7o޼y��͛7o޼y����G�&�� ��&x�/��E����8�h�>M�п���}+�r<C�����.ʛ�BQ<pö��w~GȐX+��g}�r7/6Ӥ�tE�$�s��,/��aQ�~ͯ_���(����� �4�#S-H�m�q�W����-H1�b�F?��A{K��ʓO�� E�>�|�q����5�\��}^F�TZB�����s���;������:Ϟ�|�O--�}�r��m��+�a�Z�z��~�� ��(��{��x�mH�N���ʦx�庅�J!4
2E�0�҉��t��B�:$��7^����n�] �9_	�,%h��ղR�5�8�����Ӣ)�(��}!�迆C!��Ƙф�w�*��om�3`�lS��%=� �ڈzJ�'֧phGA,�8�A�fk]���Zg}�rWΪ�&QIC��}\h}!�qљ�jW����|�����jK��1-���A!����99�����x�/�s13��#�UpRK�$(�nWE?צH��p��T*Ԥ����,�cw b��F�ڌ'ؼ^yI��z(N?������gX��z�~��%Q��S<�u�;�"ZA~H�tA~D�BZ���qPȽ�P��,�(���zD"�2U���-�?s3r��|KH���~��Ϣ�63�HMH"'��G�/AbL�냨:��qJh����
,J�e?��)?9~����뒯k�Ɯ?&����'�R㸂�(rQk�e�D.�/�52;�ɫ��&�Yg��l�*�>��_�WIPo�L�9,��
Ⱦ��w�e���ޒ�B���p����� _��b�~���\*KJ�y}CȯW��<���C���&<U����A��$��ry�%h��Hҙ��ʟ���4���hA���WdÄ��~��h����y�p`oWqU�����CV>����C2��<V*�/
���hi3�85$oH��rM~p_jْ8�����i�s�$����h���R��м���_�SF�5��=-D�x�iC$]҉��%>w@�wF�L���Q{^e~���
�_y�� ����[���C=_�%��.6�H����wI���g^�r��hs~+��f���R�7�~�)gW���{Oȭ���<�xn ��@���q�פֿ�R@�މ�]F}?�~��79��'{�<1�3��j��RL?����k�~8�%���ҏ�cE�j{M���H��d^7�}nBKz�,��X9��DRy�7h���)R�W�k���o�W�Z{�ǿ�߰H^}�)�?�k6e97u۳�c���M�Շ�+�fd����wXaW��w���g<��Q�:ؾ���K�/]ޮ��D�7o޼y��͛7o޼y��͛7o�e}$��,d�ciH�1����u�	k��3:�64��]퀍M�����?�'�u���ӎ���ӖҺ0��7�����<v<N_8'�Ƭ�,/�'����yxh����K�+x�~Zjo]?'���Et3�7c�>�����MvQ�ju)�����
���a��S�F�W������r�^�,�����`E(�j�l�0� �"�d���r��E��zr�[���"j_Z���Lb���.]��4� zJY�g����� ��-.Qx$�N[�_�OP�G-����B��=n��PKÚ�d�H'j�q��>�7$�k6G�����ۓe�ӓ�<|B<7}\'��Q���4C��L��M���?��h�(�rU<Ŭ�kЂd�h��x�BSѬ�Mm�F�4j�У��6����W�'�7gD��y���XH�%=gr�*<���I=�C�f�����(7Z��<�èů>��Q5��kZ�p�f4����~?3�\`%�S�G��U!�%Ŵ�~�ў��c�v4�f�y�e!	|@Ⱦ�-��C�o�K"S�?����j����N�z�~ �&I?+���m�W��P�K?�/�������,I@c��$����ץ@���T�F����qı"�>��Sq��(�$��~T�ũ��cn4go��E��a��\z�Y!9Ki?7.��RG?e���ۅ��P�N&���4d?�����ikA'd�9����Mv��z���(Ҹ�<�k�r��(�Qƕ+����6*�������G�9_�3�"�xB���XD;_���A�9�yڳ�63���B���Y�����|.�a��J�/�#7kc��a�Ac���D���m�gZ�$����ٟ�|�n�K���3�����hf��x�a���� �y�x;��#X�D�������}���}y�g��ձ���3j �����Z��e���������8��ߍ�V�8� �{�q|�g���T��6)�Oc
D���$�q�jf���Nj�_D�
G�4����A~sr�������D��f��I��9<��d4�Q׶��|�{|m����������2���K�Q�P�ж0c}I��;a}�,�����4A��[����fj��� p���w����x5_Ŋ���4�;2�=�[~뼼�la^�fi3'���g�y�Q�����C3' ������_��˗��~���㴀dw�uG��蠯.�
�i��+pr��Uǀu��@ƙ�{��K�����IP����?|�r�౱�v�ݓqi����Pqw�D�7o޼y��͛7o޼y��͛7o��E�̯C;�*H�uD%����C�~9ǫ|$l�`��ہVV�7��x..^x�<�ȣqz�m�#�+��	>�8�m�G�^�����M�%T}h�e��O`�yhk��͑����X�!�L�6��.H�3=�q1�N��\�QM��M�o_��/�igK�p����4|�5���C���G�ל��ojr̓8��vw�<"���-hZ":�&�E�j��	�O�ܰ#w��F�$�����5+_,?�]u�R�Na�JS<9�,<h��)�px�E!���1Dš�`bF�t5��9KG7ݝ�ay��D����q�gn�-N_}A/��+F�3�C�f��<$��������?���cC-BF�#iІMk�P#�$"5&�j��`j�������~{��t�|�9��l��!���?.��t��.P$*z)��ǥ'�d�
�Z���h�kkR�� ���ّ�[����|߅֤�RIR1��PKQ]Z�pwf��3�Jtlo�k�{��E���/���x�Ah@3*W���ΰ���4G����d��Fꃟ|,N[ [֯�v�P���]�C����ЮH䵇�Fc�E|���z�q�@z��ȫlׅ�: �� ��v��ڦL� 2ȿ��	���h�v`4]���3� �4��w��?�\��9��FW#~8����{>!d���qz�>����Eh?�P�̑�@#��w�o�O��v�j|�O�r?q���1�a�����%~��8\���>�m�ۚ��6��e,�!��Ά��%��S�8o0ZA�ߵ���V�"�y]�~Z�3fq���4W��ݿ7��O)rm�Qҿ$$�=`�J+�Z���r�%�	��_$>�!ɶ�����ߋ�<��ڴ���\������!��'��ο.Ws����ɶ�_����$�W	���ۄ�G��H��`e����|�+�EhyB�j��ko��&�K8n��+#����%	��4�5P�^�)�ʁ��q��h�)b�����褚�4�OyQx]�=I\��\�qkU��K��{��b��ro�yc�`t�v���R�����|�� D�?�m'�C+��H������/C��G����OG��w��q���J�oo%�����	�O+���7�]&oP��҅8-��,[�~�T���~��%1�W��od���|��Ͽ���0N_�
����]����?M�4��,�Ň��{Qx�$�pt����d�9<+����e�盼�v�x���B�L��x_��J�R�I�e��*]O�y��͛7o޼y��͛7o޼y����_����5�K}��o��32�����e+�F���Yx�W������P�6���H�
Ry���_�%�x�%��j&s��j0��{E�P������6>j��m�$��{W�������p�,��1�W�=!�@���h}����}��'�X(ʛ�:�}1�l-�y�B���\�&H�t�4�R$�����v�C�@��I�"�G��XX�6��]o64�a<��r�7�$x��������"�3]2�����'a>#�=�W�a@�]�mD�}�u!�ʈrJ"��}á�i�-큐��}j�2�mt=K�����V�gD$��Bc�����`(��,�=ȑ��Em=j��{A�O����p�
�i���kmEH�Y�Dca�+(�`tO:ښ�3�b���j�Г�G>x]uDA%i8dTU���0����4��M�x]�*�2|a��w�]U��؎�Y6Z�(j�ՠ-Bk ��߳���-Jt�C���F��w�-ǫ�3 �C���ƥ.�p�v`����	����r�Q[�v:]lg$&�h0fRU�y@M<h=&����>-_���Ӳ]	�z�I�����S��h�� �授�x0����C��vgQ}�Cl�ݚ5���cr{�5��������)����\O����3��\1�d�cfg�}W?������u;\�ߩњ�����Qj�3٢vY��Ï=��<(�mC`�k�N�A�>��V�<�R�����(σ��Ζ�>o^�-��L}��ѱ5g�!����ett���7H���M<ik��wT'��i!�:?� Ӗ���������_G��a0�	�dk=S��Aj�Oa�*	s�@�ݮ��3���GWh�71E�s���.��j�|���,���ޖ��ܔ�^�677���������G�F�$E�}���sܞ�|�\�r1� �a��ݵ��ln��2�CM:M�%���i�pT���	m;����\� �4��s�ү]{O�G�f��m*��<�G�P�V���\�C��Z�$R�GB��A��gd��C4�c'd����o�'aO�,/�ڍ�/&%�6Q��o�cG�n���=�4xZٵj��g��V��>���PK���YƼs�D���Ϝg�vٱ�L�7���X0�v����F��%^�	!<�>�@P������������3��d5绸�YL�X�G��I�cpV��#�!�?g0��E�u+ {e���K\o�>`S�k��S�~���^������8]�!��"�G��O��<? (u/�Z���;���/^�q�W1S�F�6�3�����q�>o޼y��͛7o޼y��͛7o�>��}�� �Sj��3�U@���a�#��6�"j#!���ޤ��Ah� �����9�iU�>��̻H��Q���H�l�3i<���óF?*I>��H��>jm��BS�AG?��>��D*��@����P���V��zT���W�M|4��_}O�IzT�z/WL���)5�� �HHD��G�A(3�2S���^[[�~g�i�t��A���k�"��(���rL��P�z(�Rju�R�	�14Ѯ�=x�I��и8"��6�Ё< �EjR��ݑcB�D[��\��';
`Zp$ۊ ����W7�@}&ag$Q��XcF؟���T��ZE��,��A��y�.]����$��ޡ&"�rW�����v��ں���)i���ܷ"�K\bv������~9t��4Op��曹G��?��8�HB�r�˫��d�ڀ�'��;�+NIZ�(�b��!a`kQN͉��R����\:A�g�c;�ү��Rv�l�r|CVhr�Q^S%2�C�v���!OA�� ⸱dZXEh�1t9��t#�z����VԮچ��ֆ��� |t��(կ�&	�@��Ѥ�4NCFYEN��j%�8�/��mu����L-�1ͬb25VQjR�4�h�8���&�S��t���'���Y{{���Kv��y�}��D����'Q8�N����vf���9��I�?hx�<C��i�`\I��GB�ǝ�K��mfV�+jR���E�C�6��| ��D�g�/%jj+ J��{XAAR��dά@A���bYC��c6?٣��nm�}{E
���u������z�%hC�=0::��y��$-溱"�)a�^\mX4f�N��#t޷P��,��N�=�|rE����""i��q�3G�/T�[[	Z�f��G�<E�H4Rc�
��k��6e�UG�5іQ��hw�#:
����q��^W?�;�)��.u����]��Z��	&;��+���]��w���V��dPRv[�JD�{`Z��"����Q�����m`%�t��ڏ��Ӧ�9¼�ӟ��8���忈��mĞX��ߓ�D�98����o$<�"@,��J8_�Ն�۸_!��fe�;$ñ҂��0�������͛7o޼y��͛7o޼y���#`c_�i (�5�Ԓ�G�ۥ����9֮#݆�� �� �Tސn³L2瞻%���:�5�7�1�Q�ٳᩡ�ZH����ˇq�M�3M�%V��c�9��G�u׼��sa�����<�F��&�&](���)�����}�7���u�=�Lj0%O�eH��d�N�O��K�g)��o��b��3��Ky�KS��(¸����5d\GBQ>��KO5�h/����K�J	��"ȴ��@�6�ք������0�D1��-mR���Լ���/�'%%K4y �� I�u:6bHY��3�]m1��c;�"z)50X΅��Q#L��&��1��ӌ����]؇縇�^`?�ǡF��<xWW�4���m�r;jY�vS����������f����h��'��H���K����U��L:z�y��{hZ�
�ez����j��JU��m�8$���u��I���D��8o�G��n?�{��Y�[� �k��4���6����o�,ˤ�%{C5����N�CS��#�Ki$�������k��>36�p�xF�e��A��lL��q6���8��Vэ�+���#)�Ǳ4��If�z�vmz��?�y%���S�uF��ړ$R{=[S���U�k�Y/\8�$�R^�+�d�<�F�̜6Zs7@91�y� ��&�&�>E�1�mv�
Ab��,�Vy�$�-�.>�%��b{����8/ʁ,L��r\g��<H��Y!+ז��/�@�����8��<�bU��5�~S[��M�|��u2�F�� � `�D$!���V�8�2m�����<�Ѷ��#˙�DI=�>'�c���I�a�W&�ٍ�}?�:��󕳼n�R�3�O`}N?�r����̟ԍ��u���t�����y�H)d���WV��c���g����ڼq���I�M��}6N���?��MD���D
-`jIs��z銨�?�����r\�$����e���o��=�xS2�}'�Jo޼y��͛7o޼y��͛7o޼����_����ԚҚO�\����2�Ȯ6<���繖��ҒhiA><��'p<�\�'}��j��T5)�!o�4y������� ��`��H>�~ڱ��zZrYz�l�/"�PCHࠣ�y�Nt0ڣ�EW ED��j�\�&$_{ ��Py~LTbS���~�.�>�㥋�Qv�58�����eԍ���Cƃ��]��@��ZV���w��8=�Ԣ����N!D�SaӨ7���I�ˍ��>�/zj�1��-z�QԤԄ���T{l=������wB�(���v�&{��Y�$��ÕQ�𻉺�Ð `y�8y<NI���!y��~ L� �[ :I���+�mͿÇE����mmW0C4�(o.c���"�<�M��)�-��}ޝ�sqs��X�J c7�I(���!�O2�D�d8D%&�pd�o\~Hf��֬��XVE˻~M���[���cs��n6�LFo�5��W��hm���He�@���7�6�܇�Z��V�.�\��5r���q��F�{,�2����a���҇3��t��{6�^��7ӄHd��S����q5:�qB���W^�ә"������q����p��ǳ�&Y�~�9a6S��Il���e̗9��On+�i����ϱ����r|h��p^��l��u�vQ�oHtr����&�Y��l4(I\q�A�	��g����mH��RN�"�J)��h�b<�~,w��`�[��$&I��9��_oH� ���o�isN���H}�H�H�������r^��~�����f�`$!�D��x�9���Q��X3��t��T�F~8���++4i���/&|�s/�K4���y�8$�JH��e�e��3�Z?G�qs셪����^I�(�������<w���!5�J�ɍ�����»-F�'��������� �'-��������>+Z}���o��ڪ�w�-�
���n�S���i��UM���zA��TM����(��bI�c5V�V^����͛7o޼y��͛7o޼y���#`{~�G2��GF��+-�`Ğ����?�2��
p�W������
�v��I�� q�{�C�'ި�TE���5z��Ӟ��{�}:^nV,g�l+Hή@)��|�PNW�3ۇn'[;�!�e��g��Ef�@L��F�)Sh�r;j����U��i���C�ҙ�	�q�m��b�P]��mo�p|h]�~� �jcF�#qI�P�=׌��B4��Ǭ*���Z��OR3����JF��6�XA�o6$����:�W6��^6g��lvr��(3Q�P�&z^ ���& �7���q��#�ik��O�������'�5�O�MhX�CL2��q�Q�Ip�$2��AEF�r0D֡qC����Mtt%�d��n(m#�� �f H���6R�WGOA��<���(\���3�6��j �h@��1��	S��*ux��5��蛣�$M�m'*�xN@Q����Qn?��^�$/��u �>ۯ����j"�ڀ=x�I:�q-Aǝa�6�`�n#j��6�$�(���{�����}�z��<4����gCF'���4aMMP{�)-m����b�v5�e�oI=��n��$�I�I�&[m@#������oׯ�J�̃�05ޫr�8v���Ο���8Er=$�j���x@����+�cjJ�ūWq<�Ǟ����9�B4����d;*�NYEn�]'�xү��`]���y�}��F��+tR����w�t��h�q��zT(QW��/�?�!\����q�1�/���b�:PF��c'�Y����TS�g�,��nc\P�i�I�a\�����y$5���]+)�-5�����mJ{O�С�IOs�=?�����>!@e���^��%���j�c��Ol��A�7]^Z�s�'��LI\g暢ZEo����p~����}���C�}
��[���ٸ3�||�$��1������������E�f�X�qjmUƯm}S3���σ9�_� �h��sZ�~�a�g|����f��{%�=��͛7o޼y��͛7o޼y����G������h���x3�g���x�2��`�3�8��=����֙�@�;{�:{��G�d�l�@���)�;m�ŝ˓�m��vJ���yoh�xf؞Pf�������%	d��[��D����%��=�.��O���)O}�w���d����2ګ�L!�@O��c��2�R1�qir
Q���}��ƺD��p\�'�<���ƞ���+ ��W���k�L��rc	�C2$�>z�o��I��$��������r��h��.^��о�OG��,���.�E�?�+I�&���ɴ�h�Ez]���>4q@�V�('��2� �JSn�~LoG�C[�e�u����˚�$׵t]��>��/��Az��h-^������P��|�P�~�Ў�K�!!�@�(�t�^VwE8�~�ՐT������+�!�&��v���:�׌=�f@�.ѹ[f���|���\;�C�m�$�k���w�R&2���>؟��g������i�T5D[E?�G��%h]�xO���+��ܶ/ �%!�e�چv�LI���B`fП2��Hl�|��j%��K���^Ծd�|q>Q���|d74���~DKr�fwl:�#G�(#��~�Ѫ�7�$���$\�kk���ܤ�Uyge�lF��0�g��{֫��m�&��ls]�\��D�-p\��I,��$�D0!�@�!-B#�XA;�����H���I!�*�~��N_��&j�ꨩ���5��-���Ÿq��s).���	��4���<躮��!�7l��m��W�8��<#�����筛���{�[s:}5� �f_r�e��AM���p^=T+��hW�2����'��c:?��/��K��tg$0H>�O����f%��J�U�s�pG��/�++Á�2�f�����p�'��y��͛7o޼y��͛7o޼y��މ�5$lM�<S��`�~��x7۫7���D��q�MoR��O�i�=h�N��<��8�/�<)CK:h�U�${�*3��-د��"�3`4��� �0��vwE�(v�R@�VOu�P`��O�)6�.�C���<��Sͨ\:��:�K���:��6U��RI<a�+BP��"	�	�5�b�W���}��D�~k��L�g�>�L��h�f]I)ot��ct��Al/���ƚ�?����`;C6�v��J�G��˱��^J��G;��}d�W.^��gO�)�#�脈^L�DR�����%Qje7�#]x��#���ڤGEyRbhw�tFk�-.Jt���K��vo�*ڋ��%_O�ٷ���ѓ8��[������E4?��PฯFDwk��c��Oi���8��4٧����e��h���Dc�w��?fsk�f&����c��G)�7�F�i�)���pb����y����\7�+5�Bk�%+2l2p�|[BjM�J��LQ��vTt��ԙ��OH��5!�ُw��70ѝ˙�L�����	�j�����$��y[ltuEA>�D�_�yn,��Y�ǿK.Y�cy�F#Z{c:�6��P�����	���2>O0?$>I�W����F�d�?�z�����7�"�+f؜j ��B+8�D�?��<^�$�+�h��la����[���%��8�3d�I;�0�'�ѳj@tk0�g�7��N�s���7Z����A��6WtXLy�<8OMJ��~h�7В��G�H�5)�M�AӔXs*���h�v������f�f��K��ၙ9ل���'���w���E,�T�vOұ����w�%��.����0O?9��M�,3�r�'����y�����D5o3��$�>o޼y��͛7o޼y��͛7o�>��}$��NѺB�u���tRo���Hx3Z�5�̛Y���<�5sk�����6H"�S���]�C�7������)�j��ljt�o㈉��#[l�OS�GG�I�C���+����m��M\���>��Vkr�T]GBʐ����d��6�)�>[�0J������:�C��LS��3'$��o���/J��jS<0W�
y��E�h���i�)���0���L�W�@�n�r��Á�q��qmQ4��y흑��tjF���|Q������K���i{�����	��0�����������겐��̹����Z�{�z�� %��h���x$�X^�Ib�OA�1c$���Lr�\��&F�'��q+���ߠ��+/<�Gn?��}�8=��h��#���h��5|=z(�u�t�k�/ӏ�H���G��B��7�:)-6��������2����N�/;��������&���=�`�Q���兯���I�����%�"H��9C#7�i��a{�G͖�h�v�F\G���%!��J���3�߹�؎�wvT�K�
�6wT�k++q�B��h��	��1�e��	FE!�g���&�H���N �_")��(���#(�E?K�+H��?_�v��V"Q�,�Ȧ_`��j�9\�k4�X��s
�t"L�/���Z�$iC�R�d#�7P���Gy�Ԛ���a9p��_ϑz�F�5�+��ɿ	��h��B���y���%���F�.�~/�>'�9�/�Q�N�6|5�uL�]���C���^;�d>����ǌ��Gǎ�Ϩ�4�朱���]W�:�.8U���~r�/���z������v%$-��S��~'�=�}�6����C����?�ī�j��:6���Puh�VK�B����.�-+Ǯd���F=k��
m�h&3�y�ϛ7o޼y��͛7o޼y��͛�����E��y!^� _a����c�'��s!Q�1��=Y�}��}�`R��}�����:,�1�3*=�ExO���)}B}�N3���&-�T4>z�l̀q:)2�����ztt&]��(�vT��ua���eԮ���D��h�����ҤHy���#�*3��ˎ?۞���W�oƱ��)�Ey�5�e���{��2A�lXEt�)D�夃:s�L�^� �k��;O��g���8���涷����Щӧ�t������G���}S8�xl�Eh�@����|�������4��<�xJ���΢���3��2���)'��f5��;3$A=���hŉ�}�@}Aͦ�
/�(��A�<"��FS<_s� !�@�$�������C�B�*By@[�J�����ȍ��N�t�"?��ΉvS!���C����ٷ�-��	h^�����i��D4��E��${xCt?�򭴻�跃5U���q'ݩ&�𭉎ʎ� =��9-Nl��F�P����'�W�W�(Ͱ_@���$����'Ǳ��$������N&:Ck?g4�}�	���/]�!��r	3�3���dC4�w�v����Ǡ4��{�B2�ul��_�\�� ��g�M�*E��q��1-DWư�0����f��q@:9$DT{�g��@��(���b�v0�D/��ׄ��wh>�z��>��9��v=渵�"�sZs渨�պ�Ԡ+�m���e�@r��!�WA,�?&q�ҏ^�� �I�s��L��B�!I����if)RO�ha��d����8�e��9^� ׳��j�)W0���>d��o��#)����N[��ԣZM���a�w����2��������>S3��nVe|�`E��r�;����\�u�&��GJ�0ʦ�k=��4)����ޟ�w&�l�������x�s|6ڻ�Լ�H�i�w��y��>����ߓ��4Ao~����1�Ik��!�"u?��U�#f��� >:�;���`׏�Dr���6�e?#�5<��������J���Y)��O���yc'��V�_ml�9���oj�����D�7o޼y��͛7o޼y��͛7o��E�����Uю�;2 �2��>�+�N�7����Yx̪DG"���¤G���R�& ������ۧ��1TQ�	�����r������VG��Y���Ʉ*z�I��`1D��}h���Sbk?���QW�ӎ��>I�Q���o��*⅟U**)bmϞ���xv��&e^�4�8���HĤ�Wf�M���g��5�ӽ���\���IPC��vu?�������/^�Ӈ�r�VE>��C-=h���v�q�i�ӌz�~���I��%��L!_���v��'��a?���|��P��#�(�ӝ�m\�#�7^\}F��'���O� �Y�����mn�MB1���c��f^{K��%��D��!Z15����+B>����e�%F�D�JE��ƚ�|�j�� 4(�N��3ZK�H�h5Vq�����m�*$�����h;�q��q��!I�r�'��E�	T�u��/�������|�#Pa�P�kY]AAA���ڎ���H?�-E������h$�X?X>�F�]��ա'��&ņC��0ڮ���\cu���t��-�\�ur{��&�U��8��~�]�o��%Q�ٿ��蓆�&���c~T��_�2[,��R�]��'��(�;X	S��?��&�y���M4��n��\���f&�mh����U��W�D[��q��R��T%��ÇG^o�u�J#�Q��5!�w�����8�q�H�o�ߩTd��I3�%�͆�����5�?5瘏7^}-No@S�1-��=1}9�B���j?�^Ѯi���lֹ���ݎ�c]��H���Zy�i!Z8�0���|���>=+�_�RkP�j���ER�W{���b�@���|���s倌�Y�J�RN���ӷ��ҢK�[�����,Ʊ,�A���M���ҽ�&�]�s��/�W>O�1f��}�@�Ct�9���8�d����8>��S'V߻Hn���0\y��=�`-�y�s���ݬ��f-HX�����!����\a�眎|��(�7]��̾>/�y��z	��Ɔ��`e��8�X�]̻��dkI�?�x����X��r�,�d���(�da�|x�ϛ7o޼y��͛7o޼y��͛���M��O��*�L��D�k[���xe���x��{���R�$��Ejc@#�1-���h��R�۞�I�cߒ �%x����aq�w�i0�cC�bD�
ւ�5�� P�K�}ӧM2R��U���}6y�7�Z.�4��ݾ���M�oCt�� ��E�z4�6��g�����.Bǔ�}%���<�z�zvT M��@�����R�o{s��|�*Ĕ�lQ��yd���3j/+<I��y�zC<*�HԯZS<7�H� 1���: �H�rv�ݒ�L�~����oo��]y�^zĻ "��<���v	�<����=�0׀����h���l	)�K���#�k��|�����V��_jA���>�jFK*��#/����U��Va$t�$���N���I�=����FI!G����4āMjO�w�/���-�'Q���O��$*�!?�����5�p��$Dk����G�F���l�7�e�����l�,����LEu児�%i���e*ʙ9�M�z�^Q_��eG�+U�В���8ph j�/�@r�� ��ě�pdnC�i"H�_zS'�8j���"�3v}ea������c�'v%v9Nl����N�\$C[��j�>x�.��Ԓ�ٟ��7�� �6�ڪh��p�Fs�̿rVj$���J��6��z��cl��Y���������Zmͦd����'9��1Z.���)<�4��v�].hfFH��h�v����n�.�䛚a8D<݀&���?F3o��������q�����8��|ۛ�����5eܟ��q���sY�	�;އ)��Dswυ���s�'ǿz�:�#��T�Y�r��e^��3*0�'$�9�����h�����/'�x����ʊ��;=!��Q�z24��~Ł��nR�3�����U�C��ȑ��5�n�=7k>;���5�M�8��|��>`��6>�,�������b;�ϩ�1� ����!ow��5�A�؟��Yh�+�o[�i���ww����I��^���uy��a�j+�zx����g�I���K7���׹R��y�^Q�{R�GF��'��y��͛7o޼y��͛7o޼y�؞_��h^G��������f���G�7����O����]x�"Zӛ��F����gј�v�x����8���� ��P����� j#L�?�1��ZN�ìI�d?1jp$�Y�OZ��zJ�ɕ�1�*��$��XJ�"���������K4�p:��8uR.	j�����B�<2�h4��!�#xJ��im�T%��5;@K-cTFj����P�H�g�X=h�QK��矏�;�'N�H�<ȱb�Zr��:�,Զ`Կ*4�x�$�:�R�4 !i��4��˨���Q#0kP.9NȖn�$�>SC-q��o`�}�#���1dHjevf����9�����<H�0�_�M�Q�#��}$������Dj���՚܏BN��ehP�s �*BPԡ;;+DK�Di�:�1x�Ԙ�3�f;��6O��v����s��!���/�*���a?�ɰ$j,�a����H���$q��r��r<�q��+2�|��1N��&��}�����~��ɷ����okB<!�T��03��'��$�0ci)"x�C{\2d�S'Nm��(T2�l�p�Yv��8>�p{�>�%Z|��9�$!LG]Nr�"]\��.I7?��M���n4�FϏR�@�H2�D���^q�q��k��<��z�ڰ��75-���#�zC���#���i���T�W�/��φp��hZ�C�l��9=���Z�S���_��Hʸ�Ӗ��4��yCH�^G�/j��v��´f���$_��������'�kE�Sk7RߧL5ptu�߮-���+5)'��S��2�����T���1��~�?'QWI��@�w0�;!���/��-jG�?������ӫ�oH~0�Ct��7����D��ؐ������5_�|�1��8�f���i��~�t�h�FC�����$X�V<D��;�� �f�0��1:�^]�1i�	�t>]���6��Z�9N�����v�� �"�8��blw�ybe[չ��?���T�G���w9n+��<�E?�uE��]�>j��vcSʑѥ������q��r'-R�F��K��i��U���=�}��hLs��z��uo޼y��͛7o޼y��͛7o޼����/��'����Rs/"�6ױ}n�����E����Q��t%NW�D#�ȂD�*a������&<�C,�|�� ����
|R��V[�0on�'�G>�5zX�%���º�$��M���Ӊ�ڳn{f�c� T������6>:=�+��s�愾	㑲&RQvI���M��i~W$5]�K����0$�'m�=QUD��X��LҎ�;�r�pt4W�!���mmG~(���x䷖o�($�(��ҁ]�<�����x��7���2�9����NW�A	k��v��;�����ڂ$��'5`y0ʫ�+�C֘AVFT:D�cT�!�b���!E���mU���cq��"Z@��\����8����H�P,Ѳ��XB����"�Ԩ�}EFZ��@Ƒ�c�@;$���5D�r�G*�Ǟ�sh��d�P�Wf%e}����6P��rU��9��B�Ȋ�D]>r�h��Fm=�{N�f��O��a�f�h�f��bF�:��qz`A�ɓ�컶x�:{	�V��G$y�*���f�y�#�q�yP��@KwVȉ�eh8���Ư��8��VRG�����$8��_x&N� 0표���v�q،�M�@��dP�h��Y�W�(���}B������>(�>����sRKie��Z�&�DY��]laa�7���V�D	�Q��4�>XK����yMH�n@b����-j�;H>�	�'���<3'�-!fH;>~F���W����>@��_�a��R	�m^��W��6U��Z��M�����~NH�&ji��] i�����ۃv.�ȷBV�K�N�\�&��A���9k�c��"��וF_d�'��m�e����3���ޔq����,���Ŀ��Zs����NK���{�r=���2nS����BB0�KR,�9Rʑ�wBl��yh=��z|:N_xV������n;{vD��Ի�^z]�!�Қ��Y�>+�3p>��A㷫���"�ۍ����J�<�pH�d�p�A9��U�?�!��zKV�t��d��+�i�"����`;.�}�G�Io��W��s���y|<��%I.I���E�0>�y55��Zv�]^��}��� Z���&����?L�}B��m�^]۔�/G�2/�T)�qW���� �/��J��7�2����^�D�ѷޖ���k�bd�:4�1���=��Bk�H��4O�y��͛7o޼y��͛7o޼y���=G��g�3��B�L���H��\�ǧZ�7��F�Ƒk���;o��������v罢M���%���<`�O��L�s?,�O�o���IL���Kqz����	�ӷm��h��BDy٣F��Xqi�I��#��o��&�x����03�\��4�~��v!�1�8C�a���G�%�7�� �F��´W"B���{��"~.�M�m]�7�"F��@�l��0�+B6K�=��Y�l�)�-F��#�-Xi�������!��	��G-��mrK��Њy�igGNdA�~J�XToS�$�@�F$�@hT��^D-=�$:T{��:�����7��̩���MR�?� jd�����g>�8}�A!�3�Ī}vQ�Ͻ)�SO<�W�)W(HΊ�`3��C�p�(Ĉ.X��A�0��	�X)����xQS��!��O4�N���Ҁ�������7�3�M)�Hm�l6G'%��4��6�D�uy���8]�.D,ɛ�
ӎlm-�ED���Q���Z�v	��n�}7�$��W9N��ˣ�jz�Fv1���{q~���=o�}=h(�<-1\Fh�O]�-��O�x� B}I�N��jm�S:����(��H�g�g�l{���	���ou�aPtL)�uҌLh�	��?Z�4)���6_دE�|9�q�4F����+(- Fy�b��1%cA
����f�ih��{媴�%h�Q����o�]�߂M���c4�<H�j]���օd+՛�~4g�i�M�;�+�O�+�H�$�;���1����?��O�=�D�d��D��� )7�'�����|`�~�m�Lh�af�E��y*I�l�ޏ+e��
���3�|a��"?��r%�=1/C��:����I�q�%���~w�=dU��D}�(�� Zo�"i�.���/)��s�B*�=-Z��{�EI�kc�S��+�����7�t�-�_�-�C�������s��!f�DT�5���z�Ŋ�4(�i{�4�I�s~�5��1���G?�h���.+{;g� ���ٿ��ΰg]O��ۘd�ߙ�V�lO]�����5���O���de��$���"�f-�? \)�
��-�[V�d�VmJ��Bd?G��L�z����e6�2���,��PS������o��n4����<N�䛝��Wl���d+)i�� ��M<�e�'�'�'澩�h��>o޼y��͛7o޼y��͛7o�>�g�ou[�-}A�j����/�1������\k�O͋�ԍ�	�ڛm���ģ�ğ�y���$?j3���8��ɾ�����5��o|�q�͌�p��~� �6��F��!��8P�q� ��g�n�������*�|�Z#L��N�;���  =7����'�5�s?��֐|Yb̧�M��p�1Ddʃf [�%шP�I���cD����;ӗ�6D[`
D������Sq:ݔ�W�g�������veQ�5[K$��E ���D���)IB23�nx�����D��<C�/!�3BD}��/���oI�6�+;��D��q���n]v�[FI��i��t�S�ƨK���~�W�t�x�:�m��M�&ߎ&OH`2Z�h�-�Sk�D��Az��R>�3������_����xC�D
�l��]��S���%DO���ڄ�]������Qh��A��L�Bm8�c�R��D��T���vVWW�͍�)<�iDh}$.L>x�O��0D��C�B��:*�g�"ǿrC<�����s+��#>�E!R�]������~�qz�"��L�6�+����]����O����K��iaZ��P�u����4�vV�#�����{ 5�m��l��9����{���83ă�]�yBn��gBި�'��~N��JK�u8�c��W����"EtN�~��5C�����D��������<�o��<N@����ut�ȯ"�6����0"Qf��^�*�$�9 �����kKҿ�}�\g_��c����+���Km���&M���R,W����yL��h�r��k����/�.�}��&�"�������I�&伅D5�y33����� �C�7ӆ�,�	}����T�K%T���1�hlm��6֥5��V`4�䄥���\���<�R���ZreD���	�
Ⱦ�<�s�}uh�M5����R�b=D�-c�x��g���%y�\^��!�G��'�%PJ�t��%!��<�>�K��b"�_t����P�%?����O����hRa���2r�ҟ�����/~ d�ND�>E�;�G\$�}�߸~V����?��<e�#��̷ؘ�L3v?�3�z��-�������
��"�tjnJ��Na���o���ښ����=�����9�\~�t�R���H�w+~�bfϷF����h�{�c����dE����D�T{s���'��y��͛7o޼y��͛7o޼y���}|�K>emGH�4߲՜�Ag ��B�|�.�Ыd�]!抦e��������xM��,.J��g>�O<�d�~�翪�3���軤��3���8�F�����|�����3N�ӻfW��`��ˢ�Վ@&��	�gj�Gc����:��<$�rD{\.FY��Z��F�Ӛ|�/޷J��7�/��/$�X<)G��4�I$x0M4,���05�-�%xF7A��Q��J���|3N5����@G�w�1@��k�����O��Ǝx��Ԣ��,bt;ԧ���֦��!�H=#١��ASh�x��6�����p��XY��64S��1�<�C;�2���0Q�v@(��[4X*h��Y?p|j3O�"�Q�1��!�ED'D��A�h�Ä�˨o  n�_��������g��r��}.�ɇ5|92�����m.��"����'!R��Ȅ�N���Fr#�����A�Ȱ�4Hq��f��n"���)�������Gy8(A3�C≼�7���X�@{S]sw�!�8�_�[�?��?�ө���_�)!Cˤ`��3�l߯~)�����0��h�Y4�
SRO"C��?R[��5,��$��"������tiEڭF��䷃sq�z?��:��ǘ"�L}`pìj��O�R8�q3�Z�v�2�ڏ�>�qM#�)�j�i"}��<G崙޴f���5���H>M�+��W/]��FM����s�;����N���yh6�P��*�yv�A����o^����=�뛈�Gԋ�BS���R-��g���>�م�qJ6j��]`����f�������Y.`}]�ouU���]��=��k+�;��L����Ўe�WF�5ёَQ�M�dCV�v�4����p����-h7��'!7X��mw`��x1{H�F��"�m�x�*4Z��%2r^jr��G��?��Nڶ���#
����_|��8}�u�N��!Q9K��`�AfzF�Ij�p�A�����I4S��$�H�ԡ���k�������E�}ڵW��ӕ�[�R�(�|^��ZQ���!� 4���q>c���`���ДܟMh�@4Qڱ?�ȁZ-�Gmj�c[�r�_����g����GxrF<�n>)��}L���3 ��Z������C��M�j�:=�:���7�����+3��z�=�����c��=����2�N4�Gb��n��q�8#D�;�D�nmKƏ�*�f�`'����	�1�9�����	5Qg�8P�I:?/��цe�8�~�s��\A�5Ƶ�{깂fb����?O�y��͛7o޼y��͛7o޼y����/��)��O�R[<;D�Z�����/��6�^_r���3qZŎ�h��'5|�P,�%�$��-d�S?���(^����鉇�Q�Z��y��Xb��,:�����5���>��ۗ�����y�c���4M`���qzqE�Ѻy�Z��\/����|�<s:��1����ߘ�x̗ԇ+o��y���gģ�/ �*в\��!���&��f�a���5�uc�><��?.��O�ɇ�����D_rTE��yӯw���#��@�ԠY�zMȖ�n���/���V�������?�ӣ ��G��K
���eGC��#��� ��ǿ��^~'N��g�	�P�U^�j)@��DQ�v�֑@aoj2�A>��$�9TQ(����Z��,��J ��=��v�]z�iԨ�v�<�j�H����
<N������&RB�?�P~h$2H�eA,����0���Փ�5�q��G���?�������a�Bx��f�ьR�e�^H�dH K�;; -�7	Q�,��E�Ӧ���_S_X�#����"�g�83���k+ⱟ>"S#F�dm0����mJ;�~���4��Ϩ�Yj�)�\���_�?���������>��8�Z.Yj��>f\��K��y��5�@N|��h*nnJ{z�_��|���m; !�5ZhH�x��ߘ���w^��uh�Pc�Z��.�qET���Q2��̨U|���8}�IY�P�V�C���8=x�u���`L:��0���x�U)���������韜M4�\�N� #���ף�ۿ��h?� �g��?�$�(F�D�gj�gί�a~T��p$��~�W^���B ۈ��,�}�
Y�����8�(��K��ُ��C�Wq�KY�;+��{N������qza��^A?l���FHR��O���!:Km�;����Do|��G�Q��N#E���9�+��0������,X��?�|s���ҍ-�/��Ͽ�����8�!
1�{�_�F���F����1��:���!�a��xcK�-�G��?��/|����!�j�9��D����*����Oη����̴�������cTv�k�z��h�^�!+���o�v��+ Ǒf�_�L>m���bV�g�ۈ�Km?nF�o��,��g@8>�h/]�y���~߽B��<-����C�u!h���tWR^���/3�GLM�r�PF}䤌cr������}�!ױX�y�3��0N[]��Q�ԗ��~@��!VBؒ�)-P���o�Y��{>�?|]��5�2���ہv%��|n2ڜ&Ls��K�9�is َ+�B5�Hq�<ČK�[X�(�a�Z̲�!�)ŋyq5��6g�����,��o�<���d�f5CbX�7b1��?�*S�_Dp��h$�Ͽ#�N�9������ydj1 �d�q����+[�O�l�J����t�9��$1��W�x�ϛ7o޼y��͛7o޼y��͛�l�>�'\��x�y�'�<Yy3��E?zS��Yh��Kt�b���$1�!=@���A�$8� �/^�7�������7���������G�_�������/X'=n|�9tmI4%��=!?�	�6�����G2p3�� ��|��;װ;P���kǚs1�|��؇����O���_xQ<�;�R/+U!f���M|���Z�4�=Ƒ��e��)QE;Ñ��7^ȹ�$zk-��ߍݕVS��]QG3�$Ȣq5�ڂ�\)�|N��vu���F�=��q��ϊ���!���|�AK(Ef(m�<�1�9_��/��|���w��ҾYaS�lOF�6��>t5/g7j��=� �v��AeT�6ȄMx���G�E�6�o��D�3�b��@����#�h>�ӗ�y@�����K��!���B}�.����o�	��E:j6H�<��ShMR#+�4/q�mh���k��L�~
���p�� ���Dۗ�15`+41C�_��8�q����~�v�A�h�%+��y���M�1Z��$BX^b�Ӗ�~EƵ�'N�~�G�z��6�A��|���i�lڡ��G��,�8���8.���BL<���A3jn�-$�	b��噵��iφI��>&׹)���[ϐ��R��@ʁ||����_��_�ӏ��P���Y�a��bQ���_v�Wc��N����;�Ih,^�$��z����;�tn^%j1)�4��_5�x��Y��x�g�#D�ֆ��RU�]g�2�Dq��G�Y{�G���#%�������;���m�����~$�����ikmS�OD��������gyQ���I�|_�x*'��/}R�<�`H�m�������ʐ�RQ���?�)�����7.�-;p�4�M����cuD��Ǹy츐tԄ+Ըf�k+�&Jm֌׬0vɚ�28OD>�%�8H�Yj���$}���b�羇�qf
Yi9�}"�..S��w�yI�*���kBz��������Q�iq��>�e.�a��8��������p���v���B#��c$!1/@��G�4��z�����c5K2��� �(jc>D�>�S�~�JS�ϟ���f֝��8�����\�˿��8=zX��\S����t������J4�8�̰�)�:l��A��x^a�\ƃ���r	���W�8,���s�����̃�����/�qe��� :��~��ٺ�/GdE��W����D�Hx�_��8�I���Ǽ82�IS���f��yntj�Nl��܌���A��bED�)�C����
�(�<��-�R��7�9��U����8��5�����&�����)�gqFc>����GX8,�tb"�?�� �
��i:{�sJ�m���&�� ;�A"�j�7Z�1��٤�8��}޼y��͛7o޼y��͛7o޼}l���򦐚{���x\�����A��mp���|��q��O)N(H\sHqb>�;���������q�
���������#�
�g��b�X\/@5Q�^��<(��'I��[��ZYb�GωG�+_�[qZ)� q����+|����}x�V��f�%1�X���5��g�H���yC�8]uW��&�E`HCʥ��%z�J��h���d�3z�X�IT�I/\�
�#M'��G��K��=�2x�i�O�ēx�xJ�\��d�!���L��N�"�RZG�<���C�Y���6��m��%!�.�)Z_�)i�_���u�8n,	Y���}�����a�cjJ����A�SB Q��^k���s?��8=Y<Č"�25s^{��ٲ�&�eOP;�ޟ�7]D��@�(���nێh��C�&��^��d��aC�W���,p���%!�n�_������7�$���^�}����u֞� �� A`�!�JA��H;$��m���W�۔(�T���(Y�� �``8��鞞�}��ڷ��L�y�ߛ}O�[����Z��P��{�ܼy����+5�iH�����&N���T{��.�?Zߒ~���7����j�5�ۇ�a �5�%���m�B[4�Wv{���2�������ZIͶ\����M[����|�<v@���o��O�;�x}���x�D?����3�^�x���_�vI"�"emAH׿�+��s�n2�	���@^�,��+�obB��ZM��R��������������w�w���}є*R�ʔ �}��hK(�R���z�f�'�����-ZZ��1:�*��!�a��(Ř?��l<H-/hq]�%�К9n��@G�u��k�>Cւ��X�J=x������S��|�w�x������g_���J
l@�Ѫ��"���e�5='�7V�z��/�GX� 3�}F��/��d���q��'�0H㊩���3��Қ�6qI2`sU�����=D+�A������u��;R.����2�i���n��\B{����a���s�"���#B�P���%�}�p��٤W�K�&&��(`�y���_�����$�m���E��z�����'R��!�?�-k�H�+$�BEU��~�  ڶ�I�����wJ�9$�$�/�'��E��ք�{�g�{���h�BC�"��}B��7�/�P����������q�$!����){��U�1D��'q�'B6���&��$�����;(I=���{�ޒ�����ɼ���0�� a��Wf���h����7T����z��|H�t:r>j>�*�;y�G��ӿ��/���O��(���_S���UQm��!i�S�|��h�51
�o�Zْӫd:^���W~�i����ȧf�h;|���Ĝ��N/7q>6B���vua^�53�2o�j�lp��q��@������������8���B���9�h=]w�}&���w�Cf�|[�G~�{�|���y�D�V>|�x�reM�$�M��v9�~|����Z�υ>:ޔDΚ��{N�<��͛7o޼y��͛7o޼y����}`#k�m�����}�<��dx�?��MhM�sU<���Mqݬ�V��������ς���;�8b�*�{���M�ӏ��lo��!0�^!��������4�Q���_��hn@�eD7��Lh@˅�҂I�qH/�bd~]H�6��ry����*=U���l���Ro��B���h�؞�-�ۓOɛ��	��I۷W�=�88Uȴ��E9P͑/�ގQ"�E��2J��âm��_��qڇ'wvL�1o�&|g4a���U Ym���W���[B�,�B���8���?���&Ϟ�����=N�'��y:��
��x>��'N�Vᡣ�z��㢽�9 2.$�n�v6D��;�չ�dt9�����h�ehV�Y-�#k4�����_s��A��QR�+@�0`���ICҊDE^&Z�7���Mi�W�\�v�!��&��MAK��c��ސ~�=�8��w�����,�zAHVAD�I���3ɉ-�krF����M��i����H!A��Q+��	��z�Q��$���2�'�Nڋm���Yy:}ǎ��G^����٤��M�׮�76%�TQ�IN�B hwh�%�ϟ�����N����S��A��o�v}cM]�]��R��o��B�>���qZ��O��$&NC��~𶫿�4�H��4$ҹ������o_��e�*�:��TBt���"ʯГ�A�ŋR��LK9^��m`<�Ȗ!�mb��I>m�z��@v���u�}�c���r��p����b�D�ƆYҲ�zZ��~��?)��פ\J�=�{�8KMO��[��d�5�;At���Ш��bd�,�´�=�e����PmA#4���G�	���h���&W{E���B`�����i+b�P��/�vqI��e�[�:M#�y��˨�G��&��G��/@w�ܵq)ǍM!677�3�	C��S/���Ԅ�Tр�·�/5f��D2�'��P�&)�@��R+D7�5C�و�����}hخ.I��*�8@���E��Ez�8��'U��J}\���<�=��nn2ʯ�wmK�1FN���v(��t~پH�1�*?j��_��>�Z����u^�-�?��I�QC�1!�\Ȩ�(��'�����#$*�T��d������e�����}D4͛m����x}�����!2G��N4Rmm����9��*�Me>�mmr�g+^f�H��y��>��)�7~$+�>��G���<���
��J7��N�8`���Y��H>6��~��N�J����g7~Z����ʀ�+�r;��y�ߐ���`�yϽ"ɕ�-�ej����ƙ���=�TF�F��"�3�WC�����Ǚ�������^��W>%��lq��fQ�?�]ti��-�/u>�����>)�/��x�{���qZ�<��t��{|�{����:�~t�����F�o���>o޼y��͛7o޼y��͛7o����E�r�+�Pd<f�#~W8� }���?��G�ʛ�<�T:�d_�Qc���/>!��fgţ���_�ӛ@Y�����̣B����X�~{6s��Qh��:I>%Fmz��X�݅��O
����	xZ�³[UP��$V�M�{fc�#�Ʃ���}�����uc#�:O��)�	>�Ub4Rr9���9c����ݷޔ���'A ��h�� M�e�^yP�����h����x��8���<*�ó�h>��@O��5ǘ���� �ifJ��{7œOm�C3B*����ӈ��ڸ�&ʯ������Ʉ�D�^F�����57�c���r�������ybt�1D�� zk.�vңU��;�#xqA��~ߎJK+�D�օ���E2Om/ٮۢ�5�����1I��$�~�W�>C�E� �#�he$�"z�������u���2D�؁$kn��T�㊇���<�|.ܒrc�S���Qɇ�\�I�O�iS&Q�h�3�"��c�<��S��t�T�0J����E�lN���Ֆ~rmE�]��X]�'��$<
9��/�V��Ҥ��A,>&���}�ނⴌ��H�%����ه�I��M e���B2��_��yOb��� ��������D	��m����������N$��c���_��C'��55���Y��l"�֗�u���8�Q0mA�[�O9.�(l��� )9Q�q�>��|��G���tM2�pQ���$z�\�l��xa���?L����.�^P^w���1�rA?D�-hY�*�Ba�!����M��	��'5�ԊS>�5� _K�~�۷W��)$�9��q��$K[��|w��%�1�d�I�ρ����+�G���������ߗ�=�(�$�9�^�&�UZ����?���>pP����t|�|~+"�V�]�)�?D�K�B���Ƒ��{�`�OI_2K����DԈ�]��<�V��+��X��^ RB	��nd��I�6A"67Y~�p��h�:jt��7�����v[���ćE�>��у�y�U#h��Z���e ���W0O	��&Z���$xI�E8VB�R�:-6.y�
(\G�o���=%��_�����|E���פ�-�>qE���'&�_�X�Jԇ[���2���;tTH�U�$˸=���u!k)�
��|��d9�S�N�����9�����+�$_�6�kC�Փ�V��>,D��cBܲ5ދy����?�a!�K%��Ӏ�n��5~��|�>���R��-��efJ��{Zȿ�1��U��<p N�X�W���~x�h+8~���ۢpۦ(����J�ݨ�*��.:����o�MBc:��oj}d�W��i	5p�}�>$���#�ߗq����ӟ��Sq����q޴"v�縻L��΃����ii+����q��gde�$ڥ���?��T>m�_|���T߼�h�1O�y��͛7o޼y��͛7o޼y�������>�Ꚉ�x�"DE�Ή�﫯�q�~��v�"���yG:��(�>�C���W$=uQ4ν/��kx��wN<���'h
�['A��y����j<A[�)+�+qJ��-h�Oɋ/�����I��m���~!m�j=my ����E�}�2�Y���q�"�B����-z:I��$��	2Y����7��}bJް;"�D;�D�������yQ�0ZU�.�p\0�w��CzMT+_��/�i��K��.�DAJtC:���Kbe�����2��|F�9O�n}���w$;��C�/!��A�0�_���ѵ�9vDþ[�i��#�BF�pmm�ޞ�A`�9&%J"���t��<<���x�鉯���A�"	�M0*=ތ��i3���sdG_E�&	��>	B-(H�޺&�Q"Q��v� ���T�󷷠�f
����od�쿲����LmJ��+<�Kr}� �r)z�'������u[�4f�Sf��l��ߗ���j��B�nA����R�}��[���Hrr��{/�*h�=�S �(��9~	Qˈ~Za�vC�#<��p^���n!j�����'���1!���Þ���aP�7�|�^�~�7������?�qU6y�d�{�d�}�A!'c���mQ�Q�V6e�ZIè�cS2_�.�?y��8�U(.d����(��{�v�4<���T����g�EW}D�N~w���k���˨�%��Jm�P�TO�����vh&W�ш���#�
q�q�D1��c�O)�ej6�9H�i�$vi����^cc6�㛠��
�^B0�9vإd��A93zp�(�����������y���*Ƨ��7��$)���$\�$�������t
D�?'��i��K1Lj�q�Ǖar�rK�}�EԂ�_>_�RS���g�])�����#���vl�J�LvhLHy�0>W�Ro+y�G&
�"g̼h`>p�C���G��xrvҺ�VW��Vb����{h����Լ�
I�:�-G�z�^!�U��+���u��7�"N'f@ zȿM�1jx���)Q���|�ق#F���H�q��y�8��*��Mi'�g\���z��"�EmR�g�ʋ�"��rk�������j8O�����Q#�{Q~Qw��R�"4.O��籣��<������_ ��������8=~\��.��h��sJ4��@��/�[8�Y��1��j�j "iq�;�_����fnV�{&d^Z�1갔k	OB�LM�.�����n?�ܪ�f��H�C���*D߾eܧYhhc�
�;z%5�˸1�����#��:����r������GEC�V�h��ݒ}Y�DѶ�`����!7;|o#�|�>鷞|P�;S�Ϙ���$Cz�%I>*|_F���*�0BZ�Ý��f,dLL<��͛7o޼y��͛7o޼y����}`ۼ�s,�qs�5=y��(ˁ��d�Ο��8��O})N�g��pJrx,�;�N�����%��� y��hI�yQH-�F�"5�L��5�:V�����'�z�a�xHH�
=�	0�*�ׇ5�,xj����oAS�ږx�ZEx�qgS�^���w���hy��G�r�:�z��Hy�BT���ǫe�d�2I,) z>�F[�!�I��ZB&
&=��h#J����hy��)�/M�Ǒ`�Qb��`v*�`<>��o��		�.����]�²ԫ3�
!K҄�.�� 4��V�s�n+w��(#9����B=��h<PCAsEh#��d��f�6�	o'�Fۣ�^����<�&Cs�&ǫT��'[�F�~	ZA!J��POp���6����;I�<�"z�0@=+Aç3����ہ��D�v`�k���&/�O�7:�N���K$ӯH�������h|[�{���r{l����HuS������hU��zO��E3*��h0�L���[�a�S>p��:ۼ��5�]�߳��6�Xb�f�C����	b�7��?�S�r'��q�d������5�����9%��̻Bn<~B�{	�q���q�gߐ�Ǐ~X����̋��$�(���6@��A�r����.�0(#�u�)�(�+B֓�њ*M�O���U����6ѧ/d��ەA:��"��r!��W��"Mx߱���K�ocM��B�րJ�q��ڐ�8H~�����>@�Cr���q�T����ve����v�$4�28�h��4�At-.Q�}�jӼ������qio7ׅ$����{_��h���x��B���h05@R^<'��&��:tE�Q�����P��� I �J>n^-��I�g�&�@���u�n|\H��7�幀�Y����}�:$�7Tbh�|+;@ڗ+r�J]R�M�G5����:�%RO���j/"�
�ȾHi�����2��FR��h��xk���� 7+�QE}e���oK2��m.��A ��dmOB���B�����*�1Wu;�$�񹇕#��?p�:4w�X��v}�9���ʭ��x� �1���>xD����j	u���f���O���-���M9�VN�}���Ο�)WƌA������CB^�f�^}.��/�XrE"�������*�����p��Y81�C�/�`����.Vpj�iS��-rw�8R���]�'�5����71Ͻ��d�x�84.�����?��'6�WF�>$�7FT���P֯[b$<��J>�֩��cs��>s�ř��%��7����"++�.��6H�c�$��=�a+_��,�.#"!�߹,�c
�l��x߅�:,��-w���͛7o޼y��͛7o޼y����:���/�mOn�$o��P"1Q݃���xh���D���?�edMGS�/8�]�hPIB) <����#Ho��x�2�n�TZ�%k����MpZ|CO�����7����(��D�Q}N��F�}�,���>�� �w��&Q�����c���v�9�B�ԫt�O��\��F�Gޝ�tY\�7�%�_yx��}�`lmA[����k`���K�)�pSAsU�&Ͷxқe�|m�3�R$�R���Dm�0��� ��%x�-�<�@�Q��DM�� �Ѷm��~��r���wJ����נ=s�@$077-:gkhiB$��<-�D|6|�c��M�AWTD=��Sˏ��$�e�tj�}�甞�2<�Ը˫�Аq���<HC�pG��d�F~Cx�z]�#�Ŗj����"���J���r��E��f`�r�D��`B���)�ó|CU_��W��S*�܏�]�H4�[0�����s8��k�Q�a���H�O�0�l/oR�D3�t�Jƺ)�=�V����FkA��ڼh�샇�)�j��/H�(GC�?�����ԏ�x\�r8b}��Y�l��ڒh�� ���4���y����vQ*Qo��BH�#DUTQ/y��=F#��-���G��I��<����{FY��c�c��������k4j���Y^r{��s{���8�ͥ���� Y��	f���:���������V��源����Sj^h�9��8�ۈd��2uC ۩>/�qr���-�Lx�ylgGѦ�3�p�5h����Y�?��S�h�p��"�d�����q!4���\�y�>~� N��D1f�&_j�>���h�9/ [��P"�2Y[�zу�n	D_D*ǩ���ifR�������f"����S���.�5�y\��dn	;{��iI�p󪴫-hS;����W��X�&&ǭr*a^��
���H�,n  ��IDATtw=h��,H�T�8�eV���F�\���7�\�5P��"�K;�m��h�h��Ø��{dep�Z �0��0��J�u�E����_9^h��hwS#�Q��Nl��̔�^�h�6S��Ֆ�}c^������K���:xP���}W4�I��Ǭ|���m��(k�@Lb|��v}��B���ZM-fEؑ ��ٶ���sz�Q��b����@i�}�_��d�.��$�c�C�5iJ�$�/Ⱦ�"�>���/� ������]��\�#������\�ƽ9]��R]��ݐ��-h���Ȋ�&���=iWO}@���1��9��ٱ��;�|9N����q��T�1k�+w��'���H�y�ϛ7o޼y��͛7o޼y��͛���2_�����=�)s-��G�1'�I������%� 6.ʛ��.N�8L>�=�&F���|��*���#5Y�~���+��I˝~$2�ɖD!����YjM��ȯ�_׹8��ɋ����I�5(��S�I8�d�+u}[�L�'�dGMD�x}v��Pyt��#����w��#�m��DA^y&p�&�"2�3m_	e��6��A#�֛���C�ǐ6$�q��S�*c#��1�����}�d�?F;z�0�#���1�~�0��[xR�#��!�
@�
��+��;Է
Zvi�v�/�4�X4��&�ׁ��U��@�=	��S���U�$Wk�*�eS�&�aj���jH�}�CF�s����=�SQ�����`+0�b�����:�B���"�w b!0�h���@� ��X���ʓ�T�I޴K$�qEk!�$����ѦI��;�ꡇ5 �Y�4! l"1E�h��d�?��e*�|�D��X�è���ct�K�ţ���
�oH���$�6�3������i���!fq�%����Yg�h�9�!�*���:phɮ�_fBms}��ΐH���߯��k��F$�a��9!W���"_���nY����/��¢x�In0?�����W7�����J��|�$�R�w�*�&�h��_��cV�N7U�д��y@2k�;,Q��*���R$�&�pB�g%�Qӊ�e��S�%�fo�n0�P�O�e��Y�bH4l�b�ZO����8��:ߛ���Uj�yo��[K3Iq��26ha@kk]@���o�<K(��17VeE���i�!�q%O�Hd�\?��\��	 �1�����l�܇A�h�������xE��Y�(�����¥P`TYλ�W�Mh8n.7����6i�ޕq:����gw�$�y"��,jN�o��~�{<N�͵M�'����� ";��u��l%�5S3B&����`�yA@pUIͥ�+��Hzγ��f4�;Z�;������׾�O<)����/��$���^5�g4n����E+���rXY���47n��f%����	L��۾#J���V��F�/����y��57��8�㳙�8;��gv�b��v1�w�|�q��B�M�l�ہ����F���v����?�R�����/�����8=x@V���+ڴ{�?��k%`�e[�9�-�dZ[��amM�S���?5+������a�|��3.���uv7;��|򒼇�`Ee�ƨ��#���L�3�z����U�L��>o޼y��͛7o޼y��͛7o���|�GO��R�7��Hk�z���L�E1<`I���f��~�t����O��s���7�ؽ@�`�z�7�p������76e}v���l��\$ �
��|�o�4|Z|��e-z���ɗ+�؁�f�]����dj�֦	r�yp`.��8��bOk$�R�'�"/X��/�D�۩z��������'MУ�,I���VC+M�v��q?�L�H�\V���#О�MB�لg;���%.L�Kh������7�^ק�p��5"�ni�0Q[g�x�zMxv+�V+�i����Q���#̨��{}���Pd>�Kã��q�}H�>��٤M���R[&
��F�l㾴�1S��4�=vv}����h3��a4�H83*m�!�oK��Z^;6���%b�nH$Bˮ����Q�;�$Z���O��m�����s��H�'n����7y}  -����$�ڈ�YF�?3%�~F���N��Tڇ����7�]��O.��QD���J��̇C6EL�;$i���u���{:Ǯ�Mrek�ة!������Fz��CK��d>;����D�h���N����D��7$i���(E�w�-ل��@0r��g�b}d�H��h�,+���|l����X�����40��A���/6����)���&�+���Ԋ-�U�f��7��[�(��~RD�!-	�~�	�5�OF��Zib ���nw�&�?G�&v;�?ϩ��+$:��+�<W>%�nD�����M#
*��r��
"=�������h��06+�*��hO,/jŪj�~s��<�X�9�f#W*�z����R�okm��1IHj�{�����Y�@�Iؒ m^�5�Z]�G�M��sD���g��Sݏ^Y�|�\1_�0��b*fGd�a>D�ʬpp���2#�#���pj��m�:��\���	�.�Ef=_��R�$� 7�;��װ������tY��B*�f���)�>򤅒���rn�^!�:]!��ׅ��vMVr�w��m�O���wr�F�~~�T��cE���ӹ9!g���ԑS{<���$�������aea����s���YI������	�h���}޼y��͛7o޼y��͛7o޼��M���G��[j����ͺ",�W�v�<:��Jh�mA���y����|8N_zD���V�*��$�h6i�Z��3�nb����O-�&��#|c����;�.�������\&�
���K��\��֨��֠q�T��(����Ѥ	=5��0Ɲzd�y���������FCN���s�zn�W���7��(�;&7����m
Q7Z��dۡvR;�9����'��Q���C�fzN��<�}�D=H�(B���?�B6���D)��IEzf�Ӯφ�ˊ�hL��c����W�2��.UMb%6��d��v;;-.�K���wAFPs��q��(���/���.7�o�Hĝ��nM8�~�2�+[[��ۈ�R���xԌ��9�#�P���%T�DҼ���B�ڊh_�uC<����u�q�D*�ld�c�Ӝ��XG���k�y�y@V������Hz�Zp�5,I�ck3���$�t���uf�s�{nx}���&��� vz��ǝAhG���r�!8<���"X���.rh}�B۰���P}�OF:L}�ۂ��)!/��-�.DNڈb\�vk�~DlbB�å�e��]��#p|�v�&�>�c�gDY!��3nm��+f���mCX��$Y�د������Ū�j�u]5��1�q�1��4w{�%(��3���φ���	r��[Д�6l���1SM�YY� �bA�S1_�u1Z5�i8�J��h�
�xe��"�L7��Kh��/�	?���|H4R�ьo���'{Y��� �~�R�6.QH(G>�������\E�tT��|���Ev9�����g���T�5��x���QZ��4�S@1�T���r����%6|\��W���em�����HwD��y�vy������I�o���Y�zu~UȾ>��G�웭�$WP�{��ʝ"����\��>=��}��������⹉�1�b.��"Jw�*�V�,�
�Z�e�z��"�T��[IAsV�����;�D��Қ�@`ee��Pji�7+W�,����'�t�2O�y��͛7o޼y��͛7o޼y�vX�>�A7�zn�G�C���˧�5�J�'�9+��M��ފ�w�������C���W�e&��f��Ni�\�7����E���=#9zPe������$��¦�i@S�����P1�$I7�ʝQ����!�yJ�I�F�j�Q�e	�@O�p-(wX�\��w�lOK!��N޴[��O#��������]�Y��J�wEjsK4@�U�y�T��̳���MN�GOy�(a�����ev4WF�=r���ĠюJDB��_v�Ɂث�3[`@�j�"ۅ��:j��[.S}^�b���$u��&y	΁M>�/����c����(��P�qT���lF+1?��'�㗭��DY����>m��k�A��	*'󈎺Ҕ���u�>�ȣq���O�)�u�O���I=V����1��#�n�<��}<yZ����z\�D�T$_j�����L��no�f��@0|\�94G'��yS^kѺ,k�q�l81�czkE��;n����-fީ5n��50
2���yU�sl�7ZB��V��*}�z�u{{�q��y��E뼉V1���h�ʉڼ��%�~QN�҂Qk�f�M��fc�X�O�r�J�R����͜���(����ѐ�)W���hf�d�6o}���#�<�d��:U_"OEj5�ۦ��s���X�)DIm\��ZU��� DMP�^�O8�U��*��\V`��B>���̼��|��|.�{dF��B��c9��x)�����ʃ�������m@����r��JE)OVKC j�W��*'���@�'�G���\y2^ݯ�%7n`�C$��`�_`;Wρ�χ~r����|9�ߩ�&�:����IT�ᤧ�����a?��>'���V�3a�T��x�y&�J_\B������qy���_a{�M��[F��W2��~������#9�ok0b�M�n��zï9�'g��Kqz���J@�<_��'$߽}���8�A'��=��͛7o޼y��͛7o޼y����}`�D�Ѱb�j�qךpZ���v���J�%B����"x��u�q�������'���Dy���*�3���	��y<�ٷ��t|n!��zN<�W�o�������JS4�Z}h��%�hqP;�.�T�����������7\�X1ڦ&�L� �R��uTt`z�ʃ)�G�H�
}P����h�j��ClG����I5�x�R��ݹ�2<�++��7U����qz��hq=�W�1h�|�g?����5N''�(��o4��m;��X�,	���g.N>�-P���لfM����3H��@�,��!Jm��]�F/�{��Ė�����YF�	yC����3��T1��+��P:`��Mk����7���:J�\������v�C�ڎDQʧ>&�-�Q���M���8}��?���|��q��.D����}|��d7Q�Ѿp����~�+q�(f�~�f��R�36)Z,F�w�զ��h�q��H���H��i8��=��Ps�;G;Q�Wr{����g��J�ͅ��c���]^\�ΟL�"����7vh�6U4� (���D��TsVXubM�h��2'"�ڐv������,N9:=��#q:;=�&ʽ����*9��k�-�����"N9_�a���)!t+�'��A���)��3d�c8�^'��prw�y�v�7�~}��?�8ݻg6L�)��X@�G6�N�:jk�ݥ�e��Ŷ�B�e�k2�����o�4[�����#�/Q_ƃAG�O�(�A��T>�+��?��������e|������Y)�H[M�a��.��ͅ�v6@9���e��̏}c�N.�>!�Ri@#d*�4窨���/�u�\Q�}1�Ҧ��C��s�8�<�ӟ����G��[X����J��v�{e� 	�_��Ծ�������6�ͬ�3��T����l?�������{���"��Vd���x��N��[�&�T���Ў�x�:�"�}�����!�P?0)�1D�.�y-�����.�Uj�����ߓ t i��8�4I��P���s�p�ޖ��������h��˨EE���:�.lDsϛ�{Ҩ�=��͛7o޼y��͛7o޼y����}`�/�H�h�;-r�|9�5E����=�4s�	���^��uxN���~�OⴑO�4�N< �褬5�����9hx�3�n� �Q������"i�%D��x�.ܼ��v@vq��w���Ã�#)e$;l�F�<wg�B�R߫rPZ����8�}y�r���&Co�07��b�(��.פ~��r8���D�SQI��}�Ik�7HG��F���)K����w�����0N���S��Sa��?�Z�.,���@�P�h��%z뇞�M��w���x�3�N�ܶU�(L�;z����v����r�M��rY),ã�7Z6���Y3�gzp�txP�-a���>�c@(��έ�[j�@i��\��H
�@�T&�8t(N����Č��o}��8}�Q��:�(f����_�_���$�*�N�eӈ���Ͽ����5�p]_�ӯ�i�Ϊ5DU� �R�9��ۮW��<���Jm���%���Q�?�!$�$���̐|������ʹ&�����t�����$y���� _LL�؍BL���d+�]}���/��qʨ����gϝ�ӿ�����qٿ�eTT��h�$���9$����~.Ng1&��n	�q���l�p\J �
�
�r`�J�Ok{�X��'�H-@g�V�#��84~zP���I�Xu0��泉>3O5�pFC���eY�E�;��Z�\�0�P^M̓H"Ai�F;���������w�N����@�#�����C���{ �M��h��J���1/��u�د�Vf�(5��!�x�*��Q���2M��	)��IiWc /��zT��Z�5��F����i��/�]�"�kn��/}��8O�:��w��i�/�W.s�=��ݭ�T��g���O����F�ЄlN�G��w�R���������Gt����斬��^����}ơiY19;)�:��8����\���Qؙ}��M����	^o�d*�o�%�_�g��w�	�+Jse �+�X��5��r��|����=��͛7o޼y��͛7o޼y����}`�/�R�$��O�H��DT؞&}4E�Q�pw��&<8�B���t{��S����q����qz`B�q�%۩|�MD�
H�������پ� �s/^�5ݭ><P� ����#�e$������wz v�&Y{��HE����h��Z |���@��380��:��Jɺ��R>��w�=�W�'��~��e�]�TE]
Q��1%x�{h/��@�}�[ߌ�/��f���{�8=�ē~��q��.��;�Nak��'��h��ӧF�ãl���}���#�|*N���%��v���q2`���&��h�kۣ��m��t��Z�Zh�`�[�+c,�;%���%~Lh,��C�ۤ���d)��� (��A��2�A��X��M��km�G�2.��7����׾�+�=��hg�����8�����)ۧ�66��_���3�Ɑ n�v�Dg;sV<�A	�Fd�_�i�P�_G;J}�=�.c�f���:��	5=��|�j<L����nYZi�fLn�].:z�]����v��FW^=?n3d8�E�QQk��ݶҐ�}�҅8]~Bƽ��D��d��z8N�xS��ހ�L$���<Z�ف��V������]�2�R�/��U\�1��>4�'&@ v9欔W��l��=��Z�F��<|E@B�/h(�AW�3p�Ajbi�C��'�A��1�\�u���4�f�ޡ��'�ꡙ��|&�7�K~/��}��m���Dò��A�_r���OEb�/:zo��l�#�ض��C��
�%Hb��!H��yG='�%�G�/���r6�I����y�o����i�׺O�<�cS��=c�_�Ұ���x��ۏ�Fw]��%��R��ϧϣI�?c�c�{ڧ���B���*l?|/ѫJ;X��|���U�P|�+�O���k������HH�i��T?�SBzD3���<���������2�.5�dp��8�B?�m�����>Gw����X��y�ϛ7o޼y��͛7o޼y��͛���F ����F#� ��,SS����؀h3)|�g�6{m�m�R�+1�I��xR�ZB୼'�3�ދ�ZI<'eD��;<Y�дA6l����Dډ�4 y�����>�c��pa�$r��ȍh��ϑ��P�"g׃>4c�n�o	�b���9��Ro����Q�����%P�(��ޘ+���L�S��$�8)�CO��NH40\���<I��Dz�!�ysY<4[R�������ҭ8eT��?�!�]�S/��/=��W���>e埞"��<��]eh�ɷDcs�%��_�b�g�u!�[�H��GJ�S�iQ�3�x�w�Q�a�htY�@����|Q:���RT�w֏�M\$����{�,W�v���s�z�p�����s�F I�<��wj&��y^�E-!j�V m;�=�Rn�ȫ ���K���'�>��ˢ*����B�m� "��C2�ڛ{��"�b���N���?���ܤu]�7E�$�M��Y��'�՚!�b4w�������ŷ[s�??f �D�*���@�j�2����ʼS��������&M�ɨ�!	�(��Ǆ|X_�v&�Ūhl����wq��7ⴌ�P� �+�%N[-�ʺ�"­[2^OO�w��hw=z�#I8>&�;��h�����%?s��������}��uu�
�5�FR�Z��;�T�DNKm��Gm6�{�G!����NM�]6U�����9�*jy2_�۟�����]�uc���(��*_^FFEH����F|H��6�a�Z�2I�kOd.!����"a$�Hl����y��� Z.B������g����}N���C�^��8G�;��iٰZ�e}w��?��>�I��g�q��� �Ԇ��Z�>Ps��yP`�����R�
Ts��3�W�Q�(�v�?ߵ�=W?��&���<v���⚐�k�t=�+#g$��L]ƏZ��ܼa��=���eԫ���5J�@��$�i��}�{�/���K�~�+�b���
��lM?��[�6���y��nO�G��G�0O�y��͛7o޼y��͛7o޼y�v��/����|�'���\8�7��%z:����6<x;���+����4=O�-�����b�:�&��n��L�e��P�k�y��~*��&Ŕ�<!B�˥���qY.4�D�<�FS1Q�@>)���� #m����
$ݴƒ�x��	?E�(�,�MT�x�����j�N��$N󶧆���+�T�ɳ��G�YL�����YnO>'�tϽ)Ѽ.]���+5�p\�#ќ<��x>^�ٗ�t�?�������c`*�I$�������Y��m!DE�zV����S�H;mn��B�ն����Ā��52�����g��)����0�YE���5��蟕���͛@}�Z<,>SS��~��1:�֖h�u5/�!b���J��"�gW��L8�~	�o���~Jߧ��|�Y:߃5�������=.�F<tL<��/��lcR�����?��Sg�����|>N'��k���E���n���g�����o��%�jGD�v�)�`i^H����2Qփ����E�Յ���w�Q������v��6Ü��Mi�����0����&���S,���{����Mϣ��nRf�A����K�y������X�1�w�:�Ꚍ��~�ui�����V�~�������M�"�$::4<+�?��|�!���׾��俶$Q�����D�]�&$G9R���!��L�ID�5�������v�vF��2H�NǞh�K�ݨ5O��t	94�S�������;�V��?g��6�� f�������9^mӖ�p�N��*뱄�|S�}�w�qn�Z��>�)j�o��O4��<��	���~+��2O}蘴�ǎ>�K7�����%Y���ss{��}Y��o��y�[�e�\����[2i�H`�h)-0E����vNPw�Vp%�Ӵ��ڎ_���pbP�+]Կ��Gr4��>o���<�tx|^2��. ���V���;��#�� QfC<��0Qj�2n-ߐ�W�\�&�uY�ql��fd�H+'�r�����$o����]�Q�l����[F���{���qzuI4�[]y~��B�'�-�VX�>%�@�/����x��C,���>/5E��W�+&�
!�y�ϛ7o޼y��͛7o޼y��͛���F~�W�S{ _���HȻ�JUސ6���la�uD��ٷR *�����p�W��������_��#{
�l��h�(��>�#�w�x��jN��u(m��^H` ȣ!GI��Q�L�CF_Vd�m9W��{0��KytI���B�A���hЅN��G��N�GM]�d@��E��A)����%!�}hlB<��΋'�SK4BΝ�ٓ��DrC.����~�����G��y�1��;1114?���y�Wo\���������hK�/"*���h:$Q��h�8Pn=DI�_��J��0js��NO{��`D���đ�.���8�i7&���A�=�ݎ܏�'>�5h(�� ���%�*N-W>h����b�@+PG�e?��(������������	�o�S$��Y�u�$�(�Oe$ˉ�Y�d����Γ������{���vw�܇:��MD�_��o�釞���=��<����
q����8=�wߓ~`�'���@��@�k֯�i����͡\��c��$2���xv�'���1�Y��$SwI�-K��g
����mF�F�6I2ޡ�:j�lvt��}��y�j��~#�<wZ��W�Vd<`ܪ������|\�G�>�{f�𫁄s�.�~�_?%��{�GqZ��~��-!��m�*�ɛ���z� 0$25�8�QKXE<2�MѾ�>9�j���N�Q`͊�Q��HMCC�)O����؏��ջ7�� �\�;w���Rͧ3���0C��~{�9�He k�6|s�8�h��������}�U���:<����ⴠ�9��[h͎���� N߹ �paZ�)�u �������k�
s���+��
|���Y]d�c��qY��h��>��ɕ�Ȉ��,������]>}���*�˃��ʈ�-heηd�tA4^Wd>9R���+M��dr\�����W~��Q}<׵3�%�Z�\I���N�!�A��5��>����q���`��3������>*204��g=g�'��y��͛7o޼y��͛7o޼y�,�E_���M�4���|���Y��aeA����H,͋�.��]�%x�� jKIȇUD��&�o�#�ٞ q{�]k�]o\��4�zS�=YQ�v������DB�H�h$1�\�Ӥ��l�~OG��iTt^z�ӒI\C*�q�z� jL}��P;����s!���?���p�����D�u�ڃe{�U���0�&D0� ����+���G_��^x)N��=����qc��/^=�o�8�����A�F��m��+��� j�mmH��j����h�Ԑ�����e	�^��}�Ƥjg�G��QO����-rD��QBƺ�T�d􃰂�@�9_	M� �����眕fu0Q	�v\d?���2ʣkUλ�o�Q��knI�����ӑ��SZ]����3��!�h$-�EP`��7��F�"~�Q
�=>�\�~C4�f���9��qz��h�\���$4�N߼������*�do?Kr��O+ i6�U�h�����v�,�7۫6�pe���82|�p6���	��K��S���؎��cN�3�7����$�W�ȨQ/(�:M �Ĩ������Ҟ}eA��nd:�ɯ��q�շ^��)ǡ�����u�?߸)�B�a�Q�%l'і�<�@��M���^�$�s�������橩)���rh�>���ْt����kk�6A�q<�q�%[ӕ���H@M8eW�9g/1=PB�� �i��H�e��l��&����\��*�J N����W�5�p�%�s]'M�\�bʋZZv4R��XF��f�+g;N��ϻS�3n�<�q!��]>�;>&D��+2/����{&��8|�ż+P6�y|�̣��#i�$�B�]hr�,�ю�@r]���+��h���&�{�w������S׊��ڟ��{Nm��Z5���;�&���&
vj�èD�..u��]f/��1+ �0�'���#:|G�C�)�A�5����2�ʆ���|���s�5��+D��
�s^��He���A���&7�|��{è�>o޼y��͛7o޼y��͛7o���E_AE�-�M~��D^<��w�}�P�,	Y�_ �E���3-��ڜ�S�a�풂z��m��#�K�n��Xz�&t����v��i���$� �{�$���Tؾ���tJ���q��
�T��\ �2Q���O
ٲZN-��<�i�=/��f0� |߇�/�z%.�������MqYT�R�C:�����0����vA�]N����HCz�ǅx�!�橓o�iq ���	h{!{��G�{�-��.n��~���>!��j��ܲ�g�a��6�C~�$x���@�� ��^�p�����e��w�/v�S��)ۨD���s4��)�\_�	�&䟚�s3�ݘ��-���:.�}iU�� D���١�kO}�!�p^fQ�h�f;��n�*P��R���������&Z�Y7B�i|J�CjY�@�;!�]���\�t�#i"�5`y����2��*�s$����������<��N!�2ݐz�]n�F1W���w�C5�@�h�w7*�1G�U{/�9t����:���]�0�ނ�_t��~SO��[G���,�� ��]m�&�� �H�M�LY�7ׄ�]m�c?�kX1��h��)�]E&�E"��k+ҟ��??�P�@6ܸ.��X��5	c�D�އy4N�!V�(�l�瀌�qܥ5!�����+�q�QCEn��m��5@���!�559?U�w`��5Ѧ��ƺ�W�q$���;7+QX�!�=muE���-hP��f9V0"���6���]��Z���x����7�Ԛ���ll����
��e�/�uԬ�#�ec�w��r��cb�o�q]����"I��7=���v]�<Cޛ��b��
�+�\��X���	y[�|�cs�i�����ڦ�Gj��[k�}@�sϔԋ
	Ю/U��|Մ�pK�G��'�<N��#�/ш_��EI6��_(��H:|�lw��ݾ#�e]0n�煡�2�
L?���t��$_�h.q�`g���H��0��@�&ڸ=>�V�>'�Ӟ��I�#��땔Y�]�hx�ާ�u72�ĸ��e����͛7o޼y��͛7o޼y���>��_��>x�X�6��M!��]��ƚ�.ߤ��+���q��s���Gt�u|'/��P�%�YF�#C���5�r�|3z�A�Od��Mή�`��q�Q�q��wɗ���>���`t��h�%����ޗ���ݺ�hq��J�eBk��?����s�=��n��n�`���/����/����kO>=4�B�:LR�K֋|jNM�s�7����*N��>�S?�����D9]_��-�=o��ȓO�)�5�����>9.���G.��J ��l_ʋ'��]C)� ����CZ9�C�&	m�����<y�G���<�zZ����֤�f��\�����~�m��x
�Gi�$R��z|��P�䉀p��ۨ|�N�/�)Ow�&<�f���a�0OMN�l''�|�gq��rymK�1�_���lV�U���O��^!-�M��돉�	�,�ߞ���	�/��L�L�M��?,i�V�=q����^� r����z��7���9�W��;�۽������?3mqmw�os#«NS�[��|�͟��_��j��*eD��J�!�4�O��6����՚|f�lm��gQٞ����]����Cq:ޖqsr���y�Ծ&e��\�[Y�̃<�g/iXG�	21̑�s����A����͊j%O�Bh2Lk�f���?�h/�~�1�0R��xڪq�����~Ht���)�k7oYǣ&�_X�t� B�M_�R>,ǿ&�m�_���' MI�7�=��>4jTq�q$\���Aە���y瑺?LI��̞�H�D��Mbr���'��X AHrR���^iWW/��zϽ��ܐ���==O��D	��$�p����jW�8��l�K��f�y����Y�7�db׽�"�ン�]G���s�+�$+�n�&[���gU~x6�8h�P����\����J����V\r�;�8��q���9��)��矉��]#Қ�ꌎ�J,��($�����Z^5��Z���k�Ԋ�}�n�ۦ�>o޼y��͛7o޼y��͛7o��+f�y4�7���s~k+B��ݰݑ�ē�����S�>��sqZ.�Ǳ�"�(��Iz`��8]�$��^]�Int�u���F츶K<�wH�ey�}����6K<T�O� �F����h����-�pN�e�Ͽ�B-�������p- ��(j&�lO͒Ƙhj<��hh�6�4��MB��ч��1������ښ��:�r�6�ՠ5r��d?���x��i�j����߯_�f���Z�-5c֖�p^��A24ƕ6��>���2j0�}�u�y�m��:����՚3nmk3���4qt��]�C��,��眵����R�_��Cnx��wʺ�̂�/�݌��gy��,���3�'����E���Q+{Ԑтr�A���hO�P-����E�z�������%B$*H,B ��@���7��E��d�ؗ��AXk3�[,䶳�![S_��)ɧ��^����C�/�x�3ڛ�,t��J+:�j�Q�����2o���ɝR�&�5�h�$r{;�|�&���CBS�,���� ��waA�O��LY];69@b7
��$$*�o�]�t��w�W�G�< i2:`s����tZ��GUS���5z�D���| ��"/��71���'8_����jlv:���J��CK��>Aίc�h�/�k�A"���p��_�k'�����RIEoOi����y~�!�o7��&�Xa4M�n�x�㙃���!ϵ����(4�rs��]o��鋑Xv6%�:�*5~o@���{�!��wg��:�{���f�b:��j���y5JV��;���h�/��q��y�h翭��㽞���݇ ��~���,w�8!�QM��*{�5�AK�r匚�(y�4�k�Hm��U����X֊2�}޼y��͛7o޼y��͛7o޼�V� @�7��+� �s$��6VE+�^��(OƯ�گ��'N�i!��Y��T��#���E��Ū�*�Ab�����جhrJJo�f�8��ܫ�whnMCI��@XBO{>��:I�Sh�ĳ���O��&���<�C����u�Ά�>k���ʳ�hy�Z��~rJ�Է.K��F]~�����xNW7�#v���<F��D �+/	��Q�A�5���z#N�y�9������xd�yL��pC���vz���8��$}�4��d��i�~z���:)�X-ܯq���DפF���޿Hy�Z[��8`�:�3�Q�"��� ��F�	(�)��My;��hn�ϴ;�bB�2��Ў�r~ɉ��p��:Ɠdꡭi�ss�t�~�v6�pxT��-] ��8�'�Qh�Պ���/�h���CC���Ftytmh�%B$@�Xom������&E4��&S[��hɌ�\!�~�R��G��C4�3$�yٳ�m��#0�7
�}�~MP8�����e\�ݎ.�jo��6z����B��訋���Cm�Q��٩M"7�m���k� �H6�H֢�&Qڸ}��o$`�M���I���!J}�8�����ڟno���h�g�=����u�\�M>�Ֆ�0�!�0OȃE�`��̟��wY��٥I>u�i"���>;Ϋ�ӭ��5ޛ�]�92d�3=�$�v�A�$R�Tkl���f���蛩|��ġ�L�_������ɸ&��@p.�ߌ�j	�}F����b�LV܀���xHb�&tR��o�g�i�5/4	ل�!�B[Kp	���wD�3'�P��'�����Ӓ��۫�'���zޥ��9�����oM+d��q>����U�fdJ��'���o�Q��[����9�C�5�G�����ѝV�h������vI]>G�c���'��y��͛7o޼y��͛7o޼y����ϼ_T�G���`o�A��v[������/���8�!* �F�a��_jT4��H���BE����p�ʯ�Ei�0�?N�0#�bw�;���W���G�Q'Y`&���P���0�E}JE��wj�Q�*"�z��.ZpԪ���D�ڵ+ =�����g�+D������O�⅟z)NK ��Ή��D�U��g�E`��I>O�,쵥��I�ٿ_�EJ��}�8}�3������"��y��ՠ�w����!�6v��8]�&�>D�~�j�v�r�$�<������v�����ŃZG�p蠜�͓?��NO�{���Q<��ĩM�iMIZ&�����g'�i�}�''�n��K�o��P{�)�]�Z��H�t���!@�G��f4�p�=��\��%E����LJa{�xƴ�i����H��3�}�������x=3��sK��v��'YG��&?鱜�#��<�$����ݔ~����(��!����l�[�;���X��&G��XP����%L2L�>�{������d� ����$�%���hǍ��ij�w�Q*�?v?��F--�K֎���᩟m�*H��n/�'���N$�@�6��2�wH�OD%�5����A�
��!�gߋ�g_xR�����Xd]?��خǠ-�}wD�{���O
6@'Y��ܐ�l�Ϫ_W��Vj|�]}5�G�I:�?y�A/ynr��Bp�&�nO��*��ڈh�&S�'��Ժ��$�f�Es�)���Y���
�6� f����Gb/�ԊV~�(����~��;�;���b���2�U���LO�||bVV�T���4�Σ>�|u�Mr��<�����&rѥ4��q�f��H�7����\�b򇕑�v��㲌����g���C����sjϱު~�1���y2	�T���mU�"B3�/i���]���~D#N�<��͛7o޼y��͛7o޼y����}`#���{C2�t�����S��O��?!�
H�������l��X�㭬��Y�cA�2޴:�#%6s�c�;�,��8ȃD�o��K}��Ȟ�n�c��$+2��s�^'��֥�ho��ix��b�:��W�����Ot��h�=�Z��']^����ġ��b/�(�����r`{�ǅ�y��U�~vJ���ׅ�Y]_��4,F�����^�1�	�"<���==%��bW�o.
�w��q����������Y�\��SjH��Ή��^�@�l�@�t�B�V*��
�yَ�@F�	�7!DqYLy��v�xT��O�����Q������l��� �OIX���;��fQ�qH���SS�:���7�nw���gF<�xF���D{����kBp��5�?V�8��XoѮ���8�xN���B����x����qZ�缹%���������qz��;r9 ӦA��x��8�r�r�^�!ѣ��&��+`����L���G���W�I{lV��}3v�8�s��6r|삘��(�D�BW��zs�C?�����N	BZ��4����G�Ֆ�F��������ـ1 R���O���-k�F;%ٕՐ��}'�S��5�1"A3��8/���ϷM�eE���2=ж0+*mjΛ�Q�z��<���[Ш.��Y�H�.C���D��.��AI+�ݮ4PP�T�lP�M��Hc����q|��O���s>7%)�`����n�-�ï#˜�{�TF����s>E��`�n��&Q?1��7�*��"\�'D�o���{�њE�j�-�}!�}��r��K�7�t*Gz S�	������`7W0�1�q2� A[�q|fZV�ܼ~6N''d~��
���w�WF[��+24��&9SW���;����K�'!�0�@�X332�_Y\��=3�b�_�E9ކ��C���˳VP�m�Fc�o�p]�s�!�t;��Q�>ہj?��%��v9�2���u�R���
���~ds=G����x� ��Ļ�N��Þ�is�gW?�:�m;�ةs;��vX~��&��t{ŷ)�q��{�ϛ7o޼y��͛7o޼y��͛���̋�ȕ�4^$����a�.Q5?�����h �`�D����r�~�])��m��9�f{�:4�TכSCD�����h;p3��.[��62�4j�F$�(�4�Y�$�w�r-�@ꕘ���=ɰ��g{���zmNG�z�hϊx�
�P�&��v��zP���	!�EtmiǥH!<��BѓM�3z�4�3�#Ϸ�OO<#�'�#��|��h�,o		؇TH�.�,�.X�N<Ӓ�'��������BS�d�q���Q�!ql��g��vS<�{������h�^�"~m�]����_SўR�K�2��iDO\Zg����n{۵���G��3�����֚(	�vT��+��+ʫZ���О�v��}B��e��A4bI����A^���ѾL4Y�S��H;���A;*�<)@K4I}�"������g��b\탰���$a[��u��+I���5�E5y�E>�ڳ��:��:�3n��e{�G�ｳ�f�n]`&
�qz�A�h��)M�Q-���aG��}w�C[���H���@ju�yJ�r\� I8`{�f&����`+z�~�5�7Ve�����02+ ��~'�Q�1\)A�Oi��9�2��G��囜E6h�@�w$M��S�K�����ѵ�<F﯆7g;����7ڲ�mRP9�{��U�h�|��?����'�J6ÑE��x���B���1�l��'�������B3.�Pԧ�$I�>�k�܎�������-���:�`�h�6	����]�{	����|j8�c�̼$P���@=��~[�ۆ�B~z�2�?�O���_�)+i�M)���O�l����mnY�q����i�� P��d��{��V�sx���~3���.C�aY�j�d�W�72)�:n��sF��Z���.��?���>�Ռ������p�MO�y��͛7o޼y��͛7o޼y�vXf�]C�� o7�ѵ՗7�{J4�3�Sq��P�t�H:Ak��͖��p�J�^�)�I�
��|���8�M��Mn�zs+�@]�]`fF2��j�}���yTCf��X�h�/PJ�r+������� �ń�$����1��9<.QJ���)V�$z����<>��&a�Ֆvq��8-W���-$]Q�eg�H�}5�JݾY�>�8<�5��T����&�]}D�-J=��	�z���D�Ϻݐ��`?�|橭HR�������� �W�+�3���O< �r��{CkH`x�Y{��t}IN^�������LW�`��	H�K������l����M�	�!�?;�ՈbmQ��{$*��9ф�mK�1����h����}�m���w@Ƨu�H�ءӱ	OCh��@R�d��K-
m��`�_f�0���aԾRَ�g�Bs���q(nF�H�sIr��R1t�VϤ�D�g���4ůCŔD#��qڔ׈Qh�s�ȴ�� R�ΐ=o�������0'���v�N���������Qx�ډ��*�a���d�K@�ZW�oj�m�w���R��nM]M�D�ݿe��v��^QY�4���o��"������l��A_E���ph��]kx�"�눮�����~�d�w��wؿ��)b�r���8�&Z�h�.A�	�Fv�:�Y���oH�r�H>��zú�m�<�[����$�&ʯ"
�r3Lp�yE�jB3y�A?�yn�+��Q��g�lQ�_���I�O�z��Ԝ�&bN�3�+L�����Fe��&@�&��(��\QI���!���?U��ΪԿ�s�B(?�r�8�~�4��6��<�R�Fuj�Y>ϕC����w��8��F�MgO=�&�j8��fٝF}O������T��{{r���zWy�����`4N�<���3�};���y�ϛ7o޼y��͛7o޼y��͛���R/��{Bj�� �H���f��*���M����������+�ZJ}�¼|��������vY���ÿN{�It��P��8-J��3q�Q�9�Hy�I���7��e}A�&G�G���h�FLZ��ށ�6�~��%D�n���Zؐz]���!X�7Q<�=FB,tyN2꽉J�v��,�++�n�&z.
�"�M͖͠$d4����-��J�Ǚ}�B��Z#W�L�;=��[Eh��A8���q��YD]�F	����J��g��6�>��o2�hf)�F��MAZ���woL;��=��M�t�� �e��,P�̌�M�q�%����sq��.Q#�@s�dZ�hk�]�¨�B�R/_���m��3r�x�����&{6Qf�tR�E�+ƳI�tZ��D�h_c��G�̡�Fb$a}0�rU�\�����V$PHȐ�"��C�@j|1Z������RQ� ꨦ�!|Q�	��:�:S��Ӗ�P*�Գ5wL�C��W���]3ED�E�wu\]^�~�A$�@(GCMy��x����RB�g�'=�,�$�&�F�d��ݿ���������U�<�`����w�����������_x�����#J�M���E�iyE��7�`kS�s���~H�I;�ki>�q�]����2���GK2nl�\'PG���{�'K����e��^���{7�@ @���(�"�)qdS���혈���r�3#�&���iB�F9�P� [��^�k�z��V��~O�=�n��n�n��C��W�ܼy������k�N��3���J'"%��X���~���'a�	(W+9Ӗ��ױ_���&��9ϣ��Z���r��xu��4}�	��z��5�/鸏:V�<z��4}���4�2�4�RF�/WI��t�:[��s�*�;uR��VK���iO;8Z�X\���ۓ"]D��6@�[���wk�jl�>�.���׳��H��ަ�X/8���>�5)�&�o\��J<�?-�>1Z�%���I�|r���P�;L�~��v<����H��gD�/)|�$R-�g�^3r�݋��vTT���aV�zy�kI2�����u<���/X�`��,X�`��,X���*�O���D�ѺF�:dTw:��X=&�zK<<o^���IDED���x�v���ꎐw��1��AËQ1��dF��Du�m��ˉ��J��`?��<�[q�e�=��I��F��zTK&_�ϯ$XNK�ȍ����y.����z5��Og(��p�F�?~��c��WM�S����#~�u�FF� ��Ӄ�84`v���u��Ӵۆ����G�0j�X�D�Iu��%��v�#�z��ߡ�`����K$����򧿐���/W~���܇�
��4UTce��O�<	�3w�����5��%�kGv>?f[���������߼-5;�R~�!��9(�垟�4IUh�!�C�v�Ԅ���\_w3껟���T���ƒߛ�V��#~�zg�V_j��e<�2�G��}!���/O�]k)V:���Yo!��+����ci�G�@c84Q<D�o�)��F�El r1+gI���7v�e>��D�~}�$��Ũ�uTL	_j���Xr�s���X��f�|7��+D���ɗ��%�y��f]����s˴��|fQ:]⽔��оa ��s���p��j�z��1i���R��-.��Cŷn��At�n�ⓑ�DÒ"6ڥ�G1�b�(��y6���'�rD��~9�M&Rɘd�YA�c'ety�@�6.�5E�hH	&�Ԝ�#j%J��l�
�~_��4h�ߗP��$�_	v괼��I[^�y�h �붥�DF˯\1�$C1��=��/�hc3�Z^�뭞<����9hݢ|GcD�1��=���~����^�f%�sd�!��~���_0㉩ל/L�r��cH�77�}��r�J����h�/ZA1����8#_���
��<��+�_}� `2=��ŎS���=Ic.�L�]�W�1�U�w�ͦ�|���_�Z ��,X�`��,X�`��{��C�8q�KM����wGP@&����k����m��49�!u[[]!8���1V�瘚��(�aV?�/�>���u��z�y��&������a0O�d�f�߳���,�ߨI�#a�0�^���E�o҂�D$��1�\�!���>jO$��)��q��vE�9'���z{�}�8��5Q�rZ�􈺤=��w��S�����П0��u�u��^���o��o��5� �눇����go��|��5s�5j��_Ȣ��~�ghb����֬F��%<��V�y�����-)��x����;{BP����f����nWbH����H�m��1��x�iv��g�Y�����hS���V�V��Ĩ����(��6�G�S-�������� �;F����j����`�nK=o.���.D���6օ���=�z$]��jfOα�b"�~�ɹR�y��<��_������#9��A�Vq�<$���Î�wH;*�0�Ɵ�����ӵ�m���P6*l�0�}�M|J٬�z�i����%!���� blZf; ~Jcj�螐�B��ql\@\0��ܙZ�悕0�GCw���<�d2Jr9��1o�T�������db��-#�*E��PB���� ��5�/��1��o槃!]�獡�m���G<�Ҋ�Y�~<� ���}\oLB�����$
c��WO����p]jb��u���>���K�"�=w��^�ĐyO�V��=íp�������i8_hV��k�e^Hm�25%V�|ؖ���K��5��y��ޒ;�!�a������)��n�{��;M���x�;^���F����v�q��,}��,X�`��,X�`��=V��ob�,�[�(b*.���j�xr��B��:B��c2ħ�	�:Ώ�q�X��詡G<�P�I�?�J���G;l��*_Ӌ�����*���J�bym���D������Bϟ%�P��E �;�mfx"��y2��`O�/
�z4�Q;Gp1�!:6���-�V&J,���יi��zA�FLZ��|���iK���N�~�ӟOӲ!�;�H��=#�0|.á�J��l�!E�K�iTa���W��Wt�\NJ��P�������K>������Ġ�� ��|���d[���4I�AB!v5�����<��戱�I�ޕ|�qi���YGR�$�Ֆ�7F����������wKرt�1�"��!H;�,x$i$tI굡�ٚ�b�ZJ59MNj71�6�3�Gl5�,�go?Gf��{Z����Ԗ�AJ�����/����������o��rV��d�Fg���������n�����f���=W.&�؏̦��z�݅!r����L���{�e�iX3>�b��>��l�a�p���Ro�m�ޓ�F� zj��3C���y�#˓�IF��F�������}+urQ����g��y"�kd�+�(���6�cch���!�� �UL�⌐:����w��ޓ�j��$K��Ip-�a㎬��⏚��=�(��������ZbK����8_=���'d�����L�����MZ�}8�DϏ���VC���̥�q�b�[�c>�k߬�{����<�^,ϕϭL�+�&�f��5��}��;�(�̆��y�[���?$����lv�r��Ȝ[P�h��5��?s��������8!�vdR���8�?`D�X ��,X�`��,X�`��{���/�d���:�b�y�'X��h���*5��Ӆ+�$�*p���=|$��G�Ol�%ׇ���?��E6�1,:�tlf;�s��ԒS��c�uu����f��xHs�f��e,���D��e�s���6��$�H&�\�G7r]5
��b��S\���ۊ]�B�/$�:�MPHz�s嚋Rd	��_Ί5��y�,ϊ�x���4������׆65�nݒ��w��NSF��܇ǚ֚m�F1��Z5�@�KZXbab5o�T�_�/.8�Ѭ�q����W���4}�Ӵ�z��?N�?���Ҵ1/��+�{��#��h0J��5 Up�
��b��nwcC����<WF�=yB<�sB�1�rQY��W2��U����<�q�^������9����G- �~4���%J���Ʋl[m@�Ԭ�yzx$�T3U����Aҍ�&�w�H^��]��F$E���P�;bz��#�����?�o���Zo����.ݛE�~f����PD����n���[�K��zCrZ�{4�������F-E�O��g2�f�]G��o)�|<���t����%=�Ԭ6�/�^-��-G?��?L�6M���6����<D��Y�����՚Ӧ�|H5�\���;�a��M�q�7�9�rN[׌��9�R�~�9�X�|���_��	�0Es���htYh>'��p�����	��+bHN�}q%�ծ5�_�?��xlW�|�ּ�[6^�GW+2��1s�~����'OKtݍ�m���� ����j��٨��s��v?������M}���A���X�Ä�َсU�	ad���8�j ���^<�M�T+eL�=�m6}�}o��9�e�m�q�F]�>䋽�}��f�~�谣j��8��{���}��]��Z ��,X�`��,X�`��{L?��>$���C�<F*A�f8fT>W� !��/��><o��1��d��ϸN,��q@Z��ClQ�K�T��3|W8U�a��~Q���������;,�*O��"^:xۛ��y�O�&�iԀ��#*,oTa}��t�"�,��z��w�KQm���d�CKbZ-�a�;B�'� GԦ�x��:v\O�z0)�Y�?T�԰����{;�'�4��]��`O����$j�ȅ�;�"f�b�j�9�9.r����1�`�������٭�+�������O|"M�5�;��n��j�� �Ir&wَ��u�Bs(�ǘ�L�O�+׮�|��U\T5���-F��F�c~]	������ZyԐ��\"`~Y�˅dE�E�:8��ը� 
��p52�׶K�7�G���(���(�V8"��jJ��m��8�&JN�H�����xtI�,��� 8�o=��Z����w;\�rԔ�i}� _���T��|���Ղ�O����w�uR@��o��Fr&6؇�Q�S�_~�����#I���y�~��9��N�qnʕ4�0W	����X!��W�&M��������G���-�wowǽ1�����ڄ$�HT��]9b+�B�_4Kg�v�<ї�XI
2�l�F3BG���"�:�Lu��'.�饷���{81V8a���Ϥ�s}A�7/�w�%+
޿-�����a�����Gn��i�J>�s2��ߖ�/����d{��77�Y4����z|<};�,�)˳�@אT@�q�\��\@��eٯ,幾&�%�P�ֽ1�VY�f\�����a9��rv��f[}%���!xǹ���S/|D˵�7�Kf�%k�v:'[��<�N�'��i��znN�w�����V�1wU�g�sߗ,1�+�����'����:��I�$�^?t�1��������_��ݞqސ�L�=j��rϦ��������@�,X�`��,X�`���X�F��n~���!��3
Ϡ�(x�MO�D]r8�$��.٠a�4?.����}����k<}G^��'<�擯~�.��g�J �v��YX�eoO<+��q�i�Iq/�ikYB`z�&��˵{%���\�7x�y-�F	�G��d�`�<��=k��Pa�҂5�c�����b�<.��窘�#���%I�N1���������%�&��S�	�`i -2�Q+'e�J"����׃[O��{��yf������jQ���n2	Wk�'���4 �$Z�_\G}E��s����A�֤/�y�e!_��i��_�j�6��O�!�ۛҿ��}���-��IDm��s/���?z�U�/��\�ݚ�}<��d��Z��D*�0�6@� DH�5I�1/�䒹�w���f�^�WvɵjՍlk����%!!� u*$�-�7�~�?�4�s�ڐ���?7�1�;��=�o������LL�XN>�Gf�R��]�0�4ʻ=�������2�y�}V�M畜���h�<A�D�K&�ʉ��2�����m�Vb������w�֒��{_�/��F���=7��	n�K�w��!5D�]!ź���J;teFu�q�K�<�5���G�	=DF�?u��|�7��~��{�y�������{=M/>�D��?-��DE�A�c�A����#"齿��������ɢ�RS�`�-7���9pƐ�^-�ȓ��_��$�[��\� �F�CXZm������<9����j�����Ҍl<���վ��#�g�\ ,��]jS�����mi��wȗ^�i�_�Θ$b���7���y3�o��|�s��!��%�
�.��f��/G�z5|�m�cv�]�6g��&���{���,�sݴ�=������a�<�j��%�>M�A�q�?����/X�`��,X�`��,X���
?��?���
���eUFT�!������3�&�S3B�����������M�P����Q׼���%7����9\=8��LD�xD2"BP��9����\,.0���V����x)ђ�@��P��r�q�ⴤ5r�DH�1F�P{_<��yj�Ѓ�#��E�����yB]�,Z�y&�@��%2@�x�&�'D���a�����Ĭ�ߢ�Ϥ��lD�4t�'-�dKH*qa4T,�j=�L�g~b�L��H|�l�r}s�n4Z8�z������f� ��z�4��_�z��Z�/��izkMH��M_�W.<!Q�>��ϥ���7�������_Jӯ�ʯ�]V$#��<�w�z#Mˈ�K2H=o��w��H	�2RJ��W�� &�.1�$oA4O>︀@��YJ��,ڢ\oeUl%�Џ�fό윒��o�\���v�Ԥ�a����ۛ[i��;��<�}�6���t���C����Q1;�h}�V��7C<:��'Ԫ���(G�� &�-[İ�o�.��q�ZY���!�f4K�(��yq��<C�!��	�-v\�j�'��1�`�\2瀜N�5f�mv������˲=����X�B:�>R���0���� >��+�? �9���������א��9�ˤ�?���[������r�1/d��h�?yJ~�7r>.I���6�3ⶳXI���<�o��ުZ�V�X	POr�T�#v�99q�Kt��Q�q�+1jC�V+���x���|�>�g�o �^��n�vm��\43V�fw�Cn�22 �l�P�OǑ�\��mV��6�q�+3�^v�	��
xT�a�>���|�C�O��7�jV�����I����&���,X�`��,X�`��,�C`�}���D�>ʗ|z������ Qi��HR���')���ܾ_���YO�}YV�P�����|,��k].���C��ԣ���������f<�6?G��wT2L����@���6�A	�3�/�� *������;I!��0`�U'F��ѹ&���C���L!�S��d�Ϧ#]�k�[��#�Y�H�mYO����X����9>#�&ĕÒ�|N���bx����m��j����\��ɾ�vB��$��>��l#_���D��w��i:��paa)M����L�O~\4��\�����_�F�6��%�4<�o��(Wb�;�����N���\A�Ș���m��ٸ,ۣ�����(Q#߿|9M��Z����U��/������$�ճ��m����5���Q�7���Zk�WK����{{Α��$m��7��q���W4��_X��iO.Wٴ�Gɺ��{:ޗf�����)����de4=U2��I$�Um-5�tW��qy�d�{}S���ݒ�j���u��8]30��t�z��H�b��IЗH�a�F�< �QC��s9=�IɴC`�!�.՚��DF6��r,���{WdHy�iEƋc'd%@��ڲe��$�Ɠ�8��&����ͯ��3��|��tb;�*��������\�Y�CS���iF����!$vI�z�4-�g�s�$挖�>N��%�>Y�1l�}M�~�{N�оW������y{5=v8��ó�}�߽�#�d����_|�f�����"(K2��u���g ��,X�`��,X�`��{l�}�v�C-@}D٥g���K� :�$��2Y�O�l_z��E�pZ(ف�I����m�nE���D�O�/j�ѣV.S����:<#�I<�"�g��S+�ռ��rK��}&2�<:����*�X����I]��v��j�D��5Q�&j5�23�7<���\��-ԍ�Y�'�W�
��O�;1L9���^N5O���RU׎��Lk��|Z��%�r�7�<�B-&�A�wmO<=��M� @.c��[�Y?�wոI"�����!u��N-��+�]I�ǟ�����eю[9&����7�~+M_���Ӵ5'���w�:Mϝ-��~�y������ �Qv���-۪�Wc{��)�~�mHF���6z��V��"1o��?˿����Ԡ�ʁĭK^�9���}��m4平�0�<���x����B-jWG&��a�cd�g7�?�0�ӣ;��LȎx�I�|�iP�h��,�~��f��2�����s��i���9��ٯP�Փ�#�l��hy�r�7��5�b��W9	hV�h��gΓ��a4�����W}�lo�W�s�ю����?���|���9��Gu�(�w�g�#	� 3������iz��9ٽ/�-��/�y�tZ۸����D	�օ�� �89�8�䫳'��C̛� �� ��Mٮbܭ7e�_Xm�f]�c9�롕8,x~{��5��d���+}Ltq�Xbl����-�E�,�Ce�>]C��^9�Ζ�8�s��ښ�s�(�2'nn�`W2�*Fd�����Q&���'��s{h,����'B^��y-N'�S��h<�|���^�|��`��,X�`��,X�`���C_b<�*=���OF���M��|Z9r2}{��W���[3}dbLq.��_�ͣT�ƽb����1f_�A�1��z�\�D��S�ʓ݉+q/sWʊOp�Sk=��Κ��9l1�����5�0b,�!ʩ��f��p�O�(�����:esb�0<$�8Ghz�9���+�3��+Vr����ГԲ�a����m�R�}ZO���{�z�Y��`���A�B��<�C�"�bbɸ~"��م$!��MAB֡9Wc>|�6ˣ�엘|�AV2��k$��e��Y^��
ͻӧ��{��������r�����?�V�s/<�d��@�^�J��(z�H4�hά/�*�-3ڡ%�,yw��&%Cl4��㍫�)���Z�F_�������"��3ד~Ֆ�ꉓi��{���}�umo�n
Γm��3���|����p��%L�5����g>-�Y�W����nTu����_�`��N�(b�	ml�Q��/�k����h�r��q��v��푰1�:�3f~�q��fO�\f����Vk�7����k5j5('�ޗj$�1�r����9���_S��GSO�=��?��_L�g�}6M��O�4M���ߥi�� %�8/�i;X���?��4}�����'_y%M����gi�����n��w���4}�M��]B4]j��0��A����8W��8q�D�K�i,?�|+#��v�]Y����>B)1�q�_l3�j��$�l%��^�M_�_L\��þ��sE{ ѷ	Ҵ�Ӳ��hF�	V.A{����ZˈB�y2?��I��gd�Q	|}As�4kw��3�ӵY�I>��FK��<�?��������ʈ^7�n��}��,X�`��,X�`�����f��7��'��/����§f��cQ��C$ ɐؐK$��Zhe���~�|�/�GU��l�����m�桳�$�x:F��HϞ��砞^�*0_��(���P��i�u��B1�hB�j/��%�7��}�w=�ER7FE=&�h=}���&��v�v�1���^�_��(W��jSe$�u���|J`j:�}�}e ��9���B�6[�k�y�˳��9��x�+�O�Ȕ��jtЯGK� %Z�l.�.����O;��NI�7���2�i5)PNc��Mh��,`�j��atӨ�!��y;��N~�S:����m�3{��9���~����+���4��_'8����J.��|s���ۻ;;���@��PPs�[�H�Q��Z}��U������a]�>�f�{�zm=��{qq1Mwww���>�o��Q���!�;�����B�5��&�������eVp�E�'��|�eߌ�V�������d��3[��4�&�٩���1[��L�C�wI�L�+B����>��Ӕ�a�z]!�]�	�e�2Ii�M��vR��Q��]���ٶQwK��#Ss��~�M����sO���rՒ���V��FrQ;)�YTDWT��<ϰ/ϳ�q�Ċh�>v�4�a����N�nnm:�/.y���)M?��'����i��_��4�|��4��_�E�R�����\��7��������?�)�cU��Ư3-\�K��ꎷc�\V'K�j	x�s���2��%;�ͥ*��jx�<L�צ!��~�F?�ML��4� �[��0k�&	WҸ�g*�����[�ʉ>�)w1�s>��g��gq��>/���qY0�ֳ^�ޯ�G�6�[�|�4x$�i���c�s-[a��$j����M���3<(;�4���-�WΪm�*j�u�`21�8N����S9���uJG�@�,X�`��,X�`���X�>E�j+Y��h��G��@�����:f��~a���A��z�1լ6I�}$���Y-�h�d*W��^X�w��s����F�ǇњI݄f�՟���'ΟO�'�n�u��Fȸ����v��D{�M!�F�x�=�����f���z�iN�����hXc���W�i�ޛRn��V$]��N"	��j |5t�JThƱ\��]�F�4��he�s��#LS��h�XϾF��j��$���h6eZ�=D��#:�u�Eӷ��>���L܌���C'�Z���a���u_��h����)�]{S<�e���8����p}9��%�����?��b\b�ޫ7���\Z�z���%�*���ϽF�8,�����FM&��|�6���:�X���j*V��g������|艷��l/�;;nv<�Ѩ��*͕��7Lm������㻝�ԫ�ZB��;��YL�s;����n�^Ԃ?$Oz��y^�mL�_ilA����X��+;�Q6���E�dtȨBδ�f�>޲�D�w�8�ճ���� XbȼL��HS����L����+A��D�cT�Z�Q1y���������_��.�M�'�a������^aI���v�bJ��t�%�u�U���+�� W��3�g6�>V�,.���AJ�a|lb���)$_��t�ow[~����4����_)��o}3M���8M��
1H��~��4}��~.M�~�i9ߚ�ڕ�y���2��9�_>E�3Ώ-I��-W��Ts�	W�Ȣ/y���VMi�ǚzhV������S�쎹������h�reQl��}Z�IN�o�|���3+fX?�\w�e�bWV�|�L��j���=���q�g}ʮk�����6����e�WNt0O���{XQ��W��
G��~-AiVF����k����vg&�rZ��z2k���-����ߡ��Lo�9�7�R��ɟm�3�ۚ����`��,X�`��,X�`�;�C��cmz4����Z��H 2���b�ӑz��O���0|�I-�߭�E��N,��=�l�E��d]�����ŧ�ƨn�f�&��I��k����dr�(��^dTy"�y��B�%�}���iz���ٜ�N�X`�j�����=�ގx^�Њ����DK�w�����/|�iڨ
�Ҁ6���jxY���n�|40�>���������)	���xf?�˿��ux��ʒ/�|c<�\�7�Ѳ��P���j��6z��>����}z�����F(S6��c�o�DΧ� �G�\V��F���y�����ڔhb����4D؏�!�:&�B���z�A=X��vT�'1�I�W���m&T�2Pdz�C��'/��+O� �^H��ߐ���'�	�ﭟH��E��m!y7�i� Q���"�����;.d�\k�)�e�%��B{�>7��h$WvIe��ֆ�؞u�#9�/��?�j�V*Ԭe�6�zU�j��W��[~X�ygKʏD\��d�0���4�c�2=Z���@vm�_�-O}U��_v���Hao���ٷ�Y�?�mZ��d��-���W�ߋ<�lױۮ�����?I\By3r�Y�4#R����ژF�3;��W�;�Xm@>o�Ch=q>�B�_j7YMK��M���6X�G~�iC�q$���s|.ʭ]b�6k<d�����ש�_��Y�Zw��s�HZf���3nB+������>����V�/2$��.���!��6(B�f6[�Q����4z�!��I[�x����R�۫Kd��op��@S�Q�IF�-�;�o��z{���~���xjL����>�9��[�\O��Pƛ?��?I�c'�� 9����4���E�B�p]��Z�����IR���p	�Hs�OՒ�y8J\��H��W�G9��`��̟+UŸ��;s�P,����[�"�;z]y��/����Ҵ�my�X�>��ry7������ �s��}1�G{D��_�I�ݾ)�A�;2?���O�4ɛ�'��o�u#j.��s���G�������qG��{o_Jӏ��?�}䯉�8_Y>~�G��N��=�6x������/��S�S���`Q��⬃yU����
ʡӕv�y��ώо������kӉ��^�=�Χ��7�%�|��|�l.?3ڬ�'���'�vȝ���/���;�;��q���]&2�E��`��,X�`��,X�`�+��7�D��3ڎAZ��Q=f�=�kR�i�ñ�|���xR:��z[��S�g��)����sg;+'z,�(U>���r�=�>����/}1M������ŋiʨKKKBu���1"����K������o��%M�B�ғ��>���O�IӓgO���杻/�$��h)I���Z(�����H�t�Aq�!�n�'��E��/��O����)�������r_�B�I��f=�Ԉ q�n����a�vXo�%z0J�qZ.V%�����%�x��F�r�v�j�уƨuJ�����US��k�z\��
�i��Q}2,���"%��r�� ��^�w��l��4}��%� ��?��2��D���%�o=-|_��/��Ǟ�ogO<�kk�uY�K>揉���Z=M����?`H���|�AB�|'���#�>Ge���ŗ[������$'<�ܯ�(��xjIY���3ZDp��qDB�¨�.Q����{wg����!� 9iH$��>�հ4����Q��=�I,;.�ϖ�c~Mt��W�6�;���@K���"���ڽ�d��7���|�ڙ'28�g�m��%��i�۟eQp�y)�:����( ��'PS�
���d%ٔ܆�ݳ��ټh:�`�Ck����wƞq�<��̷x>��%A" 6\@���L��d�
�w ��j�Ԝ�<�D�j��Mj�<�6��*闸��n�c�ԛ~�iH\D��˵#w�}����U|�H�x�ͼfC�#�#ڬ^�[�����g<t����Z�ԫr�VS��9IO?�����~[�c
`���'Z{��[ߒ��ܔ��@4�0^���O��������O��A�q�C�/��@�/�,���r`�6?/�A�-F}f}�Qo�)����ߤ�s/K��/}�+i�v[�##��M矹��X�;�7��|!�9D��uc-M7n	=�y�SR.�X�QdM�0`�W���l��<�Ҏ�ۻ2�����_'M;�d~������!��!��X�y�DW$����O��̹�i�C]��!h90�}�P3 ��$9vSB��]9c��ʳZrW�0
4+��Y\QB-Y���R�Y?��K�6�gC�e+�r�mQ.v�c9a\Օj�"�Ղ�&n;`;ҕd#�����w�6�y������g-��d�U���Ĝ_���/X�`��,X�`��,X���
?�嵶�1�����' 2%���;r�Y�)(݋��h��hB8Lrd=P>�ݶk�2�C�'�w��_�c��{6�3w:%dƉx,�Ec��_�Z�޹.��4��B����U<"y"�h����.-	����D}��ci��;Bƭ���"<]{m�d�F��#t�!�z &c]�?5_,`F�����7�tC�YN?���鳏J>��B���FI2�z%e�4�G\65J��fd�?CGb���ݒx�"�ǉf=ZU�j��i��~���~M�$5n��2<���8�z�(�1K(�@O�!��<���ݩ��G�����q�{�x�wGBhTHL*������h�A���i!\Ϝ��7�!�}#<�^G<�$I�6����N��r�q���$hC�J�jT9�o�s�D�0	=j<�����$ϙ�H	�o��{����LS.���X�s#U���x��O��@JT�n�L�kz�T���$�z^�݇'U���.���S{	$
5sQ�5�KH�A���%����0N��2�Y�S�p?\�Ϛ��Zd�^."���ߏ�~��'�I�e���t��<ڇu��c<׆j�B���[hg�R���TI��}A$�Fю��V����ɫml��Vlt�� ��y-C��jRU�K�����%lKE���s�N$J@�U� 8�(���-잏Z��Э_=`��V��ڞ��W"D5���`�!wM�z����d�Yqa��b�I���h��ȭy�Ԍ��h�����f��Гy�#�<��gN�N��^]�[�Z���c�P�������[����v��u�ҾN�����WEs�D������oʼ���_Iӿ��_�]<�G��ʓP�:�	���}������B�(G�[��" ��|�rlD��5!�N���Ȱ�7�~VO��q^��/h���P��Ԣ#A�v��u�}B���e�6\h���7v����&�s��0W����H@����t�|;����GeEPm�Gn�.
y��/��Q�C<G�Ƽ���"Vh��J��P�񞵿'�.�3\���r���I��w��^[������l��F�0a���#��p�V�[�s�"�:&����(7�4�ʇ	4��>J5�i��pi�e������j~r��z=t�3��GBD=�q����tm���H�+�=��Y��[A�@�,X�`��,X�`�����D���BN҆ۆ�ʢ��U��\Kr�9�Y�����~2>�M
2��!S��D�)�b������W��{\�(�����fkk�A�u]<j�,����<e=h�Q�!�Q?����$i�41��>H�%h�U��-��3	3-vXd�����3ŨZ�-������O)I��5���d�8/������S�]��ܰ��(J�z�H&Y��?+���j�jU�SH"�QY��]��g��H!Z�ڍ�4S�m�X-��-���6G��wz�����n8�D�4�$��ϋ6��&ɶ.�R�F+ɂ����?��?N�'/JԸЎ������)�Ei��������?F{�vK��+.y�X�:��G���WҴB���H�0ڡ�48��w��,���#��G.���$$Bm4O�Y� q�n+�6u��﨧����{��"a=�FRtŧ!iڳ�8?����BLl��s��NQ!�&:��\�o8�I���lM�
��:i.��zX�D���0�j��[����M>$@��EjI�yD��M� ������l?$Oq�}���~X�Fd����e5y���+��a{�*�SoH�d���yl�]�h�������W�]�}���J����[���h��|�.��\�4�g��{}���7���O4��5w< �����h���m��"S���~�����|0Z��[�^�Q�>�_�<�چ�?��3�=I�&�3�+B�>J��W G��ʂR���t�@���G��l�_Q��7��}Y	2�Za$�^��Ki�����'��ec]V�<��h������4}�7�toK��������#�a<��pZ���{�#k�א���}�l�<wiU8��x�e��GpR�7�^��1�/`e�
��5H=�V]�����v��<,�\���x���A}{��ǜ�漽�-ob�b_��K~�<��:�><o�������FY��D���uY�A���,������HnC+�+�o�%�������a\%��b��G.Jy�Q��+o�B!��[�p��;���Q�� ���}��3��#�wV�5�L��=�]	E�Vz��6�+�|7`���e4��C���
���+�����/N{�iF��*��Qͣ�}��y����J�r�Ē���L��a6V/}��,X�`��,X�`��=���g�g�鱡6�������J��ze����?��J�ܳ&��~������h���jP=p:A���r���A|�acH��QS����������L���=Z>TG��y�(R&��"��5j��b��Ξx���{8�Y�*ѡ�Zc&���r�G�Y�oeOpM<J��P����d�~��ĳ��'����\A��sK��4^�K�гNbd��y<�<�Ǣ��ǉ�иG�Ǐo}x3�>I���£m=g�3�&�^i�iEj
�Yc>���R��}%��Ǫ(�I�,���1�loo��V=T9Aқ�o8��i��1���_�3<�(������%���^���s��xnIޝ<%�~l?���i߱�J���֥���Y�7�����X.DCd�	���8������}��e'�k�/�]7BI��H�Hzz-��j�b@yFh_�:\��+�v�?6��t�1I��\� K������ںs$V��t��%c��d��`J�����y�|V��Ϣ�8����S��:��L's�o��_���{5�h4jZfÃ�	���5\b�f5��* �H�D�PP��~%)�v>�,f>�(�5��ՔD��ԩդ~�;+�;�.�h�$��6�eE�*BR<���7�Դ��/��!Y��$���w�z�|��|���*��,خ�� �tm��JJ�a{�Q9[B\uF�^u��j12�:n^gcC���E�lwWƍ�Yi�zv�٧�t�~ygK�a��7m;x�ǡQ�~}�/	&��Á���چ; ���]���y�@s���ҳ�B�ՠ9[E4[v����i�X��s$�����/<�����h�ݾu�'���M��]��J��g�~Z�ssX��+'$�?�\�����˟��4��/|)M��ȼ��[��uA��1p���^���(�H-�j��A~=��� {m��X�A��ԟ�@�g�`y,�����=��o�%$��V%���O�8��O����h���z rWp��n��nݑ�A�����=���
-kr5m�$�[�`��`$��|����������H
K9l�J}�Z�~j�'���^���z�y'5'x������G����5Y�q���i��g>���wQ���Ic%���{�ԭ�����ޑ����"w����r��A˰V��҅Wcw�clVڕu��<���x�$�PGF#��I�䗝֕6��,�>��p\JJ�.�8j4�Uc���.��i �O,���7����Px饾���F�{���_,ɏq���t���x�)v?�Y2sb2b�E��,X�`��,X�`���!�)�\ϵ}��_ ���̗G�R�5�G#��������Gմ�oV�x�,�dS�%�E���~��~��h|�e~��G�_��%�CN��dװ�#�8��/�����F�e��z̨Z$�*��0J(�E��bT1j��I�����x�;sZ<���\w�x܎-���S/~B���$���7E����)Ҁ�tFj]�5�$�����2�jf(�f��\ԡ{DgHz��R��Dn93Z���9�I�f�%ٞw'��I&�FdE�h-nW�akQ�I����-!j�0�.5��@�L�(l������o{��ަF�uIN�!�h:	n�͌G� 6rZ*J4q�㞻�v����3���#�lk;É��!g����a�w�mL$V>���	��엤�} M����\���/��|C�Z	�t,��W�^܁V����׷��gi��_����h"m�H=��X�
��n�A*T���]�$K��'�Ȟ��/�-�@b�Ms�IN��!�΀�m�������l����g/?)����'v/ӃN�4�����S��`t��v�+^�d��X�J�� A�����Ǩ�����"I�ڝ$+p��A۹l��$���;��45�iy!=�vO฻�0Y�O�ߨ��$
I5Z�h��ڶ*�X��}�i�q���d�Z��}��v@��<.[��a�Ѹ�L�"y��=W�ƛ��Lc����Z�+Ǥ�A�uW��@������n��z􌜗���m!�Ξ=�m�ncyoI��8!�I,�A6�~ԗ$?'�%�9yb	�aT�I>�6	��Ǆ�z�!�N����q����2��S�,��������8V�1&c��-��y�c�/�I!*yG��]>��O�弻����4�(��F���� F�ZX��i���b��/}�i��B�U�l��/���,�b�.��ֺm[;2�mb|f�Q������ˋ$~�ۓ�/@���ϕѶ�-vy^��
�I�*q]��'��1��l���̈́�W�ǖ�����������q-�l>δ� ��G����ˈ��-`eK��"d�e��X��:�u��I\�"䫉��:H�>V
ͣ]E������.������cυF�V��;X�B�t���z�c����1ORP�����J(��$�<�8~����c�Dқ��+F��k�f�;�\������VE5܎6A���%��a������q;.N�ѧ��-Ȋ�����bέ�2��Za��My����O���}�YP��l�8���~���&�0��;�l��,X�`��,X�`����y���C�g�a|a%ɧK׏�����|X�}?sVp;���SӅ�r�ri&KrZd�����<��}j�(	d�Pz|Q}�m�Ңz�y\�J/��%�@"P�	���y����ē��>��4*�F�vɧ&5(�����I�d׆���4�*�Ю� A��r����6�ϔOY5�1A��W=WF��j>�u��ΛCrd�Q�H�i�F��86�j�d6Z6���Ƶk��}�qww%�L�7dpk^��!H�~D�.���hf<���Dہ>.C��T͙�b-����K�`r7���!+�w-?f�3�1H��c��<��<�%���D��ZE4Gx�σ��ͯ�F��Z���\�h�g����#B<<���_��4}�U�r8O��%d�c "xD��'�6��nG��뿝�����?!����[�'�	Qljf���Z�[�ׯ�u�>���g���V���I������q�h|>���ɲ�������fT˵�#N��;�7Q�,Y��O�_�7�^sۼ��v���$	�Fɍ�\�\m=[��;R����%D���?�@P�����=���q��yA<��>�H8j����L�H�$G�g�MD��F����3��fT?F㕿��1J��A��0گFOdy���Uf�$�����P��f��	�yD���9�1�W�q9�*�I�=���4������m)�K�ڕ�?� ͽm���ھ#���%���z��w�췴,��19�I�0'�j���(�(�'�|޾)�>j8����A�&V���0��-�<}���X�z��Q��;��o�K�������d�!rH�޺-����'����@~o���lmɊ�7~,�r	�ty�����וq�ۑr����w@��c�"1�bly$��RZ�$��N`\%�Q�w�)�b�s��G���@v�~x�L���հ��h��a���:uh�jX4v5If�3�����#�=�+��8n�����m�Ro�@�RS���DC�+�����"s���4m���\}���~�O~ҹ.	N�_,�*�Gr��g�W� ��m��\�QE�,�>m�K����Ԫ�ڗ�VP�t�J�������}9/˙ϛ�?�g���}�\TRϵs|C��Z����|V2lrȉ
���=nR��W�؎���Xc<p��5�GŐy�ab4�=3��^�z̮P�w�w\i@����j���qe��pU�}?)��z&��'E��`��,X�`��,X�`�����$T�C7�a�p��Ճ�Vg�#��y���F�ٿR���!3n߸���Q����t�~�`"^?1P")�y���	0~��k� ��zD"�V_Y61:�x|�M�����̀�/�Z�'�w -�4_N :[�(������w��ɏ94�k��|���y�l����>���4ګ��S-ǲ��=g7zoF�Yb4r��|j9���[��;�����ѕ�i��P���G,M{Ўaq�RQG�+9�a���_}�=���pQ�&1�Od˕�������o�'�ZM�=V-���T�¢P���f�DI�2*t��{��F���z���>����I0x�x��}��R�zߜ�64�����l�v�������-�����&߳�>���x"M��K�������4���X�J~;-�n�!���e����>.����!Ow���c>��iF��D��'�8������������ٳ�h�W�e�(��T5�����|fb��x��fǍ����6�LϯՔɅw����~�(�,wj�&n��Z� j�_��%S�_��\Ɂ�'F��F�#ۿ���$���xj4k��O�r����n��FWU=jw!:i�.�u3��<4���5�&\����	����7��*�Ϛh�ڎ�`F��p��\��h� �j�&d�EjM�A������AB1{���ql���$�P�bw�O�F�xB���?vʥB�8�3$j��JP$c�+�ۘ��ja�>0��������
1F�bg�^�Lf�]F����(�c�h@�bsW���������B�e�j�&������Q��]�[{�ʋvv�h�ՐO�v��F�l?���j͑�$��\��4�ֲއ�+WƐ(��w�:�F�rLҰϨ��:;ג����%Un��on��$�ܒ�D����\|L�h�8��i�)�_�#�]<��C�����l}�D�^��D� �4��3OI�u�r_lP����2>����~���>#�/�"Z/��6�h�s�4ՠ��/����bH�����iX�s��/�����s^X���v@���g�e��Ǐ2ȣr�F�����D�դݴ���>�ΛX�����4�����yN�y�t��h�V��U���Ԅd}ՕV(?������/�s��_����t"�	g6�/Q[P�M�c$��qՍ�Kr��OM<j��J���)�
gԬ���^��S�<�D��_�5j�~�B$|��.v5�G��U�<��j��?U���V&�V���a?;��$])���!�hǜW�f�2 ��{����8����,[\�Utg��,X�`��,X�`���!0�>��6Q�˩/
[�~��~�~�\��" ��IP��Kz�7��n���D���n�:Blsm�9~fR���9� z~M���/�C�^;���?O�,���u���T��6� �Լ��wz��]O�jP*��d�rD��!<PW�n���uj�$}��e9�����,�&��xԬF�������?�+=$V�ȧ�d��J�e�/��Qۦl�Zң�膖��S��$��#�*	<�����'��(g�؏��~'A�� %!U;�4�"O�Q��!�0�t;F�"�0"�ݧǛ����\�)��X�ц6<x�/$��I���Le�[�JKǠu3t5?v����s�f�~G����K�A:�Мk�q�@�},C��ª�����o���ge�X�۟���o\��F����	i�;ץV���*��n	�2|U�o�u��S�r�dn춗����q�$c>�(ω�#��-�ݑ~�ϡOnDr��Z#�,�o�8���^Fn�@��j�Lrڂ�����6��t�y��}2"A��>ϴv���m��~��D�Q\��8���<N[�D�G$Fל�H�#��!X?��9�V���f GF��� ���$`4�����^v�(F�UmY�9�d��h����]ih��ΐũ��mkq��W��Mb�oQ⹞�}�E�1ȼ���h��U#��ˣM�tQ^u�5��f�J��0%Rg�H�ޕ7E���֡I���{rF�F.	��R+q��Bsd>�|���������s�q���e<��_��s8�/�#����J�ƊGE�hv����^M��O��po�����'� �CL��+2P@1���~N���!M�]������I�G-ۏ� ��Ǟ~.M�_�~����GM�g�/��A.�\9z�����~�iz{C������
�-�.��^N�����?�t ����C�����2�p5�*:�n���K8NN�m�!��j�2Z3�c�Q�AJ����Xv�K-D�ݕ�����p~w>����]�'OK��Υ�p$�o�<y� d;d}f��6��j<�8�lm�{,���	9�����?8�*��G��;L�y;�,r���$�J�森p"m4����F�C��:�Ej����D�YK���Jf�1�"���s`�Q�[�����:V��}�ڇ��yyI��j�Z˽��V�dW� �������~��S���Y��<���=� �}��}O�ֽG��#�?�<=q�K�>gH?��/X�`��,X�`��,X��� �f�:�c.!�4��/J�}6�A��%��Ռ+��<���?bt�!I�O��wKt�~��I����IQ�X����B� -f\���4Y�
��C5�cYq=+��0���x
�u��!�GR�ֆx.��U�A-@De!Ձ����el#ژ: �gݴ_����|0�z6�?�����g+�@3��=mx[S"���<*��kT�u��Y<vL�wZK��уEM(>Wa<1�I�PK��&�*+��#��K����8����W�I��+�}[��:�֜-?nSSJ=�
�}��I�=�L���5�u���^G5�$c,7��&���dS�ԣ���`8�6G�|��O�M�!<���D@�Mؾ	\���KM0��Ύ�o���G5x���o��\���$C�$!!G��xz}�I t�n�x^�c-���(sԬ�GؒR|��|Q���lxZJv������C��=��}C���֜Ȥ$e�.y�N=�$�4����!X^��vTJęq)���4��T���[<���k�ou^@�Y%��x43I <���X�kG�q��4)I�Nwy�ͷe O~DHVj8-A����	Y�p�;�w���]�q�� �ӘZ9�]���l�֗�on���e{���[|c���߭-!d4J)Ɵh�����GM�u�S=����B�2���'�Q�"���:�S�(�4�v�e�o�?`P}$O:yN��[�6(��W�����-���f~�gp��R�C��r�~kk�Uw��Y'� ������u�w�g1�yh۱|摏E��ΝE��菴.�Y�i����E�?�XZ�r'quю�靭0`�Y���+��i/M���s��_]��OgW���?�9�,����	����Λ�M]F�Џ=�B�~��O����?L�k��y7�=���~5M�G��o��7����+i���:���?��4�nK�HZ��_�J�~��?��}���
���wu�R<��%��d�~�K��:{�{I��Ӏ�_��#�����4q������ՓҿV��_����9�b�X�K�0O�8���:�W��}���)ls��Dtl��PF��hܜ�f��%��r�ʬ�P�QW���{5�� �y�d	�Z����Đ��S�=W�ݾ�Y29�B��y�;o�\�=��v?B1@�ΰŌƞ�G��\��-g���i�_����rbt��m7Yn{xOgc�b�/7�>�~[�I��#���d���fe�G�ܷ�/k��M�S`��,X�`��,X�`���!�J�
ߙ�����17+!xX���"V�e: �K�Ɉ���=j�Y��nǙ���s_�}��+�}��M!�6%�葇aIt=h���sW��d�F�b��j�vV^��#���V�l�dQSᣚ���X�''z.&>2�����z�'���������Դ�&Y�zL����d4ʒ�٢�@Y�55Μ��kJN�:ۈ.GO<5�M���(wЌ邼 YY�'��_\6�U�X�����reC���a������(tcDo�<Z~F$y�vM-Ē�N�xdy�SF��W%Ơaӑ�&ǒ�8�����&�|�#��ׂg��v���3BT�S�~$�9B�*��&��*<�F��@�F=�8�^O�������f��g�ր6b�my�-C%.	��&y��@mG�G}�'E{�J��� �2=�|^#D�c�3Vɘ�S�Z���LL�3��K�������>C����b[��4�5���O�i	����K��V�̡���M�?�y��8����85x�v-���ڇ�KBR��k �XQ���2�ᾴ/����
�)�_�(Q1�����)!J�g�oސ(���o�جiTA�~��n@sU5�@b��j ���� jq$z��Jb�M�γ�Vy�2\!A�vPI8��❻�6!�d��)s������)�������c�OsK?$YZtIiF���h���Yrtw[�79���T���x:������pI@*y����q��5'_�8��?n�]>��'%:�#�t#I�y5�N|T��.�+�V�_8�\��B���V�G���m�ӧ�)��c�;IQ�4�7��R�IR30�'W����{kS�)�x�{ �v�O�]/.�|��<�������|�$I+ _InQ���*�'�Zm�g+'��W��y޻t9M_|A���D{���!���⹽��+�?���sK��k :��I?�GE�o�l����+��9}���iz�~K���|穋R�9����@�������8������X����'9�F�,���hό"��EԖ�u�h�Q|Rr瑜���r���G�/���	V ��f�In�ښ ��n̓�� d=�<@����Vue��������b���jֱ�6Џ-s������G�٭m!��췰R�D$�9/���|يWK���E>u%V��;h��y���6 �v����В���t���
�����~���E֋�M�8�M0p;���V2��[[���HS�M��h��6�y�y����D��H�A3�4����i ��,X�`��,X�`��{���/#W����Gô���E�	d�I��~��Y5�|_�g���#���qhˉ3��5�ZԦ1��d����/?vɞ�~���>i��C&1����s6o����vW�5ϒj���1��BTV6��>�yx�H��u�-j�0�#=��W�����G>f$I��/���'��/ze��le�ZH�:������]�x2��r�"��D�Q�������M�"Z_��%)����ٸ#�b֏x��@^�v�!s�F���p�?1*g��A��d����VQ�����`�J�7*&�+�]6Q�Tcr��o	�۷qY��Շ随$��a�D�j����{
Q�o��Q�s�!���;,A��D
��&8R%ehެ.	�p{]�������K����J���1�1��(��(�4��D=��?��	d�S��x~�8�k�i���a$��w���zj�@�PSE��p�z,ϣ�`T���mNL�NF�&!��D*�t�8N�ލH�<��p>�&�)�,:��6f����V['��ǟeT5��^�	��M���ǛVN8�[2��r��!�#��jG-Fj\��!�s�MѢZ{_��W>�E\A�:�G�W�����$���`��1	kF�$1��(Ш�󈦇��������yQ�Y׮��H�9D�.���;2~�A��@��J�!��E0;�ҿ�@��tf�ͽ�t��ߖ�vY��Vq�\�}��7j��ہ�)���@��~W�/5�|+7hj��;�2/���E��>~,���~����+�,	��>��]|��4�}S���Bc�ُH4��.9��h�</ɾm��Ԁ]FJM��!��7[�wu�#���-!t��pD��3�mg���r����Yh�mn�y{����?�����<��'��	;�<t��Q+��$A#�shO��Qc��۶�DOϻMJ>�uhϒ�Y@;~��kr_m/N��L�zI� �נ-XA��6iJ���,�}<�6ʯ<����Cr�c/
Yx�I!1o�G=�#�~N.K�⼃$��2���e��H�%5TYX�Hԓ��@�8^�+�J?@�I�GI�a%��,�{M��v<�
	�����+I9oNt��q^8F=�_mtڥ%Ws����,�>xj�֪��%�Ͽ'�?���G患�$Q�h��$��r��H�\��s놌GJ2���b�[h�r�<Ɨ.�S���c����DW����G�Ym|�yv^��<�����$	7dT���`����%�D(����͕k��"��M"�х��H�X��Y����e����w��}��4��,X�`��,X�`��,�C`}Ӊ%%J.1a5LԳ��Qg�h��t�(o?-��g�&vrR]���/��&�@�z�J��/�\s?����k�+�=���㦶�ə��t��x��A�=�e�E���d6�,���≡&�$��@�\�Dd��'��5 ����MD���=���v�A���3%A��ZFS�d�=�1��4���XN$��ʢ�Rc	Q�sQw��k4e��i&���H�Z"�M�6�CZ���*O��9��j�sL- zd'�ߴя�1�y��%BbŞ���H�@��d"Y���	]�D��$n?A�M5z�h�.�g��� ��e�A͐{#S�=P=�4KP������b�Rk��ِ~ns[���O�п�w����,���W����ϋ��~"���%�h�Q�'���ZmH���HH������zdI�̣������E���x�ؤ��F���sBD�>ϊ�s�HS	T!4TC��:eQG���Y���(U"W��dI�:ȉ^��ĶG�HLy��79"F"7ɡQ�h8�F��`��kr�:1m��1I��%ry�$"��H���|�&��(����i:ؗ�~����ɲ����	Z�'���7�:��D	%Y�~GHFw���P�}DO$Ax�����A�i?�waQ���q�B��� R���Ǳ�%�{l�8�G��pm't�C @�'����GM��t�ڑy��ks�urA�#$����z(�kuiݮ�7���%D!�Z�x�W3[�Oqc�8G�d��!3�����HP���+K$�����w.@�v����YUh�����ǩ��+Z���	����[�}\��
4yww��|�I!	�X�ߩ3Bz�{�2�e���<�?���������u���XP���w��{$�h�Q~�� �nK�|�W��m�D�)Ѣ{��(,�R_���z��K]�����ܺ!�nsn�%�*E�؏��"����̻O��<�y�'��]��ݦ��3-�������'/��b��xQ�kw������ٗr�ِ��J�f^��c�&$�9sw��D5�%#��2�3�t���.�����8�� �P�;�\������Hλ���kA+3A;���~~woǁ��������AL�yA�-�σ�;��j���s�V�߿��߱�	"����k|n�W�v�ҏ�P��ۅ�*�#��]j���"¼ΒLWC9�l�V��c��j+S�X�����v��y����ghV�Jpb>EQ�q#3���cw���$�LW�����I!���o�o�����'�M�{���s�����8�,�y�%=���` ��,X�`��,X�`��{�R�M��$�>�fۮ-��
��,�gvω|������a���7�:g��y����Ԓ0�٢�Ğ�W>�O�nzѪ��q����2�,Q���Od�E#���j��Ux�]ף�i�1�=h4"!O8��@"mo�g��OНu��1�Q1.!_��f@�DR���������nMO����Ԁc>m4�!i�'G�Q{�z�H*��Pێ�i�K#)�M#j���Q�K5�ꌪ�Fwʹ��G�ҁ�����|4���uΗ�ޠ�ȝހњqZ}�8S�(�,�,�;6+����!���V4�Cݐ|+��S������OƮG�F��H�x
	*gà[��9dP���4}����׾�5�/4���X]��-��޻t	��.�}���ԣ���}�ܯ;$�+h,@��u���t�.K
�yy� =��j�O-˗ڕ�(��䟍�6���\�3ܝ��V���ϛjD�+k���#�7j��]2Q�%5%��h�*'���jkZ�}�'n����Źv���x��G����rIɍz�E��8�W�O�S�ڕ�c�CN�������QnI`-�~��{9D��?��r�5��t�[@��hU���I1j��N���nR�X�: 
TcG�n+�䘚t1ʫדz��(���V�a�C���9�NV|{WʕZBsK�O�{��1���.ǣ����)��y���8�Ŕ&�������z$�G�@:��\^p��̸���yY�Q�R��%N-�J�i~ڍ=�n#j*���_���~�� �6��8�P[w��6�Þ��F���矖�Df�%h>>�������k�,�D�O4Χ�W�|�XI����Ǖ6��&	��I�����;�PD���ɧ�@dTMN�[(�5�}��*{�4mFҮ�"(1/ �Z�8�2R{;h'�'Hj�_c��n���i"���B�|p]�V6$M�oA�!?m�X�xz�����R.W�������4D?;1Q�U�_������5h�wE��2�f��\����{E��w<��c�j<"!:}<��mwq���;�WU��x�#ۤ4}Ŏj5S[��$"I�Bj�M�|O���
�3��L�c��G� �G#j�reG✟$"����{]h)6-}$������l1o�E���N�*�kދX.]h��A��S�ʻ	�Г���Q��Z�J��r�����x�C.C9�����+�?���(�<�ﵬ�&ʬjv��R[/����d&����c<���s��������߁S>�N"�њIr\f�h��h�b��<����gZ]����U ��,X�`��,X�`��{�}�I�I��B����<�����.2��h��ܳ�@��z�4 =�k�iѹ�Aڃ��<<W���bD=�${H:L'�M-����)��D�]\��&�}��HŢ\"m�b�]	ޠ!�rѡf�(�f	
�mx����y�!��zF���� �ROF�~5x|z�<��lR�Azh* X��Q%����(�F��ϗ�i����]/���g�W�V�K�Z��5�q�S7����e4�聡�d�Ҳ<?��	O$�dQ+lQ�: ����(h  H��#Ĩ}[�<���է��'�u�����?k��h�&Z1�#x���h���jT�1IDӊ��5!��B$��Y�M�	3@b[F�e=[��!�	��U��G-�J�Z���Pk$���=ʣ�����3@;y晏���1�W1�������^�}d�F].c\scK��;и�������t��~oM�w�{W������7�,��;߾f��3kߺz�[�0!$Ѐ�@ ��18�"۲q�=1^���cG�'0����0H	���^��ת�%+������}?��9/_gu�g�����N�|��{����}���}�I����>["����:}?*�#)U��H������L���z�74-�x&RMG9�I��u�0D�t�x;���3h׎���9B3N%!�n�Z�&����q�~��;��c@jG����Cu|B6��o��n�mi� �W�J[�Mj���_��(��N�'w�yW�n\��X���ܩ+��_�(�m���]Tz�'':�䚚6�(����n��� �_M��~���CU�C��+����voJ� R+��Q)I�Mٕ�\���ƅm��7�Z�"�EEE�� ���EN)�`L��"�_1B���$�*���#�;{"��4N��L�q�&亢P�aF�[�H���Ǹ89c�#5�E��4�/���� �y�(�jY�T�l'NY�|�s_��{�v����G��+Z��Unh��tK�urY�c�8�|�_gC������|A��j_���H@{�����c�Q���8�:�H�e]�����i�mi=�FF��պjoW�$�k�mH;�ܹۢ�6S��w��0��S'-��i�1�J<��?���2My�Ļ�.#���f��M��KF��X���N��(/O[;�Ԏ��I�֥58)�I��#��&�����uc^����Fe=�I����Oи�y�,�5��ˇ�d8e������TJ����X��y������a�{�s��WS��ڪE�F�tw��i��k����i��|�q�V�{�����s�l�Ҭ���O4w3�箢6�Ç(﬋��߼�w�{�R޶��Jk�u0;�$N�W��w�A.�����@���b���ʿ�G���3k/�.��G�����Q9�H�0��5��|N�^��A��BR�A;����uiY�{��]b�`2D���,��h���c�r}㚍�<w8�E�}_Z�	���k1�[l��[l��[l��[l��[lo {�}>��ӛ�>Aݫk��|����d:w��6��t�"~��d�^��d�ebϽQ�bb�5��޸�~����0ڦޘ�>g�Mۡ!�ʒ��]~�e�.�N��x���YE��O=��6J6/��ގ�߃�ߑh#[ �u�9��`�j=��#����U��z��ş[�EQu>1;^Ꜵ���y���2��G3�����~��mH}����ܟ4(2�-�V��<!i��	;,��#T��!����<�)W�h	�F�?�N���|t:~�@<ѩ�ՃoC'y�ڈV~h�,,��Ȏ���`Sxl�D��sg�tMQ$���Z�r������[���}h��_{*�.,D�i]QK���t\�i�)���/఻����?�'����(�|ϠӬ�i�n!)+�/뷇A@�VETT�S�pٗ�u RwO�P��짭DL�Dt4D�f&�d��%���n��s���S!��=���n����v�������'͝�_��dZA��~FQLu�|?�8O��j��S�,�dݺH�g��{X>��e���<�� QP�Z�1.�+�M�C�uq�y\a�nNn����?�2�NH���=�JN[-(L7n�:g���v哔C���I&��?��(�$��l$Р%"��~*�B�iA��Ԥ-63Q�B"�� �|u�h��=�|G�GM]���Wl]4)�\���<�y;-���}M�N��D&�|;zR��5��JTն�ɔ4� �׮�q]VD�&:l��S�/�&�?��5�����Ӫ��C�K��DZQ7��w��@�4^N��yrB��H����f[�~�c�Q���~�������.���zꙧ�ta޴S�Uh7��Z�h��Ys���[ȩ���|���G�l����K�����~��/ݸ��و6����y�� �"����Ż�H��H�����i���˺�cj�hh����N�toC����>q�PQ�f�4R���#W�Zw^|��(}�Q��}�7�3J���Z�������O=��(-�,�hOvz4�v�#5�nf��v��;��詓*�{D$�h��Yw�����EK;ivm �XR�e\f��<{"��h$�劈�?Tf��@���Ne�_�2n��#����k��{v��d���V��;n��f�ʇr�8�?�z������7�/d�^~��.B�sF�����KQZb�+ª�v��96�ܼ���������v?-r�zO����(��V ;۴S͇%4e�s����H4�P�m���J��!xtL�
;�����sڭq�"�4��=��n��ml�CK�e��9�U����9��"���6q���7Eܝ<cd(��}<�#rme%���w��WS$f&x������!/.b�/��b�-��b�-��b�-��b�-��� 6�E�0ʮ<����D׽y�ǀ�f��y��Y��8ͪВ���#�|�4<�.�7�x�jz�WVo��d�q2�}���>���o��a��c���"~QW�Uis4���zV��F��Ͻ#>!|� �]u[�M�<�y���y2Ҁ��'/'MިWk�F�Ѱ7�h@B@P��r.�D�!�и����$�����i -��H1u�l��������=�)�>4
��0����'�o�� �)��f���VyU�u��i��T�<oCr��mHƘ�]4,?���M6�Ct��}�#����5�R�iD3YX0���+�N��W��!�_0" ���W��8y��I�c� ���t�gy�!9��/d���^9�=\C-�ԁi[dZ[Q�:�O�h��H?���8����?�DIUO8�>߸n�*���S�=�v��w��Ec[�aZ=���v�y�#��h�P~h�L��1LB*e�]�vr�]��G�('�<�� h�8�%yB�EEsS��톍gD��>!ʦ�[�7���C�K��!	mi�c�Mf դ�~R�s�]���vN{Ek'��Ć㨏\�鄼�@�Gk�����q]�>%M��)�G���OSc�!�7t�W�D;uV��0g�xW�H�����:/d%���2uD�L�뿚�.-i�u3 ��'>�&�� I=�g�Fkt�Ə!)o神�d:D����%�|�+֯�7"hM�Y䳍Ƨ+YP�NKX$J��F�O,8�E�Y*[d�qQZ'|-�i����k�n+��Ut���u��4J�����n~�1O�ׄ��*�)�}h��p�54��P�-�&��y�w�E���C,���gR��ٴ����H�v���vSG랕�V�!������"Q�]5��Nʊ���d�e��¢i�H{�!#����ϬO��;#"��+"�榍�j���]��_2��mo{�>��3QzB�K�G��=i�]x�v���X�H������.�i=>��\�KiF���C�g�nf�'�/�fK�����1���)�8$�u�i�j<�r�H�Y����l>�}�9����֏X�Wm��ٖfYCZY;�V�%7)i�]|�ȾG�fdߩ	���Ț[�N��a=@�I;Y�i�e�xy��e�n�8��mw��R�u���srZ������K�\�ϐv�[���=�O��+Sv^�hR��g���i�\5�@���]�����@;ے6 �)�k<$��_^�u��'�<:�N�VZ�h�2�B���M�G�]h�nw�������G4��ȶ$ϛ9�=�#5����=����<�-m�v(S"��K6i�/�0�F_N���{4�<"��_�������h�i]�u�@ot�)����K&����i��hC�3��"�t_N�;N�\��xS�g�.�����3��{^`�M���"��{hj���3A�q��h�7�qy_��(yG~&5�C��6�ݗ�Ʀ�EI��U?Jy�#d�@��$�m�����H��s��֑x��sc�/��b�-��b�-��b�-��b�-��� v��>X}D�u���0�}O�|<�#$^�y��8�ʽ��E�<�h��Q�P����W��Hē��3�E3!OQ��.&���ky�w�q��?���Q��G_����jh&@����C� ������p�g3G�q<�Ґ���^��x���7yٜ��IQDˊ�ɭ\�ƅ^���1��'~]�6x��Ȟ ��!ډI[��r�dv�Fͮ�G�<Q�ZD�S��d ;sʿyx��m�/^���t��WyV�0��ˣ�4t6G����!b�6�O@��PU�'w]�X�8��db#/�"	������oEOD��b��ac�H�T�߈�H��E�)���Jtd��_����м9z츮c�A�@�m��uD�l�;oC���-e��h�)�V�'W�n|�>�?�(o�ı��-����E�-HKE�JDG�9�W�4�،�J���h��"��w�{&�v�<���D�Y)��~�r�ƝEif������SI�����\]󮏦d�4��y;��5#J�v=E��ˣ�	wk��OC��*��nد��<�hr�b�� "'!�fda�a��Ii���9E��q�?���4,UOmy�D�,�}���mJA���]t��i}3"�>Ѫ��ߖ�qNjH��{H�M��� �8dBHP�m�
�lX�h�h�Le8����ӰO�������:����`G��c�?���A֑�%U��&���S�s"�$��ϩG�\� ��B�˰��[Z�feK�h�AX���a�o[y͉�ʋ�몽����U��#Gl�h��Y� )L�T���(���h�J+yg� �6�D{c^�� {�J3+���pF�͡���\U�����zG)4DI�ݸ�G󰃶����~����M����=���ӊv�@b"�^It_�O�EI���pǝ��%md�BrW[9E5f��?������dfrZ�)�S��t���ܾ��sQh"vU֎�V��H�����׌·VdH�E�9ͽ�}�8�ٲ�:{.J7��F�:r?E��<8='mV�/v8��YOY��A��$^����KQ�~��I����E�e��x4�uj�U���j�_G#ʌ4����⩋Ft.��Y�[)�خ׆�STU�+�?��{ƣ}�h����v�+�������w��D�f|��8¯�/�_8b�S�W]Y�|K������U?��s�U��;��.�]�߻�Z��T4<o��Nc��jgNkW��>Ƴ��v�0;�Y�h�'�rO��o������Ѱr�% %}�bv����)Q^Yg��y��f�AG��aN�\ω�`\��{���Y뗤�\g��섿��c~�kݞi2�ZaG�V"�+;��!Z�H9��v�h��&6.&�m�g�Q屾�����������z#���<�B$@��9Md43�>�������0l��(���[l��[l��[l��[l���_y��}�M�<H�y�u�j :��X���� ����o�:C��%�b)4����-^a��w�8��h�4 ��9���b�<Q!�袷,芇߅ZIAI9B������V��#z�ۼ��+� Ŷ�eÙ3g����1�{Ҵ��8a�������gEi4�혇���|�J#�v51m���~�^~H8<���Bn7�:y1.ω#W�!�_?�=�N����H
��ʔyTץM4u�<mx ����Vkv���("%�E��$`GoP��<1/��>Ci��D?����Û�8�����%�5/O�1������S�hƁ���g�eCv��	qh�T幞�E����ۓG���ѕ��n�Մ���O�=�ז�hr5�����v�IZ��ZeD�Z<b$X6k���K��-�%z�~C����G��q�h�ݖ}��+��V]יU9:�O�6+�X_�KF�\Ța����ܨ:��@#$�!�!/I돃Do�|�Q�rj=�{5i�O�Ɨ}_�B��Q�FCY*��Ҹ�=�Qw@���&���yt��cNkב���DB�5!��v��g��*�B$*Zg�N3"�.��b�NB(�<S��"3�5��~�B�S������j��S�Ѽ�m����+J[�7�r��A�=��@��ku�dN��p�/Dc�:#R8/b�$��FԌuU�����fݠ㯏�=� %����< ���dԤ�JӒ~��k:C�͎N�����B"��vrd��=h�%D"'��"'�a6�j�<1�(�:��:,�1�����߁�k�9���~mmU���Z���1U�x�����Ҭ�`����=�hM��O�@&RA�{�N���:�y�(�XS�x�G�fY�ɐ�hƅѳk�H4��޸a;A��u��o��ť9���6�e:I��$d�����h��y���!-�,��s�v�־�Ê�亨�2��o�:y ���6ڲ����0n����l�����1ފ��8�B�\�*G�j�ʨ~hO����4��(�lA�Di���-BT;xXq5�^h�7�v��%G!Y���d�H���8s�l�^��1�ڮ����g��[a��}Gڵn��gV�We�_����������Y�Ή�N�|l>�_u4�]nXb�~��+�|g�Dg��?<�ծ��7��<�u�0zx�����\����Bл(���N@�k�9�ND_������Ӹ4�9���������%r"P�O�|s�۵	v�0�3ΰ�kZ���joE����������9wzʏʛS7�hݩvו�:�?�I4�sD_�v�:2����*Fk5?��$�1; 1�:"�ᴽydh�E�u;������Iv�4�>�f��y���E��\��R�����U�ǚ_��а�7�zٞ�7; ������a����`��U�߃(ǔ�##O�<�.�u��I��Ez���-��b�-��b�-��b�-��b�-����[f̋��� �	{�7��姞���Q���G��X(=��Έ�A��]w�88G!I�3|������LÌ7�GϙfĜ4R0�'�����:�7J&&��R"�6��z�+O�>,���`'o�|&�����:����Ɂ�*�iE�}�ًQz�y#'�&Y�5�ܤ�Z���40�����Qr�m���l�>Ѯ?%͎�9�@��ˈ�_���@������(uъU^��Mif4��t��i�]��{��t�_AaS4�@�p$�$�����"DDA��z[Q_�v��}3��g|UљE�Ֆ~��[�Q��n)�YV$�ɳ�9�����K": t�i��lHR�3p�i?�b��G<�Ҥh@&�1B��'���!ɑ�?�ylZ]<8��t�<=h$���fd�7U���ѓV\�<�Yy�h>{�5�nF�""l����G�������oY��LX����x�I��>�T�/�%&GV��(��XUo��4b�����Mc���(W"�R"r;DS�В<�i�)bH)ڦX��h��VohF9�9q����=���G_�D͌��ߩ3Fb�N�V͎��Ο7��UE���Y%�L��i��R%�h�HU���<�=c�zi�*duݶ歎��W�O����^�y�i ��E��"�����Ξ�ΥU��|L�D �N�D�h|��E��}R��� �-?;����4d��Mxǣ�E�ƺ楁�CG�Sh��J�
҃��h�@�n9�2y��������h�S"��{��O=i�̈l�+�$"�U�ry�]�9�/D��<=�Gr�;���b�n^W�e�w>t_�VDl=�j����D�~�'���vm^юvW?\g���KD�GsV��L޷O\P^9)~N;�j�S��ٲ��Ӂ̨�dS"�,Hӓh�Y��i���ZC3Q^�o�RѸ���A2��U��jQ�?�"D��i�.)
";&��̼0Q��&h�=a�ݖ��ci����(�.�!:�v���K�t&�2_ۧVMi jz�m���3�v�"��+4�&��!b��������	4sC�v���Ȭ�_�Ы��%; ��ZOo�z�[��sZ�3��@���C�q���&Z�� HC�薔sUWM�(�]�h�At�-E�T,�=B�NXQ��];���<a���9J���qaO�$�)!�Y7:�I��M�O.�+$�H��P��~'����u[/�4es�D~�W�(��[�wDӞ���D�Dde2tk��fcV�E��p�1I:�?�Sڱ���9"���%����q��;�煭��M;���1��B����R��:U�/�N4�#�i$��C���&�<dw@������"��>;b��gŘ���jF�u��?�웜������ ��k�7�{�g���~�u��<��� �Y8�έ�OEv��G� �I�K��M�>��R�Iǂ�dS���N�C}4�цU;��������!�N��{kWݮO�a�_!��"͸D�C 2���Nay�ڳ����;)�}��7�������H�c��Gݍ-��b�-��b�-��b�-��b�-�7���>޸-m����kW��r�"4���K�y�;jc��M������.-��-�222�7�yCr$ሖWSZ���[��`�˃�䔪��#�vw�÷�oo�!"���f���/GG2�-����;�+���'�ʅ�-�}��x��/m�zf�����ʡ%䳖Q������7�7�ǿ�]��u�"��F�W��?z»Oބ�(�Ⴂ��I��}�m�#)$D���"��y��6/M��w�����{n���Ӗ��`l��lL5�)�Y <A�Q�О��_�����ۣO���Qz��w*�9�I<��#�:�A��Q� [���}�}���_�y��6�~)��e\�S���O�fm�E�OH���-&>ͮ�ƍ�����<�r�M,�����~��k���q_ǧ��t�Lؔ�X�`��'1#B͢3�A�LZ���#8�6EQZ�=�+2ka��OI�����6�M�^��Dkv�d�<�@x��uE�-U��8k��V�Ym������o���ā�jAk+!�~�n��r�ƕ|.�8�F�Ź�E�}�GL��|-O��	��ڰ�����ь��T��GW\G�j�ݼ����h�)ߣ�4]t<��'�9Ȥ������}Χ e��z����F���>3<�~9��gI�W�}i�Q h�u�)�v��4��E��(�*�M�l��m��V��miw�?��mɔ�M��QN��8��Z$�ȌBُ~Nt_4� b��~Z�`d��Q#��/����ĉ3���)k����}�L@��뢂��g* ���KG�Y�	�A�r��I#�.��R��4�3�8�O�vU�C�=�|����Κ����$;fW[�P�կYA���&�H"0��G;D����u3��ޖ]��������_9��k�k6�H������u#%+"�o\�u�'$Ӿ�PRtʺ��I�ݦ����t�&rG�k��=P��Dno���J;uʈ�kWl�w����г���h�Z�$M㊵�ZM���v�|�"� >]�m��D��A�}W�.��ѡg�}��D1�8�R�)B�
�Ѫ�;IG&^�t)JK�e��rگ�h����񐒗_��1~0� ��٠��;�HK�.�﫯�����]�~LT̎�ˬ�}s]d���]5��?U1���g��Z�CJU4�e��)h�N�����u�i�M�~EǙ#��%ͫz�#7.�%�Kf|��l�~�q����z-g�s�$�d-ߔ��:�� GC	^i�A@�tsC;���X�V���UE�g4����a/<O��
+���5.k����W�ls;���ؑ�&��m�׬�Nh�]0Mk֕}�7(�]B4�5ʺ���T8��ܕO4��V�=��)xUѸ�WE���(̌v�t�u^R���+ѴфO�g\�9nd=���G����.��i���:�b��ΦE����4iK���^�,F��R�i<w����>�Ƭ4��9Q���)<��hB�RN��wBDx�哴NY�>��:����ο��Cyd܉���b�-��b�-��b�-��b�-��b{���E�8�`�5o0��1�[M{������:Q��F��>�|�1?���Aou�sw�'�(���M��"z�<�S5�hƸ�0#�1���z��;�t9u��8{�"U�^�-i����gn���8IA<QAT>��mJ�@]yx�?lځ�=�p�n����d��-���R����"���{�L������vT��7��	{�~�#���^;My"��yRx�mA��ǣ���-GY	����y�gD�D$Mɣ�HX}��w��<(��|NAw��H�b��ѥ�x��V����<5���ЏFi6K4bE�S=�DE%�~��iA���/ѿ#�H�S�Kf���W�c)�+yx�д��f<I�o��k7\4ېzc4�Kl�E�2V��8I�:B��x��5�5��0�����H;���"b?��EiC�ҔȆ�ȃcG��)�'x�\�\�m		�hl~�B��И_i'�xeb�|"���8��u�ˈ�;��ј���4���뿖q�L�94FOGF+u��n3��;��"D)Q����� ��J	����Z���4OJ{��{����we�	y�j'N�N��o�8|�{�c�W��=j?��
�T<�Y»}�~ZDsZ���/Zc9�?��O�1�WD��t�>r�
H4ӷ|�D��� ;!���m&�jI�vy��.�?�Jt����w_���@E�E��Ag ��頉c�����^��'#�d(�
���G�p@���#ى��g> ����A�p�nןO!�Q�z�?"�u�v�<�Rҿh5�(�"����u��cg�bt[�7�OS��o+"(�#"��A0(��Ji-A�&r"饵�IG=M�r�\FV}��d\�Z3�q�h��(�XE��icň,ȏ�mE�M�� Z�GEA�TE�5�M#�/���W��l.�e��Ѐ:{���N�sK��DoE[�yZ��tج~?���3N#��#q�A���ݴu4���򋗣t�l��WkY9��vֵ^�0�u��]�Ry��<9)q��j>��EK��P��Q���07M����i>]�������q���f��sC�ᘕ�[��V���vd�eZ)�;"���/3��՟���uڨ�e!}ہF_O�Dq�(�6͋�����K���4Zݎ,=wi�:s�v�4D�B�m�_/�̅���,_;�_ ����w���q7���;h���f���i��6De��q��#�\Xz'a��WZ7�S'�������	wR�X�j�|�6r(��&O�ݒڴ���8/�^���tf�(H���~3{^gm+ͤx�Ԏζ�;�uD�*�yEگ����UM��y���v���i�8vV F�Q}�%9$��u��Y����%b�-��b�-��b�-��b�-��b�-���6�E�#h�^@�I�PU���F�o�眢tu�h��%�:������Tp<�S��*:��i��S�'��6D4Qw��[�X���$�\��H�|�4c�ᱭ�U~}�`]���������]*I�!��ԅ��V�4����cߒ����-�픢p�.IӍ(����VT�YE���N���,WP�\i���(
Zsg�ӲY5������7�h�(J`6k�[����vGtR�h��v�)yn�$ܓ��ǿ����o�����>�Gv�i���AV�tO�:@��(:�5��A����x.!����|͆�M��g�#�w�yv,M)4��������=0���PN}�㝶�}?���ȳ���tͻ���
<���6��h��ڿ��@k+(���I���͔ym>��_��\�C�Ǒ]xd}T��z{�}�Di��O����[;��c��4E=�y�o��ģ�SC���3��K{$�kc%�2J}� &_'�x��h��k�G������_��P�&$�n�0<����r:�:����*HM%�K	�s�I2$QCB#0�G�	���-��ƾ�#4�l�2k�Dy<�EY����^~%J��mo��XC`��&���#L�D�/,��Y}l���˓|�]wF���y��V��~��
��f��V����B�Yf�^�qC�7i�͛w<d�}UQW��]���A#��"!��GT�a�9+`,H>�N�>�h�p�/��uN��R4���/yoW�9��0�����#�Dj<KJ-��z�H�L�eo}K�'�Is�Ot�D�����hH8�^���,<��Y�}k��p>9� qQ
�덌����r5��>.�A9���f@���G���{��`:f�qI��ݲ��i��Ҍ+I����@D�#�����	���P�͟O0���#h�&5�@4���u���Σa~R��F���=�
��1�ϵ#���Rv �;UN�:(l�dr"y�ׯp�����t��:\O���,庇�����w��>Q���Y�h��ռ��K�d7?������L�wb�x�|���V��5iS���mJϩ�n좹��4��U�����L`n�P�x�!ZoOdhR����湮�r�O��\vV;�������і�����i�p�>�?��q14��?�s���.�ƣt�/�"����~ډ��j��֙U=�O�\!��Kb��!*�X��p���DiW��>u&JW�V)�xޥ��5��v|i�x��	�āv�ϫ1�[l��[l��[l��[l��[lo ;�E�^(�7�IiX���D �,Q^���5uk��C���*4���m��g�&G��v�i��H�[�C��K��<��)w�B�0��ܢ���)�-O[���8ඈ�T�6I�d���f�P��ޜ�W���^�����ڕ+���i2�M}_�P���*�+ICF���<�m�x��N5=3���q�++Q
ɷ�dQ���]�������I����(����q����o�����s?�Ei�ML���bX_��es�dR4e�#K"�HOK�)h�դ5�ٔu�CV>[[�:OY��Hl5���Zi��eс�$_H
ɣ$1�B1���!æ���	����%
��}2���eH��I�~�ǋ蜻���T�xN�d��"�[��G�	��4s&5�!4崇�I凇oo�'�C.�0Z)��PӉ�)�����5kw}��.�vJ�M�K��|S�m5��������UN9��ŋOEi�k���G��(��c����F�hEd�@���:��}�V�Ψ_����x�hjҖa>rQ]�����L��i�(�=�Q�zB�v��
d3�E��Ei�Ѿ�2��B,��A�E9x���<�e<����! �D�r�Q�R�����8�y[���jD-#z)Z��(����y#�)w�yO�M�c�kw|O9��h��}+�'�y6JO)�g{Y��头%�d����g�2J��������&Jw5�о�j�u�g��Ƈ)�Q�]s�ʲ�N��iijͪ��+JyB��b��M9k�i�l�dC�B*XgD �QD�4H����,J�o��E=���Eۅ �([�C���R~C������Pt�L����g��]�1w|�*�A=�ny�Ο��NV�pK�Wu��rE��y����	���mD���/��qc�X�$~�O9�O��~}����];��u���ʇ��c��v��Ã��0}G��'�I�E�Δ�>�hrJ�����74�>�����D> P�4.�z6�@�����l���@jH���РY�qV�:)\��V4�ϭ�!$h�"n��8�G;�%^�FȾ@[x�>^#	?�h��4|y���|ubk���a7Լ>���yu}R+�W��������\�3�ٸ�k빐��"��u���/���S��������J4D��>��|Gc�h�U�(h����q��MB�}8�[�8R��9h��_wvl�4-�k�`��JX��C)Q�O�n�T@�1�0?CB;�U��9����� KtY�Y����v�f;�\�-�����N�U;2<�g�j�u|�:��������#'�:XZ;�%���x��.ؙ��:�Z@�_��G]�Ĳ`'l*�k":��I����.�9m�1낡��M�[l��[l��[l��[l��[l�m�E��{���RJ���IR�0�e���jJ:�s����^l�s���٬�M��	�Æ'��{h	�!5#Z`�qo^����U�әฤw\x_CM�ק�0��r���sza���;ܾ�����ْ�	mFyj�@Lb�.�8�8oJ��Mx�%�K���vo�3xP����g��7�d�vEin������oE�ٓe�}���(}�ɯ+v���Z�B�eD�ԥ�u�<0D���~�:Z�6��7�v���/G�v®��m�닜��3h��5#U��L�՜���ax���e��� M44��V4?+դ���@KOH����g�	Ab���7�M�n�iD�܄E�:v츝g���� ;9�~�g���!@��k��t��l��S���Wԯ��m[��*2�g*ӳ�nd\^,�u���)�<�կl��w�.(m��H<�Q��};�tw{[�dG���ɒ<]oW��5�8�ʖiF�V���(�e����b9E+�+ۣ������ݰr���OF�F��בXO�:/C��/�i�_��떏m����_{��hY/����i��������x��Ugf���\���k:vĈ���<�y�:����&�n\�q�D?KlZ�?bQ��.��6~ů-R�#�v>g�gO�ډ���%+�Mi�UW�K4�J<�u�+H9�)�WЎ����}�d8Φ�d����y~���FrҎ�Ԏ��+�74^���J�qn��wU�����c"�y�ߡ��g�O�MV��ӯٸ��[��M֖  ��IDAT�җ��h��I�2o����U�d?�}�멟T��Q^�d�{_�ADU�A��N^DaQ�� ��4c
�"z�V������<�H��W�,��PC�$�h:e�N��.�q��y�;�&�-��tE��4��߻�>�����>Q8e��*��?������_�z#�d>1������dȀ��B�I�D�Ps̏�My���_`���~�Qy7���mCH�L���|��V�҇vǺ�uΪ�n�5F��Cn�����Y�(k�v=����c!��5?��Fփ�
vI8�/}�����D2��h�rp܆�!���iej|��8�fXQ�jI��~��q]��������z��2��ﻨ�<���k�SP��d��^h�?��ѣ6^Q_�g�H���Ѩ�|���
	"�!�d<��h=3��ˁ�֐�g}�4ɒ���)P�v�$Bq,重#}C�g�sg�!.<�f!IN�QjM��3x�F�kɴwXKdUU��\|:J��"�!̂�&�Dv;&��>PS����zޯ��{��vsw[�v���k�����^��C^�x%c��լ�Oe���v���ǎ�AG�$gi�秬�g����I�]��k7�"���e�{�i�~�K[�nI�ҌuV���D���|�WD��NCOZ�����~���r>E���%hWO�h�����=ʃy����B.��\�AJ��G���!)�i���=;�Ҥ�%[��O���������6�8ϭ�'�N+�#�έ!A)����B1�[l��[l��[l��[l��[lo ��olʐ�#�S���<�1���k!azdj��c�G9�k��xI*x���?�w�#	��a������%�Ƙ#��G*&>�E=f��/�w!��9$�_���;�HP]O��V)O"N�A��	(���/5���S��Ӷ���W^��?�/��(��6�������#oz$J�@�l�]Z��}��iD}�3�SK�9ȕE��~^��//_��3w�uy��A��������*7����@P��vW�$m:h`�E�e*��>�:%��no�H�ꖕ�^[ѯ�D.ueY�:U}O����I��K�1��c�K����y��舴��}���[+�Zn�ݪ�9I���D�E��
j�!Q���[�Vf���t�fഴ%�~�/Y=�JK� �;4P��Q�"��ڛ{vޝ�=�JKQғE+�.�<�}�e鄈����bm?O4ZV?��Fv�iѧ�xܕfaM�pG�Z����ᗣ�����|=��=U�����#�)���X�O�[���R�e~XY7Bkn��qO=���E�{YD�f�f�������$Q>f�,�W���(�s����dD\^��<�����8�U?Ȥ��6E~LIS��:!-¾H�ڀ�w4o�G�y�1+R��bR�M�J��k��Y���Ɔ�o�?v��K�a����|7�=�R���o����������D��qq���Vޛ׭ߔ��Q=�������w�e�s�ƶ-훧�5����3Q�#���`�nY�9�E�}Q����_>J��[��'���Ҟ��4�'���s�q�[eRB" ���gT�U}��znlUU���!6���|hqe�g" zզ�C�EҒ�H���(�}y����o��!i�5_������7��l�`l���I���s�8%"yi�H��$����X4E5��
����OJS�'r�/��#C�O�9��l_d�d��fdm��Y�Ǥ�EU"�M�뉦�ǖ�P��Ϛ4��I[��U�R,���쩾�D�S�sv������/�5Y�6�?!?��y����¼��ū�XyZKS�Zm�>���DB��&��'=�;Z�sڱ����vL<��3v� �.D�����_32�� �����F�W?�Z7���=��Q��O>O��7E�����4<�}���ⲕ�K/A�rD뵄�g���Q��`�"3���J�ٗ�.+�~TRvh��UU�4n�=�g�E�Z^��۩1��k��A#��`�����Y�Re��B+K�Mo�"��$�k��{��se�h�M��GC�3 �z�u�}F9GTRY? �{���
�?�(��;"�w�V~^���i����IS�}���B�[�\�t��@L���K�j9���[f�U{�>����h��Vw؏�������ʹv�h]�67�I\�r�L8b�'ӆJ�EJj]	�}��ȇ`��q��uf���-���A��N�`��uQ��N �]�G˝ό�{y�Q��3��PKmB��{?��/$�64�2;N;�'�!�8ϐl��S���v ��}��5��\�8-D���݈�ph�����}��[l��[l��[l��[l����[~�2i^a;9N5��{̽>�o������s�z#�ߘ����&=5Fc/�o�q�HO�{�殣��B���hN������D�eh'�wp`�� ߈����.H�Ԉ���=���ֺyR?�_>��]�@.,���3������=]�˷�yDh�)�S8���hR��a�m�H��G����w�/J�������'M��]�{o�^�g��~�cQ���ע�"ͱ�����U����R�jh��Fãh��3Z,�'d�*2a^ui�\�����y �f̣�	<!xRp��1�X n{"�f��(�� ��M�1�����%�f.�Y�h�I�/��}F�v<ZME�<"-���P4�6��8Q��TJQ-5Ra��Hx~���i5�h�MTϦ��*"�zF�|�S=5�v\U����[i.m���m�����S�1ٷzɈ���%�+OZO��z��ZC�G���M�KH�j���)���(UX�Iif�!������8����E/�rA���u#�N����h�P��>h�|�?<�%hA6�R��}O(�j�i�{y��� RQQ��"^�L���(bcM�.�Ǧ���Ʊ���-��#��>7�8Q*K�Vb�(e	�(�BQ�Nh�ɈFMJ9���n�tV�]Kڎ��?�ҋ�`|ࡇ�������y.J��<>���������W;5�D��[~�>y��SF��Q����_��?��E�Ʋ��~�o���w����?E�]w����Di_�|C�QDow`��i7��#�l�4bܭ+�^]�Uș��O�U68س�<�̖94a���XWM��k��� K���ϝ�y��wMڡI�CA�����CYѿgJ6O�LHcv�<㗟�z�뼑����~:J�-�&_t5\�8M������g?�u������%��8��^UdK��O�D�MrW�ߜ�O4WY7B�2nA�1O0~A*��U�,��WDTA.]�b�����|	2�qAL"����^K�gu���f���T4K"�ܺ�i�&t���y i��vU�%�n6aY��r_ݒ&s�����/HҚ�5Ь�:Y�4ԿN���D���N��Vʊ��vޱ�=�����/D͍u#_��!�J*����4q��"^�Ӡ+�P��74��.Қ?!_�}�b*׺޼��"�\4� /ј�H��&�rj�/N�����aJ��AHҠ�U��qH��e�u!d���v0슈-����h���gӤ����u �k7����P�c��4�Т��Ӟ ����
41C���j���_�F�۬��>�97�Ő]�1�����"*n�K�]%�iN`<�*Xy�}δ�ϝ�y�~�:���kS��=�=�����7l��2D�@n�hM���l�޹o�GB�.��nK�(�����mLU�)�?��a`<��E86Sv�t���:�,����Q>��9�����0F�͞��o�6�����@Qi�f�#�����|�;���=�s&ч!���M����
Q�	v�5n��N�a�遗�P�-P�Iy0�:�K�ܒ����e�[v�`e�'x�Ŷ�����=�ov�voq�d"��b�-��b�-��b�-��b�-��b�+o���7$��7���`rmx��_��9�aQrÿ�Qn��\7$�0��ׁ����ҹ�ZxC��$��,(�D��0=�<���E�	4	��7k��!�Qa��8j�d����AX�b���eK���:2c�-O��D���O9p�Y#L�Ғ��c�ĩ{݃]<CBQ�H�L����a�����v���o�z�~÷�+J�����_���{�2m�{0r"/Oў�K%E��hPZ;,I[m<�Ey�����҄���ǥ$CG��޴<�8���bO'Q��ј�;�v�Ҽ�sxb����%�0��x5��%�1���$k��y&�댴t��W��"_�獸��W��<yʢ)�)���}O�=�8������@]�b�d�>y��"^�oX�m,)�p������*����<�hB�@q[\<�D]-��>7c���<WG��T���j����n�<��}�&-����JZ�D�#��<�����g��+�P&�5������}x�IC�d��}G��Ƴ��,-(i�M�Dڕ'9��0c�t�r���Y^A�^���Ȃ.d������&����ω���n5x����]%,Ц��eI$ڞ򻨨��?AY��fu+��4�.�|)J����Q�t���z8J�����ҹ	�����Ҍ��.��nG�L�5[A�����K/E)�[��ei�������>j��?�o�M���o�7����v�=mZ_>a�`�e���q����#���5x
y?j�3"eZ{���-�Ͽ�;O��f �쌰�����qoRx�+��ƺ��?W�F�����S6Nlt?"�J�x|�1�o���?�w�v>Js�^^K�4ddA@t3ޗDr��N�7�Q��'?������o3�w���bAQ��vH�v�+b���~W$�Ҍ��+�4���6�ȏ��C{��
w(���y��F'��E���ȑ:jD�f~���$�5�'dB*�\�Ni[��D�������yrC�ʻ��S�_��yKF]��1Zt2Ss"���ۡ ��}�1d`{���"��kV�k"A�:��N����H�"�!���?h�-r3������)����|�:�@���Hʭ�y�r�,��Fk�H�Mi/C�Q�����-����6��y���űSډ�y�u Q�!ֺ"Z��2Dc�(�׾Hx�����HE�iC�k�������[g��Nh��`vD�\v$���:3'�
������W������[/����:
"�PԸC4f�k�����cG���t�(=����ַG�)=Oe0:hW���\��g_���F�?z���O\�眯<��GB|�nw��~sD�4%k��3z�,)znQ�ڹA?��������)��"��Zoe���hJ�P�^�(mm5���!!��7�hK����(������i-57��#�v8�ѧi?��Yw�;��?�Ot|a��\D۴)r�߱^%�h�r?h�����v����h���`�Gyn_X02y[ڒ�7���A0o2^�=���H9&|I>�y;���v���&g��[l��[l��[l��[l��[lo|ˌ�� Bɐ�
�>�c�Ά�ܭ~Cu��Y�	���E��a�'��<�ej����E:�F߸#��l�������D��I=�h�z����x�A%W.cN I�u�c��lOdK!i������w~O�>�)#C����|?�S?J�I{��e��� �����'������i�q��Mo��F����TJ��Ⱦ��F�|��L{������s��F�Ҵ���>S�@QtT��(/<xTrx��h��q�iy�J����Y)+O�j
-<�ui�q]<)x \TEiU����q)��wV�E&O+DiMyڜ���Kso�s)7!O޶<�yE�Dۨ�
<(���uEQ��"��F�=i���l�։���ܓǨH�2�۠k�_q�Wq�����q����F�{����WL�,��λ����^L��0g�9s�<����JOn� Y���ŋ��E��<w�m�]@n6E�P�DguZ��E/�A��ES}�ӶL+js_��DZ%i]�����eW£���pEZY}GBA��E-e|�;��/�h�X-GEi��s�ȥ뛦�W{�?��Q-AF��1�4�T x>��;�y��VW����#'���Hs0��ϣ ��NW[��E� +:[:E{��~��	}�v��ǌ������(}F���ߵ�����[�������;��]�o�a���t�����*���\�.vet��1݇��#?��Q������k�v���pB���c��������(}���Y�mib�8?�(���G;�BsV��d��u$ڢl�������i�e�(�{��� ��)�њ++��ޚ�_�9%�i��3�FL-�d��g��oy�����n��m�Z_�Id�e�F$D�#�4?��"����w=�(}�^�|��_�?�t}����]�1�U}��r"�Z�������!�Цʤm�����慣���O�O�ͤiE��~����SF�C��w\������͉��s��D��ܴ|D>mJ㳤��G��������!$ɩ�c�� ���i�so��?��H�[�6n�Sf��C��ɵ�Uݯ�dڦ�Z��#y�c��hB Q_��h�j~#�vO;U��j�O?�T���m�.�7��D~��v^�}�khcnm����P�!.RRM=�V���� ����45?CC^R�S�C��u�J�rʹ#��fVD�J���G#mw[�%�N�_rM��aZ�UO�7HƵ��1�9�sфu��w�w!O1�S�VU�O�fCT_�g�\��������Za:u��gNd�MZ����+M⹒���b���ϞG�Ca����Ħ��,�P��)K*"���4Y���_��߰��t�I������U���c��4�Y�$|���1�������)�%M�1Qv��5�]"����x�g]ѬӖ�\����I�.��h��ϴ�c�Ţ��r;�����0Gz�g�=�ۄ��z\�Qj��=Ok~�4������m=��|  !2A�q��F}i�3�65��E|<��Ŋ�5��y1+���\6��_]�84���|)�~�V��0�K%�"}��[l��[l��[l��[l�����}�<�W�)�P~��4���;� ;�F���w]w���|�W�b��'���&v�1�H�d��_ϝ/9&�E�/� ��=�}��E�d�����3\�����9\��h���mQ���/E��|��!�f������Z|BGD.Av����O��4��%ؔG�!Үط�g����ed߳ϚF�K˯D�g?��(�St�O��ǣ����OE������DƠ��Vмȍ��'�xD�f\B�D���y*�=;�5�^]�bdd��]xz��\��ܓ&�8�R_��s'�$CC���NSN��<f�C�d���sV�/_~ѻޔ���D���Q9o��O7��ڲ��;�hc[V��"9-��^��vİ�YE��0h��d<���
!���h^xɈ����vDP�U�E$�ܠ-ĸ.OWVI4�����Թ3�oy7_2M��I+��|Ԣ���F��a�$�5/���O}]P�9��C4D����I��5ieA�@�BB�ѽ�j$0���<���c^Q�!��츱���/�y�͞���"[��U5bijjZ׵�ATD��1�I�ov�(�v���W��f`:#�u����m���x�S���P��\3B�Mo3��b�����n�ҫ�\�ғ�Z�!�蛅��（�\VQO�v���?��Q��È�_�E#��5N�=f������~��WW^��C
L�ӽ)ҧ%�jG�Qi{N�@[P��$Y\��]W��ǭ�����(�'�����q��c�=�r��'�4J��~]��3/m�?� �y�E<����Fx�8@x���%�^��cOd��+F�A��uD{bxe�uQ��:mߣ��8�Vأ��ė-��ٓ�^��}F�m^�~IԹ2�Ԫ��<��De�����ߎ�q���d��8��/@w��c�������[��DWtϺ�UǴ�����4ZER�h�vT���?�Q�3�~BZ�DK��}��6/R�q �ꁇ-Z�3O�ڏ�sC;\�M�Sq�[�x�	q���w OO!����B1?E}E�����5���;��� d�����x��V4�������mw�%�3D#��].��D�@~dn������@jB�L�ڸ9�?�{h�v�"r K��O �
قA�좡��)e�B�M�5�Q�,���ycb�׶�,D�(�D��<���[�[~ Q!�јD�֙k&�z�v�z���T�id��z����K��
��Bn:=�� �k~?�-wi�	�n�_�%��1Z��O�}벍K?��F�1���.�v�'K!���vޡ�@2U��7M���o��(�؟�zqW뱅����h Y�I�;x/A&�9�h�����/�+�GGojO�ܓ��4�Y/�k�f����T���h�g4&Ѣcb�ω<v���d%�0��c4�B0��V;�x�`�#s��d���N+�E�{�Y��uJU���%�ŭ~:9�'����Ϫ�;����~:#������/1����iH4�w��T�8��ؒ�3T�~}}��[l��[l��[l��[l�����Qw���8�G�B��_%���N�����]'��9:ȏ{S�z�^�%�^�F=���8r�v0��1�?�����G������qI���y�y�ޕ���]����Ƚ?��OD��9#����y��x�\1���V����k���5�����z?%2滿�Q�淼%J���v�!�!�Q0Ɔ���������ҥ��ɟ���6�x�#Y�f3���<3�����<W�@�v�L�~��F--�-E�]X�Wy��<��g���P���'�V��{��5�j�nZ��㑷E��5Ӗ�����ue7#� Ay�r��v�ݝ�6�iQ���	yX�~BS��Y#��^���6�͆���@����!�deQ�>�^����x�E+���V��SF�<��iG�A�u��ǫѷ�Y��	؝�YTɯ�{�wQ�\[�(������G�G�MAy�4�Oȍ�$'Ф9uʏʖ�23e��S���T4b��>Z��N���Ԥ]��뢵����zDKeUDڀ�C45O�1�Ӷ/R���sgL�kn����Y.������i��~�ӟ�r��2'�,�<�0�R��C��"��Ƴ�^~!X!	�"�h)������gl�;y�L��t�ℵ�I�g�/[{hUm|�]�e��OX4�)EI�[��w!�D��N^y�e�zy�K����f��m���{��O<�O}��Q��8J��}�~��l<�j�NיQ=OB������Z}|�c��K���v��sA����M���׈��_�k����zo�~��������(��_��Q����7J��l����8J��=ߡ�g_Q���
گY9tV��y���x� �vK��u�8+�h���E��'}��q{J��wj"���H�/~�Q���S����oU��?�韉R�ZX3"�����n��Ɔ����/J_x�b��D0�]��d��7�E�_����-ߦj��z!�y�{�k������һ�l�!E�ǾO��Q�Ɛ��ֶ��2R�8h.A@B��ğ#R4^�TOժ'��c���P�:�ǑHiE���x���ꬫ�ZK=�e�|��e�Z�3o������SRQ:��Ұ�!��z���4W�?�W���C��|N�"�Q8�	Dye\sQ/���-E�E��i5+�"�!P8���]w���HӎH�.�:M��y��._��PV��NCXe2m�/�nG�Z{����=Z?@���Ƣ�Ƹ��#�=�;��!�14����톴�EP��v�W&��|��[�;*g4��_��$$iHn�~[�ܳ�s�5���ߑu	w4��4|���$QN��v:u;���<khA��O
:� j4��y��Eͦ��n�_;UN/.y����K��Gc�['��M��NrK�U��۵�Zy]�f���������-Q��m�}u����8w4�N�z?���]yh�C����o45�%\;8��s�f">;�眕�~}������N���Ɇ�mJ�Y=7��;~�G�Y������q;�X�N����"�)�P���SN3T�=ż7`]���0�`l����H=O*��������W�oG꩝�����B���+�1��{B�E�UK���y}��[l��[l��[l��[l�������4���n@X�=��մ�������u��4��Hr��.^7�7Εt��_�F�qȕ�!D%�����ى�X�K@�%z�V��[�ڕg.E�����[~G�ANsm�<ƿ�[��_��E�D[��@��Z���_��(����Ļ���(}�o��,煂<� �=f��o�������mmN�e�kF6Y4�/|�"� ��E�#���(�y�"t ���AIQ���F���,�h(��D�����0k�K�ųn3~�їiQV�Ү<�]�)D�9�h}hk�;�����	#'fJ�PT=�DT�v�D�k�#L9.3����gR�f��5i�MV���˳��_�b�jB�%��>���G)dЖ����q]�ǿ!O��3g,���?i���]��y#�J��vV�S]E�D�:�*�XW;��Y;�e�Աz>}��|ٴ'E6^���4��D.^�3#��}�c���Gi��wA�(�9H��S���GTF����oH��	O ��.M��4�^T�N�<k�-`q�H�)E�k���A47��sy�A��VD,N&E$H�cn��#��[V�x�Ϩ�פ�F��D��:m��+��E�S�p�����7g���3ߛ��S��7��s"��T/�`����u�v�u���U�OY�~A�J�h�5���k<8�d�άη#2�i�I#�4m~��C�~�Fn�3%��?��������>���/���{�h��G>b��h������|Ĵ�>���{7,�o��wF��i��3F,����v�9�)��"b_�Ҭ�/&<�m-���n�O����.�xC�C(ϋ��5Qx�J2@��ԏ� uO��غb���{��*j�DA��H� "������M�_��Ж���g��V�k"��G�v�>��i>���k�p 6N/Z{��iO�E��k^C������y�K"��B+�7���?z#$$SMDD"Z=�!D_[��xrگy� ��!���j��>��Ww��{�e$��gD�V�����'Z�y�'u�Wc۾�����䓦y��(��V^�h�%���w��k�5?�фV)���^�E�<x��]z�4!YoBhP��K�G�py�Ʊ�v
}���_|̢N����!�Zu�N�R�Y�<��xh�A���� �^��h fE��=��N�q�c^���/�z�?Q_Dy�]���D��J;��!Z��f�`���N�4\ݰy}�����ڐi]�YEK��Ƌ��h��Z_�ad��w7�39V��iW�Z�S/�w���J�5 !.ER�����״;��v$w�<h���#D����Y?���m��[�O���q]VC���u��h��X�|���z�>��s���'O��
�ײƟB-h�~�;l~��O2JgO�����iH�Yʓt}��9��h�Ss6�B���j����U#|Z N�M����X�s[ʏZ��u/��?$F�-PO��i��{n�q݌ӊ3k��Jh��~վ6�N���$MJH>��Ḫ��֩h������x�-蹉�f���u?��Z?�;�\+�J�gw}�E�_I�ʺU�c���h$b��4t��s]�Dyv$d��,&�b�-��b�-��b�-��b�-��b��`�5�x�{|�S� ��X���}��v��α1�5��k��s��s������C�;�8|���q�{rp����0�����7��z���l��>�fc�����H#2�{��2Bc����I�E�3'm���̓���=}\��o���D�S�Xt�xL!�2�P�e(Da��_�U��D��"��P4O怨E"�>�?�?�?Y��(ns�fx�i�<��E���xf\���\ ��@$��z���ˬ<�;��S>k���M�-��h]i���S����s7��öy� �
� }�Zi+j.�gZ�?h8���RN�/ h9<U�W&g����!
&oGf������r�<��[��e��FU�>hƬC2�O��Y;﮴�**�4�V�9���v�6%��3F�\�<�h��f̣Z��޵ߝX��D)#z�<fD���<[-^f'N��vVh)i�5E�V�靓'v�<�"֮�Y9..�:1%�E�IF���r�·���;�42���']��sF\�Yޯ<s5�ߔ<�D�l�rV-y{my3�ʑF��~��JK�����L#.� �<���94���� ���M�TGȪ}�4ϊԫ��ߐ&P[Q~�^��Y�Wq��I]��o���oׅ�J:�M��+�G)'��Y��Mi5��?��(��o4�yU�[���\?���A�BVM�Z?�Y�)r�|Ď[Q�L����e�.Aب=fRD�����׌4���O���~�磔�ZV�����}آ����ܢ��vk���&�*V�w�!;���ȇ�v�Q6̯����{ 
���"��E��v���QӚr�7�wD:��'�8Q7V�n?g���i�i}��������Ҭ|��M����h����Qk'��n^q����:bW����oLK�'~����>kQhzд6�h͈��Fi���W>��YE�)���`�J�阈�Et{GC�΂H������!��l�1���;��h���I�C��I;�-�z�	�����{�I�Ҳ�8����d
�h�sT���3w[���5k'Y�[�_fE��̆4�Xc�Hí+m>�R��)#�]4�@k	£�q{W��I�X �9�Ԣ�Q��4~������Qmvd3롲�T�Ǝ�����O�|�����mu���Һ\	:ϼ��=;��V?DK�xw�v�>N���S9N�p	T4>�:t;O47ETe�V�1p�����L����?�򓖟Ȯ��s���ʋ�^+��Qy��3Q�_��s����Һ��nG�q��H�72�vjB����%�k�N�fgD��<���1�$�	Ĕv�@�
��<n�}V�w?������~
1�փگ���_����y�f�ϱ���=p�ާ��s����g��ME�=�qd�"�S���#� �z������;-�<P>Ш%�}K�";����������2ڡ�!*��G�c{��Q�q@�Y[Z߰��E�V=��>�I�pG��W�"i]�w����N<����������F�%�	��E�V;��}2�B�A��	�q�l4^�;b�w`ǚ#�E ��m5�����bv
����!(7o*0;����������w2�=�����y�]�]���-�M)���J������x_�l�鉠1KCC�x��1=3��l���K�01��Y��l0c6xߪ�]�JRIJ)����_������s^^e�������CG��}��{�{������{�O����"�-Z�hѢE�-Z�hѢE�-���'� ��>w�7ۇk�=7͸��|#�C����7�,ȺN>Є�����zG�����,���ddM:����9��u80p�g Ҁ��"z�u���������@�b�`NS��{cRZd�6���$�zUkà����ߟ��>�X��m�&2-�0�]h{�C���W��{���7їǓ�s]+��9�D�9iZf׶��y�ސ��K�r�ز� x�l��+�����"R ��`k�sU۾�.�`�0�)k�,C�@��(�����0�;g�MтA���͑�h�#�8�/�7��3"R�bN�����a���E#�GP)�gM���2��i�aj�#��b�	A9���k���g�"� �4��O<��(x���Y�簨(}EM�e�����w_��%Rb�h�9�+�J�z"��j9)��U~"	��B�>�(�s��]��R;,�)A���%)�����1&BI�QȨ˗��X��d�����'l�8w���=��
�F�i"��ooI�eB��Q��m���	&J밆�ݏr��7�'�h��hB��PQ�k�[EZiRuzv�޾����}�5ٔfI_�Ah��T�SU;o^Ԇ���0ͺ���{�r�ğ}D��淪��r�|ň�i��?������sK:>���f���cUZ6��%�g~�g�������| 5���������(�s'�����o���O�y����AS��g~O$Ӿ�",��^�L/���!7B��77|� $���Q=;=�J{"*���3�@���w�*������E�=>c�ڢ�J�yԷUS���]��1�s�Vr�`�p����w�3I�'������G�*���ޛ���+#��?V֬%pB�S���l}�G�m�G�"��֝�z�N ���O?��`��H�fj\!�������F��k��W�#Bb������D�k� �pޟ�Ӡ�J���Hǚ�B�Dǉ���<����k~��Ѷz�����5#��E��X�A@�)
9�ѣ��	燸pQ)OE��0Ķ�=����e7���9�ň��Zg0��*"�wm}0.M`���u��<�hO]��h
2�4��9����Q^�Ꮀ�@���5�^g'g��[{�^��7�����������5����^����Q�Z���e���}�J���S�C!I�v�$�|JNi�c"�z�����0߻u���](U9!h�s�)[�w��<� .k�dGѴ��_�ȿ��k�uL�p_;���s���X?��O'�5=��猞�����u�=Z/|�ˏz�m����<�@��|-���@C�(��i�$�>"�G����He�Ӗ�%�%�ӳ�CS�In�H`4�ѧ�R��*W<��!����: �_�M)­t��g����Z�j\��x�}B�Q�NCx蟗��3k�;�O�+�r�H?b\�����s_��_֏.ր�ۢ�}mA��s��7T�ż���ck�o�敶�p����D_�hѢE�-Z�hѢE�-Z�h�;� }	S�A��;$z��&_f�B�.C[.��0_�݊9�(�(u�A͐лu��E������}TB�i�ȃ#6�����r)�rwx8���I7��	/s0A���=JSn�<����rN��Æ4�N<bd��h��o���П��wWo���fVx��剧���z�ޔ�����T�Cpr��Ⱥޮ�Z���y�7���۔fX��ڑ<{{v\���q_�"�M+K�n�hz��������OL]�TU�f�<Sx��]Q��
�)g<�S��#jl��
�L��k�}���wѓ���#�0��V;���wY�t!REk����/[T�{�5��֮�}FZj�.���`�� Ѯ6D�8-y��my����rر�e�_�]�Ӧ�V��aR��z"f7U�}�G�o�Ѱ~�ٳ�a�&��w�ݔ4/_1�-�Uᙆ蜔�������z$��<�"���Ex6����ui�}�8���a�&Ȏ<����G>4��*��"�����ey(ъQ=um�X�h�f�+<�9�DUs� �U9]�FVcBZ/�R�Gz�6�ʣ#��$r�,rʑ&�O\���qD���Ad�WE4+�ug�ޅ��8#���4.f���u���gD��-�O~��I��h���������4�������%��ےtj܈ƹJ�����[�޿��}��>k����؅d�b{.*���.�-i���p�|�f߽����#�k���o ��Ho�U;m'����}�M4B��(S�C͊`'ztGD�}��xW0΢���ҋ/$)�7��G5]�g�ؘ!O��?����[���$m���y�d�uN�Ds��T"j#��n��G���" \!�#�XNA�C��!|��u�-?h�B��T̷h�,��iF�#_��2;cԎ�>�1�A ��˟څ�挶�滪�$y�ق���i�'�(gw~��7Ђ�|A���v�,,,x���q��!�\�{�i�)J�ͻ�fԖ�wЂS���E���#Eލ�����9����.���	�QeѼB#�h�����|f��C�#�B��i�d\�r�j���w��y���hZ?��_��G5�sD�������uF�'� ��$��Z��>*�����s��s�H-u��SXސy�T����8j���g�^�h�/8s��K��"�75�@v���Z�6�}�֎��*&G02?�1�h�H C��S���FW�<WQx�ԙ$��Ӧ��s�I����z����+ׅS�Y�:pR���j�9��E}����NH�ޫ}z+o���j��9mW;hІf�7��&D&������)��?�*x���K�h��ћi����=��&͇ՊO�BB;miU����yR�����j+��sZ�?�Z��%��2��_ߍ�Z/A����[��������3�D�v;�D�b��Q_#E�/Z�hѢE�-Z�hѢE�-Z��e���c4���j�=��������I��=ߣB��-����$�8/�dY7� ��{��|8�o4���|�r�',��C�|���)��~L�K���0�?rوDX:iZa7�H�iyʗ/����c�:�������(]xT8�VSĮ��0s����,(��"�>��E=q��
Y�|��l*�����������!OrA�TW4���l�сt�����=y��!���h�a,��g�EcR���]��u�BO��}�/y�S� 3<;hL�ZB'x@e�C�V��!�5)����<�D���ў0����y�M���-og��~w]�\���(hm�}դ!wr�4�楁��f睟��lKK�hN�U�DY�HT�(�Ͷ�.�焈�Ui0n��]��'�!CQ�%O��E�ߚ~w�m�=��-�Y�D�P��	E�C��-HZ��Ix��ת~�jM��MRO'���
�p��ȧ?��?���v�آ�@�AFw�YĳITż��>��6��<���<��vĵ���?�ݛr$E3�&�p_י���4;f��Uk�'�߬�H|۷}��/�W���ӟ!�nuv�����";��.<��/�ߢ�t�n��@Ɖ��D������b�z!ܖ��F�"
T�h�U�P=�;-t4<77Uq�@d�h�h6�E����kG�i�B���o�F�o���#!,ׯ�8�0��Կ��D!1g)� ZV�Դ�����9I!V�~��F ~�QӐ����/�1]�r�@�h z���Ț�@?x��%�p}Q � Y�|���xj>�ј�}brjO�ڈ]����w�a�h�ME�WYɡ�*RC�Z�[��虌��E��"���V��v:"{N�x��y�$�go7B�b��D�����!�.Qk���TX��.vE��.Ѻ\I��`��*
1ZO~�w�<��a��SS��p�Vv�@�q�"�����(7HC��i�~(/G���d���"��͐�[��=Q���o�M&RZ���3��yͭ��͌r����ʇq������i	�_�[��z���[�I����)$���KݮO�i���/;lJҀ��P9CHr5���W��颴/���4DdJ��pj龫�h*s�u���c�.�DZw'�~�Ej3��#h����)�����
2rF�yn�'�ٹS)@��\@������c�u �q���E�z���sj��D6;��3z^�P�x��N?U}@�~d��1�� ��N@:z�j��;��gZ-�Ṑ���WZo�����@�� ���;l�����K4l�ggDߩS�|}]��'ϳ�2�Ե�f�K��B-�r���O���qQ�)�����묬���hѢE�-Z�hѢE�-Z�hўv�/�2��{��9 �B����9m���<W{���Si�Y��6G�� ���!ȨC�6��N#��!�B2$�\����4C��m�exv �7Dy��hS�h�"G�	�+�_o�<&�~��I��n�Ar�;���|J�Lo���*�����D�O:���e�mI{�3����I_ߑ���b��C:��������{�	��v��('���y@u���!������3V���Bs�VF�˅9�Z8sҚ�xv�?!�[G��d����C��F�	�o�Q� ��;��<�NSH�!�lN�d��G��h�u�	��j�ړ�	���_��I��O�2%����4CZ��[�>����H�9��h�u�Dy�NI��m��Ĺ�F�]�t��'bBcF�Ʌv��[<�w�iZZ�V��:"�.���P�r�Ǒz�_>�i���Z�vv���æ�ie�8fd�~��1.�aLZ ���v�l�>�D&��#gԏ��GK���|��v��-���x�Y$&Ѥy?*YUR��Y�U5%i��58���U*�M���c�$�����}%�ុ���E|N�q�����:��k# 5!C���~����_��sM��8d�p��#.�Y�ٖ�g> �Ҩ�h��T�|�:cd��e�n�h���L$��k�F�h�NIN�v�7�I!\0G�|-�Mi����E>�?:�D+��V���Ǻhp��b� �^�����j�Ds�2�A�i��L�M���"�"�R�b��|�����"M����"�1�o�����pQQ!�4~���
���l�\׸ I3�6�l7������T���m�-i�4���ztw�נt�Q�i��>��E���a?Ц�,�O�m�*��]�E��:i�|ۍc>IuE�9�AQ�At[��+��w������\�ߝx�I�:�/�Z������cYSA$7d:���J��d���=/B���<����D�E�D����9�v����C��whS�n�$$YX`��$�4;c��~���G��)�٤�)�%+'���7����T���]���io*���)d��6�oo����,�P�u�5NT�C��-�C!��Z*e�ғsK����zz���7��`>���@i�W+����1��q�*"}���)i��F\ϟ��xN��Z�I��
v�>���6�����X'�|}@�ܖftU��)o��X��\�ovu���:�v��<�!�y���F\t���DIf�wQ|��Ƹ����~����?�=�z��٩U�����h��aż���0���s��rb>d�_Y]񮿯z@�?�hF�E;��Nwp���z�Wq�Qŀ����uW�E�/Z�hѢE�-Z�hѢE�-Z�灍��K��g�z��>�L9$
�-G���!�7�� _�����~�'���5u7 �F���d͉ �Ǐ^���y<�Ywp���>8�o������EW;����n���S+�BD��M{�����nY1O�l�<0��ȥ���G6<��7�Њ��T��F��π8u���I�OZ�e4�uE_�Zڊ�S�g�P���]Q����d�\��ݗ��D�bK
�����-��)y&���M�/�4��D+�� j�<h����6�뗺�����L��9�*��+�g��j�m�a���6Z)�[�a�#4I��"77ϱ�u�v�}]�����D��NO�՞�>$d׊�>#���/?jڎS�vE�)y&gO����������<�k+��2l��y#T�f=��V�"�p���m,�*�^v���3���C��"�%���՞��0���O|��E�=�9�h�v��E�ݪ�,��	��9��ø�2��ĢOj�D]����X�@k����G(�Ů�G�F����۪<�xʻ�;�߾�L����f��Q�xT�'�.'ѕ{;����s�g�}<�e��!����v���(~�fK{���E�>�z���C���#_�H���}��h%aY�jh�_!�D��$ږg�� B���3���!�N��h����t}�";8o��V�o�ANc�y�	-bt��/`�_84a��5��4!�D���Xv��;��|A�о��(��5��<u��wǾ��j�ᄢ��N��ŵk֍��Z��aخ�y(��}��&馋���/�G�-���`�����ճ��9�?G,���ծ�Hxv���6�����YtRZA�*G�:�1�?�Z��J!� ��_�q����/>��m�h��c���,P�"����}tE��;hQ�$��Z��g6!�w�i�UxOZt�%E�q��wd��}�uE���#z%�(�Ⱥ�O�3�Y��pZ�/�����xS�zkW;�a@td��4YV���N�MR��ܺ��I�.�11��U>)2�4� D��)��X����T>'R���g����G���Ŝ�E]�Aв��Ǘ/�x��d_�B4+�@�n�:�ʽ>�1y�X�=p]�}���s���-��*�p�t���E]�跴��#��)&bvj��EmG� R�����d���?�P��%%���>i�xSA�6Ĩ��E�f���sU���z��`�^y� 1T��|�z�u v�����vEv~��|B��1i	�U_�O������k���Md�΍u�nK�)v��㢤��F�f�rv.Q�`����8����������c�t[�הc}�v��]����*�p��>�t{<���r�]��|���6;����-�g<�a���^�v������N)ʻ&�f4�Nv�����v�1^��@�?��[��9�@xǻ�3}���H�E�-Z�hѢE�-Z�hѢE��<�^��T�OU�koD�vͳ���i}ȓS
��\@4�� q���A�AH���#O�g_pW�u���sx#��Ͷ��:u5�Z�]���x��B}2��]7�6Fû�7M��� �x�v��|_�x k����L������CH:�5�~O�^k��q���
��Q��7������+��E��ܛ�'��Yi���vT2�0Cエ�xF�Ψ��@�@6�f�}���8���}ޓ'�Mt ��т �V��&Zzjf�	iџ��W���<$*�hHx6�gLc��%i�-(�(Z`��ڃ##!���
�2��K4#y<W�D�9�B���\��)\RM�� �v�&��6�v09e��.+4��U잻�p�X�re��-"a����C��A�<<>C9 h��������+n��O�5�=��'���K��x��h�h�������h*�| (�Q��v�1T<��O��k3At9����h�X�g����K.�L��#BiC��dO���7&���5/�i��w���g�=���>k�Ԓ�s7��}�)��P�	�A֓G�hn�o,�E��mE#t��@6�5h@��S��}��2�h��A	�${݇<���G���36���_N�-֧Ux�]�Ҹw��9�?�?w�@YU�:|����/�#�`�_c���O�OR�f�Ͱw���V~�����c3ʯ�+�'������m>�	�Y�55� �r^
�E��`׻k������k���Q�z��+��h�����^eo' LB�.���]����>�GZ�<����yYW}�۾û�,���W�u���H�]�9�;[�֛ ��I_ۉ赐b�� |Vڥ�g_������Hݎ4�zv}G�B�i�i�|���eǙG��D�M����N��D�m�R.�4o7�G=%z)d��G����8rA�k�hmA��4��4~��Lg1V
��R�K'���["�{��d���L)J0���~��K�����#�\ �u�u�4S�$q�lBK�P��Ę��vF?`�b]�z��$YQ�S`>f�t��/�脤�u���R�Y�����|��M=Տ
_�
B	҈�׮N��vX?k]��o�v��_����N����M�����W;��NNN�zv�|����h���*��pC]�\;`z��r�y��R,�%!�+AT�Ӯӷy�����[!o��4ֿAN }���O��}�]%J�ʭ$�<��7��%�q�O��\��MӰ�臌c{E�9��B;C+}���j����4��Q���/���|1n���_�Y8_B�Q���@$?�/�HG�:-O�}O{BӖ�΁�9�rR;�y�m��qƎC2����=��ovX�DwZ�:?哾��w�u�C��6�2Qʵ^q�~x@�������s���o1�E$��E�-Z�hѢE�-Z�hѢE{X)�t�	����s�)�O�y�_��7��.j,�>�,�a����E��(�O��fY����SI�/�xM��Ϝ�
 |�j�)WA��a����a}����K�}��:���~��MC��ܣó�ǌ���Q_�+ϛ���>uDz\�h����\����N�mD䔢=9�o��1#�q�;���,���� y
�h��qW���\x�H�)E�9>g��P��1iZ͌���3i���g-J�W=�P�~��Lҷ��Mv~i+]o G����$��_��$]:���aі��Ӛ�7h`L�CF=k��wQD�o�S���5�K�k-Z��<t�&A�CD����A[�%�x��O�<]�%;�ܤ��6ݰ��.���#C{�cJ$Ѡ��]��-O�*�Z�fL�G�/OQ��	]�Y�_ʽM+��	EMt$�H�-+��1�<Ë�LC�(N-�Պ4��k�Dh*�&�і��M�I�BQ�*y���yk����g媴���Q-�}'O�����13a�.�Xn�~5�vz嚑�*��M��}E���T8N�7�E����k���Cy��}�T��-c��c*'��%�����D�ڱ��Տ+i2?#Rl���.�y��zUZ��,���r&�־��씑�m��=wF�ɞ�so���v��ל�#%�����K"����#��}��E�7������^i(_x������G����B��{��93i�ay�Va�a��=&22�kJ��ڞ]�#͵	�K�5iF�]��SP}�:V��WE�.����	����$����O�_~ׯ%�O�������C 	_�b#J�\�:-˛{�1<��-Z��}���}F��y�%��G��#I�|U�>��'��Qqj���5�'�_����z����k�S�/�Y�ݸ&M��j�]���E�@ix��v�{���.���C���Љ��Ut�]�X���FOA�znI+wjR�Ȓ)�����g���/��w���8g����]������ Ő�|K�Zch�1޼��&)ш������7��A�eRڝ;[D��س�b�~?�|���fR����VN{�6>�:iD�������'z�������Z�ķzI��嵳�Q�v��Q�U^D��p�%՞F�;�O��"L�wٹb�&M[�g����O���֖��z����6�Ԫ6^1����֥M(��!�GM�֍�ʄw���������貊N?���!���S�v�&ż��<�k��k�-�/~H��!�A������:� ��h������ 5���ǻ�]+�fӏ�{邵����A�B��i�]8��ϊz)RiW�z�`�MNY�[]�yy^�]��x��z��Dƪ]�$<�vu�+67��d|�������QEY��GCݧW�������jE��Z�B(��D���T��8iX�&n�9�F]�;��a�*���V,Q��i)Y�u��c�=�[{y��3I������+=�i���o��$�����&�j8B��Q;HSd�ʅ�X򉷒���~�����^��޻1;������STgV�i���m�h������T!}mϪ�E�c�%�� (���gںv¤�|"LU�<�e��j����C��ۙ���������x��gl� �0��m��2����5�X��7D��e<G3>a���!!�p���BQ�:;��	Dy�=мL�bʍ��� _��BB�E���d��d�<Y��>÷FX$��E�-Z�hѢE�-Z�hѢE{Xi���\dx�f���R,h/uQ$�<�����a���P,�1�2�J<0��K����{�D���o����7���go��@pW�P����ʷO�G�m�iȳ �0=!�KQ�c�y|\�H�{s���	�' ��qQ� ��h�)��ȓwܙ�h�oB#nsW����Ј���F$~������u��y!�m1��������/�7�D�|���'���%/��y���-?���'��������u_��h����7���'O�{��V�h6���^E֙څ<�x`_�����jWE������c$ˋt�/y�˓tK�'n;���I�~x�>��?���<�e�`<���I:�(]y�'�!٫�z't�\�wj�`�p���"x�!Y�bX,��R?�紑]N�:�fD�.,�q����B��^������<U5�<�X�l�0�p����u�����(^h(�Q��*�1��������<�hY,�r�R�k��Lȳ���o�ӟ������yL�r���-��	R�k��]����F.BXVk�ώ+Jj��{�jo�I���ж�ޘ�!7�����Uij�Ox����/�ey8��h��W>��H���c�����4H%28�#�.��T��QT@�)ren����5�y�z9�"Nw�h^�XH��O��9D�-��*;z����p���Q�-�/���E�=�������ߖ�UnI�w<�x�s=������*�(Cä.�cf��oW��6���F���Vߚ����B4ϟ�ɟJ��j�~��/�}��{>SR_�4h�,3�ꕯJ�Yy�!^� }�Y��,_�N�|��'��n�н~�%6$�rV�c��\��.�"����=y��C�>�����Oc>q�����Oj�E�^]1Ҳ+��4ן�|�{���Xш9���e[�lI�oNQe�kv<�}�kv��W�h*��,*
/�Û5?o��y���N�B2�ZD�Â���嫶�x�ˌ |���n�� DG�i'��_Y~4ϣ��P�r��C���|���+�	�a���Y�S/���*Ϲ)�}ii�{6nw����v�[��}n����S&�ZK$��e�v�_�kT@��h�Y[y�}:/rm�e�!!'?sU4-�Ҭ��d��mX?X�fdYZ{�tc"ٯ\��3�`�p}��9_�v�a>�pF�v��|\��UES>q�擩iia9MX�����	�n|����u�A�!�F����pS�S�ŚHj�{+�v_L}'����GH,�uG��	�#dI���4[!�|� �XT��r
-Aȗ�k?��ϝ���%E7���D�$�MM��x{]���]��v,�"e�F��N�t��]�آ����\��N��[7�+�a��w�QN<,�}lh�i��R}A`;v�q�hr1N�Z	eKJ"&Y��lk�HS���zFk���zgG���'-Y�#�]�o�I8�]�|���}k�U�w,��u�|����|0I��c�Ï~�q��=�|y��Y���:��N��z��x�!,w��k�6_�n�}���]�k��i^��@�vv��ܰ�Cs[���n��5��jW�kz�mm'����?lJ��u�#�s���zD1G�Y�RG�DC��-�,�>�_�@�\���zm�0:op����c
����g�/!�8!�A��z��f;"���#%�q(2��Ah��|���SC���cgEH�B����ޣ��4.
n����_�%��v�pݯ?��0@���dH�E�/Z�hѢE�-Z�hѢE�-Z�灍������Z��ֺ�Y�_o���mw�|�__�~]֞�4:.���`�GП��>9��bK��އ_��}Sч�\0���<^�e����>���e���qUJ��G^nD�}A�fѻ�\x6Iǥ��Tԝj��]�Ѩ��^� ?��v/�!R����8y�����uE�<~R�=���1�y��"�j�hÜ��� �{,�>4�7�;��}Ó�FE�f���CQ�~��������������+rSo�g���o��$E3ᗤ�w�䒗/����cq��]��	+��72��m�iN�_���~�]�Jҗ|�i���ޑ���Z���k"b|~��x(��5�y5W��l7�:���-~y�3��~�^�_��̒��-A2>78Ϣ�yJ�B�����z~��5�>����'�������/P����׉�A���9p�c�X��[�"�s�9�{7|_����~0�=��܌��7��M�2wknv�w)5ru0��k�p����4X��03;h}�H`yԷ%b�4Y6���C��1y�[��;RÙ�����>I/I+v��͇�'��?�C�,I��nd͓O<�����������=I�{�����*�����e~�$:-R���?NR]Q��_hL����I�]���tIQ@����%�%��.*���<G\M#y��������y��o�k�}�Km�|u�R���#�^�f�wZ���v#��;Q��߷�oc���F$�*
���%����Mһt��o�z�S�|hn��ޒ��Ҿ��خ/��i�i+�1Eq_UTշ�OF�ݣu+�8y�{�?��&�K����yi֊�B3����wu����)����F|���������ζ�/�fڔsV���q�ߏ9-تw���ֿnW�JH����z��\��S��1!�ɉE2ϓ������y�����"ԏ����)
mC��&�n�n�Q��|lHK��1����w�p���xUd�HȞ���ʾ��v����S����j��آv
6t"�E��7Bb��'歾���q��垞�k�(���ʓ��hTm���T�-�7D	�D9��Bkp_Z�{Ҁ�Ւ�����wAdg[d��SF^��I���{�V�S���e�Ѭv L��~���7&b�)���Y����7�>���g7N��(�9��u����І��iU�t^�u^������n7�t�z�bT��HEx�ʹp+���o[���|�HU4,���x2�]���Q�"��� I��5�H�Ӌ��ÎƍG~$I�"m���+e������>�Ѣ�V��{��:w�9�S�C��ի6���VE�Vdf]ڙ�m�7�׎.o��iX�{��֯���~_���CF7Pp>?���m2�j�rQ����s�;dX��O�_ƴ�A"-}�d�׺ۭ?��OC��W�Q����ܞ���$h�Y��$_�w4����sd�u��vj�/�m[;� 	��9�y�zA���y�EaVF�aE=���	�-���x�}��Q���j#�qF_�"�-Z�hѢE�-Z�hѢE�-���J7�&O�uo�W�2y���%󴧈�����$o*s�(�x���(�0���3migw���������{���$�h�>9��"���G��!�^T4#ʃ(��#��ɤ��H�@�0�f��1�V�_IY׽�y@т@kk�c��G4"��(8��f��ԂDn|�yy�sq��}�f�>S�۬@�H��;���$����_'��Ư����]Iz�Yk�8� ����e��/Y�~�s�K�g/�GzW�S�4B���c"�E��X�j��?��"I�y4�t��B5D���h\W6_���0+�H�~�D���9b��Z�'.yr���B�_n^���7���Y5� n�G��d�H�@��=p�8��-8"4hO"�9_��]�?�2�x�1��A��"㟫�`-\�a��i����b�A�h��3>q�i'�3�/2�A����΁?|�iz�F|�={6I���W���i����zM�����������6�UE*�.�҇zQ��k�Jj^�f�P��2M���F��[�<���8�P��92�e�D�D��h�Z������ĉے�N��|ы�w~��?Kj��"��H�+�ͷ<&M�����K�yQ�~̢?��I�:i�����������oH�����Iz��Ԁh�T�����?��L�ǍT,����h���TY$��RyP~�o�R!C;�����Y�����j�绾ȯ9�o~��\A#$T*%�� �h7l�������sλ��N���7k>v�?l;"R������!yɎ�`&��Kzix&��7�3I�:����8_R�c�y���yi�;R�Ek����wD��!�:�8������]0���
�k_���w���a�/-kȚZ��A�_�� �0�:�t���5"θχ�~�_x�/����.����Yg��j#�%���!�o�Dh�6�ʆ�i����t��u��������?|·��A���_H�뗍���c6�K�~i�OI�ri���w��FL����$}J�l> �R�܏
�ַ�5I_���ݘ�ܖ���c��{L�g?kZ�/{�iG��4�Y���*rB���;~tn�.48��4�৿���,�r. �Ќ-խ���1ч���\�1�!�0�m7v$@�wEp2���MY������ﲎ̚|vF�~F{����`�}ȴ��y�६���g'��*]Q_��;� ;(ى�)2F�D�&�}�YW�x����w<�#�}�;Z}�tu;�����܎��	>������s$��E�-Z�hѢE�-Z�hѢE{Xi�;س�޼:ϓ}�כ�	yl󇼚��<A۬�7�Ў�\n|�'�&�h�A�����`bR->}1�HJ�8�5���h��:�%ˀ(M���#�{����8ώ�xW���r5ȟP�=E-&�!�Ct����y�O��<�=.<m>�
N�~t�:nI����(�?�Ӗ���0I_/�4_��L���5#���y�+L��@�'J��i*4�*lo��V͓@{��_��$���1;�@��a�mg�{�1��a���\	�ê�iP�|Oq
��|���j#�>��(���?n�V�-�Α��yx��Z,��C����xȸ�$�����?�'=�r(���ȓ@ï�w�Q�g�m��c�|�!Q5)'�C�^��tf��P�yygU���#4�^v��	���Ûw�׿��I:�h�?'lz�<�=d�]w���'��k(z����7��ܧ�g�p��DQ������?I��W�*I����#� ZW.��$�����~?�??������}�p]�u�ߡ���ݖ����7}˷$������[��>?�9#H����o|�d'N��t��o��?I�4`�9�$�(��_��EI�������'IZbƈ��*a���×�G?���X�E��v���^[Ѻ��1dMA堜��y���J؇[����0���ŵ��d5^9[!h�e5��]���j��ܼ��#�HMT������p�z�߃!S��M�/4 �<�3�>>�v�qE�|D�&j�;N?�**/ϯ���}�2'$p25���̵ �7$9.gnc�HU�~\�['�8�X���WLo�mzGxgNݞ�m���ߑ�_iQ;�*z~lԩEK�w�ەO�V"��KI�䖢����=Ҏ-�y�i���~k�1E��6&�o���>�_���}��j�0!-~v@�5�t^�d�ȸh�B���& ֔`Y�m鹶�q�� ��C�}��1�̧�ݹZ�e�z9����E�����#s�w�?��Ra�}���J��q�S^K�@�M�j�$�Y�|-�d����1�i�ǅ�v>���\H=����큖!�������hѢE�-Z�hѢE�-Z�hўV��(&��sgM��ҚE�1O��Z�#W�=#�,O+�;��W���&:؞���rB{�y3��u� ���ΓmY#�h�K���u�s���u��,g^w�0:�:Gdj��#����y�{�爻�_����V���#6u\u����Eg��S�9��<y�2�Hv?�~�#:�xs����;�����**ߋ0b�S��d��Q����T��N�q@���0/�y`�|�4$���,�aE�����$E����e���g�{#ړYh������,���߄����㞳3>��)<���!K���-Ϳ��QvR�a���ӍH�1?Gժ	��
��C-&׾�Z�pA��P�0S
��;�w���DG�e�'�ϊN��7<� �N{���8�k���3���`��@u��69s��$}�k_�����'I��H��cFzA��\7m��O?���M{�4��pk�,��~�&��~0I/^0M���JR4v*U���0J]Hv�]q�:�0����/sw��"Z��]�-���/7M��/����2m�7�id}�Qӊz�!��6�5o���!�Hs"����_W��|�ֵ������[I�C?��'i����E�|�FW���q@T��y�wG�\(I��6� �NS���2R-3^qZ4&A��95���� �u)�
��!���߉
����o��(�z��W����v=Ȏ��}�U{�hO��轝ލ�5Bhg��H�E�}�kM����u�s�!�Q�����P�}��<'�A�.,�~�;��n�2����0����#;���a>����m.����[^�|ꓓ�χ~9�<��sɞ��g�&)��/+�m^��~��CCQ�W�=�ƙ���w߭�N]^� �G�%c}��c_����3�m�i���I�~�w~W�V 3{�'h��i��n<@߻��wR��|�ps�kjw:nl�H�ͭ}�q��WlZ<i�vN��FJ���Y.�H��.;�j�J��0����<�sqHB:�ύ'�xDq������9��vqZ�~Լ������e�[O��	E����e/_�z����P��y�$M~�n�_�9��T��=
��)?��N�V렾?�P���y��?���z>�9��j�D_�hѢE�-Z�hѢE�-Z�h�+���H*���_Ko.�9{cj�ތ��ۛ�~����Z>����(Dm��8��S�F�7�k}d�KJ2�L� ?��0r�H>�F��h��[����r�nH�`SdZSQ늁KOM�Io�!K��6I�F >�%����W^L�DLF���#������iɍZ�����`���]�J��*�W�ʴ��7��v��MN�rz������LT�� ��궴j��g~������5IO�v&I��-I�v��Ҿ��yv"sQ��4ؠ�#���Ѭ�N���<VD;�E�o
�e�䮟���v���>��#d�>��4�2<݅B&��Fk�����?_)8���/Վ3+J������s�v\օ ��,O�p(��� p����y�@��W�G�}��0*���oƴ#�԰��oxm���g~��'�w|۷'鹳g��T�t��O��Iړ�tjʈi�R�ע;�G?��$���g����$���?�g<��,��l�V2	���^�`����a��������EH�r@TQ��u_�uI�����$���{w�����ɋFf��>���4YT4ޑ����&��5E�[�Fѕ�����4��{�����$m6����8�E/��^Y��M�ӿ=����٩#��������'�RMI��-_�F�r��:R�mi��c�i�gH*��o�l����:��NKQf�}���0_|����y��E�9D�a�F_.�}a���s6<��I��χ,���9���p|������;J���Ӱ�\��'�a=U��ў��4m�?k��e#���q�8k���hZ|����{N/I�R��z�Fe�����&�ʊ�3�B����/I���7$�;�F4�}s$����,����0 �CR��}C=mZ%s�Z�|v|�H��-�|S>�Ǹ�F�ւ4��clYZ�!�G��Q@sY~q�u�ΏpG�Qǅ�v|(Y�S���n��s��݆�g4ƍ�����y�x>�A������ǌ���P�Ǹ�$��; �B0кU.�Ҥ����<�f�|e_�/+Jw͛�����#�-Z�hѢE�-Z�hѢE�-���Jm}������d���*p�Fi�U�$�|��ѿU�w����_|����ҨY���Q=kx��e���9*�Jo����|i�<m�!��Tn�Ga}�<({M�����[D3�B^��	����m�/��7f'%�xC^�!OvI��~�/H���W�(F�h��҅Y�<��'��,��w������?iD�˾�eIz���WVA@����)����T=+M���ȇ����y~�?�j�N�	�'�y�(w��}[��i��5Z��,e}�#RQ�2>�Q����YZI%y�:�l�KS�-4���G�s�}�c�u�(G�!𜦞g����n�!�/<M���@�fg-j趈κ<��]E�R~�-͡ɉ	�����I�'.K+�M=fx,u�.7<�Y�W> (�,b`$GN+$��O��k?UNU��A�n�F��A�B<{�H�gy�sW&O��'��~�����? %�C�dx|������0 �B�/%q�<�i�.��nS���I��G����_��EI��_��$}�^#��G���~w罦���(j�V�s[S:�rG���>��$��5���W?���>k�y�c���-�ۘ���n2m��2�?��S�Gx���&��z���Ҥ�lIÔ�Q�4T��8m�K�'~�{�q��r��{�l�\�d�TT�����N�w��?'�'�l�.�Ɣ/Ecܵr.?i��}i�1~��m�a�j�|����|>'���N#��v^޴��6n�A���;8Y��GD.���˝�͛|>�H�۲0�g��<B�4�2�� ��;gc���n�	H��/��I��e�w�FM;,�NX���5�8��x�vDh��t4�e�[����y!�׎D�sG�)�����B;?����g�?�7=l�?F�f�F�F���\8��;ڎ�#�|�|���Dmp��7�P��>��j��v��=��~���}#��/+�|��H�4[~}�ί+�=Qx?��O'鎈����0I�kz����"(�#>�9l/��u����D�zD�������l�����^��w��N�NH>l��-��5{�FӯR��Y��x�\�q!��|!��C�:��΀�M�o�?���9����j�yC��t�x��ʶ�onǏ�!`�v(��IY�q���汎v���� �xn��oX7��1�:��%�0�-����^@.:�����D_�hѢE�-Z�hѢE�-Z�h�+��"~�ܻ7����B�z��7���E�|��Q�[%��~�iR�&� V4�8GWJȄ����Nώ���������h����D�䍰#�<j�؊�V�7�3��a����o�)Y�6݊<��yOd׺4p^,����yx���f{�*Lo�!�и+JbWd�EE��hO8 C"'-`�<\{֫l��A��)O���4��z���k��u�҈h[�~��ߛ�oӓF�z���A���&��A�1��C������M��U��v�鳦55�����9�l[Z��n�((�D���=�����6�hV�JKdĄ���̜/�`c�<j�[vݢ4+c��yVZs�~��i����WW$@O��
C�S�4A�K�%�WH�"�F���ew{�+�p��3�
�jծ��M/ȏIy�:�֞&fEʊ�I�=�ǫ,`��1�~�k�nD̚�ic׈��	��"� &՞�hIU�ʡq���XP��k�i��6�iYṤ��QD��y"U/x!R�kx��9�	�P3�z)��Y�6(�[iT͜�}����x�T�U�Q�F�aK!�A{sJ�7�)ζ�.�����y6ԈM=���F>ZBiT4�0a�F��ɱ�(l~Z�D ò4���-_������k^Z4E���g���~�ǒ���iD�����D��vI����x�sZ:�ϞJ�j�����ͿJ���2��&����^@��~#�����{%u��W�s�.�<ϩ���D���{�lbn=�Ā,-uU��������o�)K�}����x��Wt>K�E<���[�qr����IJp��4�js����������!���yyƩ��:��;v<�TM��46)ҝ�0/����[{<)"u{"��~�eY��ظ�cO����u��O��!�紫 ��,f5 ���[:L0�������W��^�uĈ�h���I��CH��Rn]��~K�i��fD���D���AX�NJ������x�I��r%�s�����	H�0?� ?YF�5�Ӂh��.��v�����:����+-r�KG��ܼ!��A��nw�ޞ���U�m;��.z�����\J��so��>�Oq���RE���κ������]���I���F��s�]Iz��I��+��t]�pw�士��{���c6?��i���,
���7���F��v6�hV�k�`���|-L��X箮�|?��q�kg.���H��
����Jsxjڞww�u~�����7 *{E�e'���5ƬGˊ��A��y������EaV��z�uS���V��N;N���0c�����/���u����wO����.d_M�WK念e�S�$�ϵ	g�U/����5��y��}O��������'z/�TO�M�!�;j�+�$�{�`G�{n9D��D_�hѢE�-Z�hѢE�-Z�h�+��;]�����P�)��=u-�����������C�gf���l�F��?f�}���Ͼ�!��.�oR�����*M����I�F7C��]�?��{ܕ�~��*���Q=�k\7Rox�<�h;ml������p��/�=��=U��-��3���-}�������|R�,��v���ڻ�q>}��$��sx��{���e��s�I���yyho�w�,�x���˛��',��+^�p�nK#��5#U>�E� :q��I
I5=md]�IQ��}�<���~���r���Ė��7-[��Z�<�N������4�	�}���ɇ�z^��bE�[�go��o�%�;�þ�oK�<�]�9(Ox	H%��V�<�3�U�������?��@��<�y���8Ry��X��H��R3O͞ʿ�h�S��/._��Z�v�����&R�!T�b���[9��zWZ(��S��jD���<lx��h9�-(y�  k"Ww��[y�GM�Ȟ��mm+j��G5'��SȄ1yĖWM�����v�vG��h`�lSŠ~Br����b�w4�9��5h���\i�ơ�<�h�AxM��<n��7�Id��ȳY8��X_]��}�b�t6�r�u}�1Hl�!<�x2�]���h����`}O�(D�㯡�%�g��w����y,�}C�ݞ���42���u�%"vF�㛿�[���H�+�6��w��%�o��H�����`��KY�BM��^kQ����v����IJ����_���M������}ߟ�8t���O�wр�~�"�I�b��X��=�ۚ<�i��"�i)��9R��^:ھ��~VZ���4g�ڭI���qO�eR�ә��!zZ�ۺ����a�S;�yM��E��Z������W	bݘ���e+GW�?b[�._���ٸ}���0U�)�G��Zi��}��E6���h����e|�S�45��(��ƭ�������ag<�n�<��#���+�/�b?%�-������Q��5�����ma}=��͚濥%[glhG	=Z�R��eE�BRA�/�������ܹ3I���O&);:Zj�E=0�NLZ���|B�\��zW�@毴�]�j���<��Dָvz�\[���!��j��o��%�~BB��R�uh?|��zS�ACzQ�c�s��i���[�S?�s��������Ӷ�e�ڪwn޴�!�77��H�1~���+�.lgחsG��������/;���t�9�QS�T&:(�%�:KI�െ]fʞ��E�}�S�I�/^0��̑[Z/A
�0?i=Z[�u��]��O��{���"J���?O��?����{>e�u�ʑ)h������N;N���u�,2Z;�Xf1��I��Φ��n�'lg�Fv�0�r+��r��a<���|/��q*����Ar��7�����]���PGD>Ĝ{.`}��>���N��Nmw����Eܑ����L�v:�y����ow�`�y�����g�m��'܉�������hѢE�-Z�hѢE�-Z�hўVjuy�xfe.�a��}��
�7G ��/�3C��0Q����{S�A��;{3o�G\��o���O7�/zb"���.���\�ɐ��D�K��sxf�M7$__�h�@ïi�F�.�����<ЅΎ����;�M�y�+"k�94�DfIà�7���%�
�-_�}�Q]W�wѿ2�5�'�vħ�<U]yf����|����g;���on9��-1���=�Ϧ4�N�m���{��,��V�.�sӔv �ڐ���Ȳ���"�*�DU�mɣL�W<�.�/Q���Ӵ۴z�Z�f �-k�=<�D�T;pڑ" 4N�u�bUdZ@�����=�>M9yf&���h�Ṭ)z�����n�g�6ET�/<�uiw�9��hZ�s'O������)ݗ�7>m�Q����4��V7Vtb����}�b���'�.���(�r�my(��w���V�[M��@�k}j\��z@���cCc"ȧӪP�:�;�=����h�@b�՟*���Q���LY)�GY�c_��W�H2��y��b�c'͓��lܘ�3"aK�@�����l���W��rQ��|4�4����H3����ۃ�/�C����R��U��p$Z-���cҸ��vm��2�"z����r�ָ�}�ʕ���W}M�޿��$��y���pƈ��#=�D�\��vݿ��G��ů~E��݈�=k�ݒ���+F*��[> �]T�P�O6;=����Es'#�p`��X7�!��G4��@�9�D������iO����Ĕ��"�t�=���c��4�m������+OIi�S��u@�n�Fl���Ꮗ�2ī�m�@�G`�M>���X����|���f�S�];Ȉ�HGR�ƹ�Y;sϮ�ݲr\�<_7�.�C�����V9�]�xi�^�H���8�~,r�;�lQ�ȣ�d燴��tǈ�1��|�굥u �Tɷ�r�^42��1�g�Z�D^i! ��\O���i#��	16�֛���n�Eۍ�����k~A{rQ�QEDjS�՞t�;yi�M�[>:.jo`���yN��e��#ڲ�B̻h�2o��E���0�C����Ԃ�?��o��-]�nP�&�@��P߅TT{�׎�MP�M퐨�!ר_l�whfj>�XOX�f&��1nH���4�����[FTLl2 7��� Z��[E;}�0����=���E��ݎM��(�}�Á깭	���]�Q{��z��w&)ִ��<b��3S֮jm��Iv��������@�EGh���;*��+6�絎�,/MH���(�4���A��Sϧ*ֲ��Y7�*v<�t4�w["R5_0��N�3��~播3��6��e����D���c��G~�Ɲ��� ���|���7��L#?�3��G������;�'�-v��x�O�>G;F25B�� %Y�;,�v-녀����ב�|�������p���1+�D_�hѢE�-Z�hѢE�-Z�h�+�F���ǎF�|�����*��+lo^v�fy�C7G��$_�����F�v�a���0Ъ�SzT�|�u�/������^t� v�z#�H�4�Tp=���}r�|���niy��hB�L�\O���y* ����fO��s�Zx���3�7����\W��*��pHT��w_�P�J)ȕ�T�=OׯK���kM�'�+[9V��zx"���|ٴ�Ф@c��<*xܥe��Ҕ�g�*�eQ��r�����h �䱧ݸv7b"B��Gv���˳� AP���Oc�O��%�A���jWD�͑|A7�����Pu��4���[Y�����h��s{���<��Ǭ��<�x���Y[3�ozFږexEѥ0<Ɍ����<�.z����uv޴� ׷֕/��1����>����> �(��Y�Ͼӌ�#�j�8���m_S�d_�JQd�ˈ����Bָ��h^x�'����e����J��㴨T�5y�9>4<�U]_��>�Pc���#�<��oSd%Q�U���TK��,w�<qО��c|���y��Yã����86%M1�������㝟���g�����Izj�$�tF#m��_uO���hl"4���}I��Ϙ�Q�J�_�6)ѵ����c|��;"��jG��S4���
ڹ��
tĽs �s���BbRQ��M������� R
E�}3�tE���"Q�e�Չ�Q�_�V,Z{��Ę���}�4��M�W�R�5`j��Td>��BC�Ku�%� �!� � ���鹽g�ȸ�u��)#��<k �}K�iO뵂�ϲ{\��斕Kc-4���$��6rčo"ӯ]5"�z�:̇������K�P��T�b��"?�W�#�#���AO0_*?D1�&��R��u�"��G����ה=�ћ��U�-�2�oYZ{�����WyT?MEud�����j[�褈�~�dH�\`>IrY�����kZ��V^�h���Eױu]�{�y�c��<o��z��Y� љwK" /\�$R�vʺeU��⒕wm�ʉv��$RUG<iP�|A:�g�)�|eٴ4��E����mE��?���5?i����M��<��<�f���%hmBxӾ�ڊ�F�[oh\�S����6_�����|ᴂ����:L��=4��-��pAv<���h�":��Cλ����&���$���Nd0�$��]����wx�);�d��y��W��K�8�S�����Iw_�����7�9��b�:x[�܍Aj�1�T��V����GF6�	2��:����C_�RO������~�R?
˃uMC!͆����V�C��;-��0��r"�-Z�hѢE�-Z�hѢE�-���JD%b�o���J�ey�����7���K��o�..j� �%����G<������g����˝u���_�$��f���z����d��;Z�SH΅�*y�����7 �-�O�A�8-}���4��ǔ����;$��Q�,l�|B���35E�U�j�c�ȃ$i�`ZL�W��\N"1�d���pڍ�[t7lI�o�5(mHt ih��G�(JhsM�ṗ���;nQ���a�4AT�7���FT�1y��-yU��䯯�gpl�<�����_<a�ҕ�����F�3OR�i�X�O�4� �mg�$�{L��!O����q'�^�G�y�T�x�&���
�=U�tN3'��� ��*D}uڒ��iY�4P���+���J3�^�A4ki�H#�EU�p<q��_�d�`A#���J+2%��Q�a��z���0��*�ª��t���A�ST<�ѕK"P��!��C�|Ҩ������B������E���-�V������u�|���T��O��8K{d�{���G_���d��	�M}_-���iG=�[. �3z4sڇ��� �1�N~����qJ�Q� ,�|�$�D� g�?�d�z{�6�v���>��z�?`�t�Q�O����"r�E�Q�4FՐ�EECUF (f�WBQ?u��j{j����u;���(�y���c�.`ti��.g]E�d��A�'�`���V�6׷�7w��"�+%�i�D��:e$&�/z�)��]kGx��ݺ��m��������\��7�C�rs@�?�[D
�O壮vyB�W�FdFUт����vѸ���R�!C�Bx���x��F�.��;�%��_x<Ig�n�~c>&��K�$�Bma�4�!���
ͺ�H�t�c�HN��;Kh�M)ʧ�G�h��{�������:q���-����t��31�zD���w�3�ݢ�;k6�/�n峫���b|w�iu��"�Q�}��~4)���b}
��H�!;f��鹚�w�R+O����~ʸ�r��E{�V�wÒ�[��~ǏB����4���u�_���j���Ɏz��h�쨠=Ҿ!d׵^v��N�+&�~w�v�;�䚈OG�@v�h���Xυ�{�V|� ��0�Cf�E�A�B�E�U�\ �<��U4����j:�܎��,�v���\_���ʣ_΋��q��p���eE��a^td�Hq��) ,b�W)��Q\�0�!����7���ʺy8D[�1mګ�ê�"����s\�Ǹ�&��<=W�h~,Kk}R��c<(z}����(tчej���t|��ߌ�ཀ�6Ѷ�!#9/#�}&�����X��3c5zB/H�6�5��#E��4J���R�>��'�$}ѢE�-Z�hѢE�-Z�hѢ=�ԃ
����<D#��9��{�ƽ����\��X$�@����t�ݵ�QE���ycD�K��(ψ�N�"u��\��4iBbNW��P��j��o�۫N��w��7-�������Oή��S괮��4z/�՜��bv �{��>�S��m�~���wC�MD�Tu\U����_���G�s�P��f��yfz�z��=5g��|�Lҫk�9�L�#F/
��,����C�ȑ�Ei��8t��v7�u�v�֚<x��@�*�
��ӳ�Ds��I����LX_���ꊾ�����z��MÂ(�h_A�]ij���B}�h�xb�8ɹ�oh;IsLw$_h��gk�����L@��h'�9	�k�όg�=i/����+"� 3VW�(ĐL�֙�[�FȓYEk��x.��5��±/x����K����� !�x
� >�nf=��i��no(���G� $�Sr�}����g�1���� :-�ݬ}BjAJ��*�-�@)�B�d�������pwZ�A{sY�<%�䁇T��?ў�v� Q�x�Xt��-�Pm���O�	_HG��9,�D�۬��>d���iM� �r^�!5&5z�Y��O�:�K�왳I��&����z�����߬�%��y��r�nY?��7�hw�Z, ��1�hz�j�D������߱ra�D�v��Z.4'� 1�/��������q�&��e�'$����ꞍGhv�5��KKv��u���H�V�Ҏ�u�khU���uI���ɓ�� m����/K��O?���aM����HJڡk�DU���"�y����~S�Ͷ���|��eU�*k��g��Ҹ�xԢ}���N�p���ڰv<.ҧ�f��kW�a�%z���S�Bחm=�xbɻ��˗�?��Q U�kv������Y����݂�'�d˾4��t�GHힿn �kN�w]��_	�q�ui�2�ML��e�ݓ�������k����%�n��agD$�KӰ�G�Za�)�T3�'}w5^��>v�-_K"�]�� ��l#?<���ʼ?�[9�׸@��i�����)ճ����n�����es��l��·����%�ߺ����|����}�����|��Zi'F��k���B�R��F�e��>�~W�m%C0ո��O����+��3N��l��Ӭ�XWҞ�&�Ɖ�H��+G�ϲ>�0�[�󅋶��h]>�uk>�gg;|hϬoWE���q��EW���GƤɺ�)⻭uF^�aa'��%E��y�v��Lh��Ze|��Gi��X��A����Zۻ�o�^2U	��<�vi�2﫿�������<��[{���<�v��^%x_����5�v��=����
˛%x��h#17����D�!�hןݎ�et/���CT/�s����D_�hѢE�-Z�hѢE�-Z�h�+��MpH��$�#�ܛH�x��8	�cR�Ao�{C�sjD2�֖y��7��n��I;��19_��i	� l�y�fo�ui�T���ey�+ei�T �|OL�Vo�y�=�ͷ��3�����GX=�	�FR��d_���~�&\uW����|���l.`@B��и#��]O(d_A{�y4�DR�]��e�my�%�WAQ^����7�6I�ݿ��C��eH��T�v�˷~��)�o=�syi!����/�i�%Iv�w��[���wuUO�3�Y��"� �C"�&QɠA3�}�If4���� A3 	q������Z���3�Eh�}O����qofVuw�χ򺑱xx�{x�y�=A���Y-z�JJ<���H����?�=�2x�:D�qԾc�A���O�z
o߹��x#q������7eh�b��Z�k������������OE��Q+���F-;�j���e�������T�~S<��0��V܊�ܰ$=�$���<���ϵ��O���W�Ԥ6�1�z1J�j )IO�C����ISMM��(�$��4*��N�ƨ�h�z?���	�DI���7=�5F���<�$3y��U[��D��PSʴ[�FAT���Q�U3��*۱ԧ*�+��H(�������r�ڌq �M{ߪ��������5=�3$�����]�z@>�^�"�G U�@{�Z}?���?���8e�hTHh�u�)�dT����5��Դ�{��hK�@#3��p� ��}پ�!���t�j��<�6ڮ�z?����E��h����4��T�$�	�k�X�I�s��w�$����K;#��~�����Hd^�"d	qj�u�p�;��z�P:�W�2a��*h���gN9���{�ۃ��ų
���Cy���l���}��1,-QNӁ�S]�W�ANRs��eM5��zON��2އ��7�BF�a��|l�J�:xBR�R$�v�
�[��B>�Ϡ�!�=-���Z­����X�X}�Eh~�\-1�`��p�ə�_Cԫ5��i���x�ϯ b�h�����7$���ҭ�?#�I�Z�hc�L֧)��А�}<?j��+ե�{�P��F��:W�`{U�{�#�g��~\9��]��L2��qr��0	B<�q��?��)�˃��s\�&����ǉ&����8�ڔM_�������H�&Vd56������T��ݎ�_٨����JSk�`,��ޖ�IE�5�#���$���������+���y9n�xZI0��[5��~:��U�ö@�S�ߑ-�;I�s�tY?���u��p�O��=1��`���r<Ir�$�% ���iJmt�W�p���;����^���$��޻]j����c9�<+-w���0ڭ�?�|y�~�1�b���=9��PU�|���?ݕ�W�-?W�J���J6;�wT�ھ��(�̮DȚ��X�hcG��)��u�a]I������7b��d����E��,��J!�ԞA�D�7o޼y��͛7o޼y��͛7o���S	�MT�Ό�33���gf�2�c4S�W���c;�(���d�cY����z��h��'e��r�$.��сx*v��d\�.��V[<��6ECbeE<�p��vCh�H��弰��'�=n�F��SSH���r�?� Mu�=�C� Q��Jʗf��0����W�H��hC%ծ�2s=hEF��i@B��u�S�G8Ţ�<�Ӳxh~����8��X������9F4&��;z�H����3�&�3�ѧ)Ғh�a7�_D�Y���<�����])z��LA�⸂s��C��Sc��^M�A��8R����.IZ�Qw��`4�=i�x�E�Z$�x��4ѨlF��ZiԬ���j��|1���l��/$I�hi�O��Gz�x��}�2Z��?����@�G��Y�!�GR�!��&D�h�n�/F�܂Gs��h+��;A9�4���{�b��e�7�ȑ�a��Z+$"5��d����d	���Q���Z0�j��Z�IԮ�?ZU���9n8BtV�Q�5����������^���'J-�F{d�P�x�N@��P�v������D�|R��-G���5��J���F1��x�'[�-�J��ԑ󐰣�əR��2���A��`8�ј������X	U�D��M+�Qo�}{�w��o<^j�"�W6e��Z��q4`TR4�|��"�rj��/���%��&I�=��{�*�� ���h��H�oD����9t���B:\�\w �B2�
�����kEY����{�+ם�d�FF= ��lK>�� ��U��U�h���s��\��~t"υ�{�H?�q�
j�U�qv�Qӕ��~���ҨȒ����NIw"�58a���α�W����������Ԁ��+]�*'�=���ن���):�ݕ�9I�v�}���Ղ���=����P[d�'�w����}R��(��Sb����ԯ��i�h·7U0��H�<��-)�c�ʓ	W*���ۛ=�v�?ܷ��Z\��"d�/����� ����:4|�dU����]��(t�+a���D"R�O$�H,s���������gc�����p%�����q�)/�=[B�24�,yr��*�������X�.�� �GmĪanys��ͮl�}��'7쓸��.F�Ǌ��j�x��=˟���#	�*�G�2����T�~B��L�=����8W��@�Qs���h��s��oBss籐�W�?B?�9ݛH�@���#hL�;^�3_�M�x����Z�x��%7I�?�x8	�.��t1N@>�ղ�����c��w5Z#��x?�+�b���e��dܐ������Cv���R۳5;lOi �����<�"��zݜKp��h��hV�Ӟ(�����|���۽<��͛7o޼y��͛7o޼y����+`e�p3�-E(Xm"��WHj��:��8=;r�+�h99�wF�y��?��7�|3N�]h�l�������o ��i8I��p23O�\�hF3;|"�KW@����U��>	��s�xJ�)�A�A2LA=�%�f�a��'�}#�<�:	������/J��/�F\�O�	=�	�|���U2��Y��}.Y7��]���f�k�@�޺s=N�y�v�Np�!<!����hCI&�#WpɊB�%]�eFSO�*�@˥�DF �0:�>o�"�����X^��^�3�~�P7�j�x�<��P�
j��HZ�'�ѨH�G�D��MԐ )�!�-ʍd���c9��l;��u�9c���nP���5訕Gfm�ո��]-�CQ��)d��<�c�m eg(�&��Nݡ�o�y�G�5j�� SO4?���Z>x\Yvx�S�u�2���F#��c�{$��I�QՍT�
' �JFˏ�COr`�q1�z��E�Se�}��>��V4Z%���_�h�n�EJZ�R��|>$�J�Zd�4j�����@-�F$�H~P�h�ǒ��e�d���X`�btc�E�gE'_,��y��{��Fo���$�[h���)ن~����l���!=�5��̾Iq�T5��H�V#I�V{���[���#z��t*8�����	�|*��/��'2"17&a���Ѭ��*9��E�tw�#������ǌ�-��c������%�pԿ��Y5Q�W�d���h�����uG 6V��֧�$�#���Ix��^�i�	LTj����q)�O:$���)�Q���b��c��(��4�oޟ�e�{�`,c��s��Y^-�o��9>ܹ'D[!\�?���$��9f��N��Dg���T��ǽ�{?���F3���9� ���6y��j�f������l�D���%'$h�q��9v5�����@9�LZA������E{������ [_��ɍr<��u�i��M��&V>�l������ZG4�1�W$q�P���b|3��u�_)Ɋ�:4���!�3�n���E�H�r;�����P�㜏��)����Aǳ?��^�v@22	H����zL"���ɧ����֕���5G��9�V�ύ���ԧ���M��=|o$+��~}���|�>ۑ�4>������éU��{w��iI<��w�oe��VL�d���� �XE��uT��\�Rs�=��qɝ;�]���q�kפ���X����5h�1_e�V{R����u5��a���̼����ُۗ���$�rl��xvB^c�n���%�f&z0�" M�BCB��3�AAF�軶R��y<��͛7o޼y��͛7o޼y����+`�0cF5=c8q2��zZU�̐mthu����\��?��8=�B�"��C7�y���׿��8m��_��c�	��Df��5�mb�~�hkex�۲�&�9�c9Ϗ~�8�L�F<'7^�����	g������8ӝ;A8ǩg�h��3��E���D=��,�HV ��a��?�H2�na�>%�B��H������(� d�^Ex"�6F8����mh@�'�,��	q��?2�s-2D���CY�æM#��<;uW�c�b��ܺ�;D)K�.���ݿ�#�.f9/4��W��R���z ����sQ���\w�|�� ��� �g�}���X��~�!�Vc�!�xl�1�f �c+���SL��l�?�zʎ���~��s���HX"�(<u$����MM'F���y�����}�/�F�;�g�!��v��F��'p2�Ѻ6@$�Fʅ�#����D���8D=N�4j5��j��Q���E�����h���v������$�����P��j�Г��*!���A4�WMDs�g�d�Kj/��Q�T��a[E;e�BK�~�S!TXf�K�ծ������2*��O�)��X�s�'������F;�ɣ8�"*�U�Ӊ�&oH.%�r�7���x�#�BV�v��
�1�w(ǣ#7j�����T�Ԓ����h���s̸��RLE��d#�_;^H{F�u��d��x�m�������(\�`��c�5���أ�Q׹N�����U����0'��S����%,�v3>Q�HX�1:2��)F}�@�bē���H`Z$YQ�+Aٹ���3�y������ETv��7#@��M�z��s�E�dW�Lq�	�����H�}��ݻ �h�|��6�Z�chH�#�Bw<?�	H�]�۽�ch'��}/gf���l�Ew�Ͽ�<�q~���ߣ���O���
2�pc��q��ڊs?+3J|cZ�x���KR�-5�$�uܠ��Ԡ�;��MHx�렡��=�sHl��#9H�k�+3-�%9�X	���:V�p<���$ʍ� ��e��V
���e����m�D���f\I��A����UhR��Z�$4{#�gQ�����"A���㑐�15�|��^��$�������d��3�k�ߵ�ys�Q�1��r�
���8�k@S����h���d���;�����p�e�ı㦬�T*j1L��l'�Ê�]�h;��s|�G���M��1a�g^げ~$4y������1��Le�eQ��{y�ϛ7o޼y��͛7o޼y��͛�W�.p��k��!� �2�ə�)�� �����8�\��H���_����'���~r/N/����@���]�\���u�;����e&�R Q�DO"��N9����Li�,�_��w���{��'B6��q�M!����rz��GR!ã�b6�i	˔V^�of[IA����Խ�nK�C2��g�E�7�A��E0j+��0��C�x����h�� ԉqW�d��>���AP��w~��8��y;N�%wGR�>���8}�#��Z <xmhv�Vb!��BO(4'����������T��Y�2�pp	j	V�Q��	j1��èNS��\���o95Ȩ�Qbt����8z�jh�$Ҏ���F��O�F�����Ƃ�ɴ����xZ�k�3K�!j�)IǨQ!��1x��$�eh��Ө�8n�0R�?���_��i���q�DL�9z�
�y���Q�����"�И�Q�"�ρ�$]��ǩ�m>I�x�9��!2����ymt�ѐڇ ��7#��H���2��_C��^G��p@/�fj�:�l|>�>��kׅ�+��(��B+����=R���F9��j�U[�Q�(n�Km�H��u)�������6���h �P�\˲�R4��F7\4ʙ�0˳4Y���"��G�ﷄ��wK�����:c�H�=�}l,r�In.�罏�ˬ�l�qBV��4��k�qAV4�I�%��K��}_����1�Y���;��W'���o��wQ
n���Z	�ML.y�~j��+|f�S��>��Ө����b�ƛ�
H:�w�)�q��U�^��sK&��~��~߲<u���@ml��
��|������s��K2��6�pWƍ$�=�x���ie��)ߓ��'ۇ CI�3�-�A�0���+C��(��-72����p�R��s�����X���j�E�)'_�GgD���o~ԡ�����B��7_��l�Τ\X���'���zY��!�h�n.���R+	�^�yD_j	��e�����j��gn#vA���F$�;A��]�f�����>�ϤVD�ۓ��>�|_�<��͛7o޼y��͛7o޼y����+`�e=���QJ@�`-�ѕ�vDmQ�v����ZK4�~�ۿ�?���}[�������D������;�g��!9�"��0Ŋ��!y�5���.c��^��J]��Νo�i�.�ދ�����L�~���O�Z��1��(��]8��ǟZF$�2<�SC0�(1��.!�<�G;�3n=,�t;$�f�P���$��{�xxR�C����haժԫ�1�@��U!L�!�ӽO%
��:�x!�+�%�h�J:��$�9�B�E�Q%K����?��8}��O�������}��qڼ,��ăU5Q Á��F������	<W�ci����#Dy[���O�S��G?�߈����|-N7Ut�F9�A��?D?�U�'jv�'w�<Ӑڞ�,�_��/j�X���D#�=و���*廷/�"�D�D3B�+�_�7�����։�̖�餖�	<���y1jn�N-S9�w��:������[�a=���ڤ��گ�����ΛBt��_��k�kJ@.�a�Ll��x�u�j]��JU���O�=�}�^��!�ݻ_�v�Җ�����Ԁa;Pr�����g��Y�mB\�ha�2I�餦	����ۮ��4B�M���g'�}���)	2���nF=X�l�X���Z�/���\M�e��-k��?�H�}:�u��jU~^��8=��J�q�5_T�̋
����hp�O���[͍Vg��\8��I�fY�˟�D_�e�W��s<[>�+xBh�C�O�xt(ߕ���G|��
ϟ�!WL0�:�q˓+��[5Q��~��R{lf�W�Q� �����0W��~l(�-{��$h�1x�|Ws%�ѓ*�{��C��d<�����~�]1J5�gu��8_�I�V���]CB�����1�ߍ����%�8H4[�ȷ���Vs?���@%wEL�eZ��Y���9� �ګ�W�J��CY�X�Wp?��
D)�]뎛~: ����&	C��3���~1��[콝�{��ǋ���~h���/�����>��e�<����L�4�!�3��̊ˬ�5}<|���a��2O�y��͛7o޼y��͛7o޼y��
ع'��L$=ֽ�x��i��v��E���!�n^�-'�!j'4w�6����.Q"�ί��O?��K � Pn\��� e*��Z73�SD�%�85��Fs�F }�]9~�)���ߐ��?�/Qy~*���?[W%�A9��4/�mZ�ȵP�d�ZY�K�=���R��.ȡ�Pv�;CY�0A��� ��>�zئ3��x`�³G�ɭ�R��1�L�� �㡫�քg��^�Ԁ:U���mE�W�Q�$�w۟!�h
���H��֯��8eT���ܵ���jۂ��QgU�Q�ww�#E�=��qҕ~��(`���џ�U��UF��>4���F��꒟qW<���?�ӵKB���$�Tp�	5GX.{;BS[�э�$����H�&�V�v�o������9���>�r)�96�-x4����T.������������c�ք���.�A��}�T4�6A���H�6��<G�r]���&*��d�hRZH&
�B����*1Gm����,K�O[h���g�/+��%+"�a&�,Iq>�V�%e����WM�!4�v�{����i��y-N�����^���ܸzɹ���������(��-��_w=�hO�#iG��KG+<�$�53���������2:�řK���I!K�[B�DU�{0+���vkY��h�i}6D���D��E(-i��s��I��b�3ky�i*�.WZh?�E���r�׹��p�al�yD̗���&h��eͯ7�ZfŒ~p�5�1[��[4D�	��+�1���Ͳɳ,����ݏ�]�W�A�<j(�p_6_lO$��z��]D�-�~I�3\	F�D_�U*\I'�
����F3Ǘ�G@��>W��m�;���25�48�Z�r� �k�[2���Aَk8 �2~����#˅��A6�Y�z��k��؃h�d���c�ԯ�\�Z� R�\��a��Ϧ���Tk��sv�X�d�Q�Sg�"�r�+%�3V��X�U)�<#���?S�6�g��.H�����f�5;o�,ឧ��X�o����͛7o޼y��͛7o޼y����sO�i�PF����p_<�>�/�O�i�Hf�_���8݄�ٰ+�_�$�ܻ�HT�f���u�{�@�w����D�a�t�nقG` �N�V�23ނ�g� x8CrI<�~�5�P�@x���[qJ��w�O�1u���猳���?!K٧3Α��(LSD�;�l	��.Дet�飂�����F�͸z�l�=���£օe4���><��U!T��
�BC��m�X�/1%,�<�V�%B���I�=��پ.�X�*�՛B��ɶ�+d�pO�'����z��c;R-<D��vM��u(hj����w��އ��YB9]�y3N���W�NI���/P��+�Z��a�\j]t���]l/�e�$֨	Im�<��W���V���w	}>��֖�܂�ڏ�F�(������ܤ���η������W�"�j����tz������:<��=�{{{�gW��.�\���o����|���Ir��V�p}v��K�ehYh{?ciϟ��z�O�&�$ӳZt�D����9MPLneC�� $^ϯ�̭�������� �q�o
͛F[�3=�z���5[Z�	�~
ϻ�B�!!	�}����_�ߏv��
��\�$�X!P4|懄Fh��L �l�_K�%���%��5�h��e-K�%駖��E~����c���˽���l����i䥉�Cn&�ֿ<����'3�w�J�s��8�j��/�/J[�$�j_�1ʸ��������d�ǔ���M>��k�}�v]��)c%
W<�H�E�?#8���~a��{�����J�.V`P���4\�B�)�o�{��w%���Z�%�M)o�'t|��}��ӿ㽭d4�0��5WlT��yWg߆K�)���5�	ڕ1�����?4���KYՄ� =�ɽ�a$�{ �7廪M�2�����&4�Gc~��Q����U���;�H}��Q���hF?2�zy�(�/y=�b=k� 񺬕+$]9ބ�!�e�40z2����}�گ��;P��-?�Ƚ�"�.>w|��P��_��>o޼y��͛7o޼y��͛7o�^˝�[4Jg�A����n�~�h�������1t�5�J����8��e&��h�}�;߉Ӄ]�&�V���B�52C���ޏSzm����߸!��|��J>k��4@�0��C�h�3��>��Q����S���o�'Q�?�L4��o�f�ko�.��42�Y6�&�7�˙���PR���Tg^Ȓ~; ݜ�5�F��3%�tԠ:���;��gᒕ�F �&�Sh����ࡪTI�����x����kcC�˨�G���D�ofS�?���<�e�m�_����i킚^�������vv�-���c�����5@@*�2���zw;��/_b�+?��L��R{d�@�v�����8I���Z�~Ch V�h��qC�P�Y��q��>�|4qF#��0d=�ҳ�&���+U�3���?�ǉ,�}h�|��t�m_{O��}h�#)IRq�d��gz�����x���q���̣G�`��)�C$y]�5p=n²mj����䍶����d��u��)9k��n�h&��n�I��g;�|wv�=�P����^�~��Q袊�tG�o��#���B֯��߳cr�.y��� �Գ꒑����$�H;��7���o�|���X���[���;��?�ӏ�>�~32"����/INC���}����Lf��%������_�F]��:���(x�E���ZV�l��R�b�Ϣ�Uϊ����?�.�����x�˝���/����k�c{QѤ���T��,�L"�}/8>ȫ�c�s�GR�U�xD5p�%��5�D�j�r<��� �٨������M��]��^�R����o�̻zM�Cd]o��6�b��5�o��r�Ns�p���LQ
�������د���+KXiT�J�:�֮��|���)�;C��؞��7��{�������vkk�~*��zS,q��vL��)��_��G�v�K�q��Tc P�/r�%��R����Sp���Ͽ/֟.��)�4�擁lg$���\G=�vR��	5ڡa�����BNCF}��aƌr\<7�m��~߻'�{_z�ϛ7o޼y��͛7o޼y��͛�W�2'�t&ެ��@�<D4��>C�@D���&��{o~-N���7N?��'q��G��y�"���-�ޱs�GР���!�"�~��8��@����m���.5�����h�q�8!�0��hr��3�+}hu��ƕ�8�����Wq?����Lyjy3����jJl�-t=�V�(E����gW7���$哧�a=�H���xfP
(e�_ O@����ǈ��zu�O�_���< o+R�5
X�DIdː|�:��O�F��#Y�U����6���$�*����A��F���O�;���}�D�䣡QG����D-jk��>kU9�`,Ej�Ex.Mh��QF*=���RMRF�e�2jFУJ�ْ�Poc]HF}h�0Z1��%S�8:י��|"�����Y�ёr��B�=�2��vڊ�V:��}���\۔~rO5=]|N?��ǲ?��6sj���S��bש!�a�89� Y/���{���9�Z�6�v�"��3�1d5���L��l���f"��@�S�Qw���u5��ciwmA������O�@o]������[��Q�]��+	/H�,�q�FZ���b�������}�ڭ8�/��cO��7~F�	' ����)C��Z}�� 6�gՄ�z_gi��y�%͢,O�������je#?ί�M�2���Ȳ�j���K��rzQX�uu{�l�m�|��d�XGg$��Ym�m���ڎ/ݖ$W�~g}߱%AFK�s�>��/��n�������F�Ğ��Qy�u͕��@�>y%�H�2v<������Ƶ�.����ka�̕�7�H��^Yu��+�@�u0._Ÿ��ԭ�-��WQ�p���<�GI�x�pZ+kx7��[��+�̊3.���V�sO�M�P��?��E�[_�H�deE�	��0+L�`���"̩y��x���++#�����]�w��#oޒy��PʽV���O�$�v̧��h4�����aG�[�S�v�wC����rוz�����c�����<���^�}޼y��͛7o޼y��͛7o޼��;�g=C�Y�3�O��f��vDC��K|��o���w���@f��B��?�f�M4k��	x�Xȟ�O�:� ��_��8=d"xD9ZA���MYK|(3�����3/=7��j�Xr���S�.�cx:��y�5!q%������mB��,�Xk���3�e��?Խ�I�T4Bzr�Q�A��k�X,{_���(%P�tL��"n((��"���w	�����P@�'�̍ t�Zm�ـ��|�I�-����
C�����:|�Sx���OeD�lOd.;*�ث8ס�^@mhT�[8$��]�%�R,��@���
頇��ի�h�}z����Aj�Q�%�&*�n��{ r�����w(�y��7���������!�#x�����A`�(;���r����!��1�3���-F���a�5��`��&^m0z[褴�u!����$$�f<�F�-�N�8&��?��q��`�~��1��l���m/eh���yf�]����b3�=�|>Ծ�M#[�����:s=�I�w&�ܶ�a�y!uR��*��zF����ϠMD�J>�R1v���O�lo؅�E�_lyq��,)�����57�w�hA�,K���U�
�g��W�5�j{.K Z"�=��f��W��ug=����^��X��z �vYb>�}������2g��}|?��d�D�UD[=�6q��1z+I�
4�H�����W�$d��#�7��aYߔru�����ʮ�ܨ�3%�eFb���s$�T���F��V�5��I^o��.�'�/�d?~O\�&��\i��t�.j"�q�	�R��e|GLA�a<[�8ϡۓ��;I�k����������RȨ��{�|����{w|�)�S���OY_��ٮ���ff|5g���n���l6�z_bќ�ZyN\h`eZ���uz�g�bn�"D��|���wX���P��O���AS�ۓ�A�K	?������j{�ﱌ��َ{q�o޼y��͛7o޼y��͛7o޼}�-5їx����3�Ch�>"����^�5ό�����^����|^ٸ�?�sߊӓ#�y9��wdm5��~����M{��$N�߸��D���hb]�"�)U\Ҥ����p��2�ZfT�	~+�(�Ae:��W���,I>�c�0|��~9N���������t^m��fQ�G k�����x���!��^E�HO�A�D���7̅��q=�S�K�Mv��Ӏ��X<\�c��԰���jBM����L5?�iPQH��3e��Z}�|l�W�|�~�*�@�>9��ishxL�a����eI�M��'>�~xF�-9�u$
��2���:FC��CR���2F3�b�C��:<�$�V=�|U�P��J>�8/��u!�N���j��c[�tU<�	�� ��l/���*����G#!D��,_�r��ב�bt4%��|ݗ"FE���$4I@%��/֡�8��i��h��z�=D+�K`�M�U	���Q�3�Jk{I��Mօ`��V�1$c�	,�E�� =�%�����J��N�9��e���_`-��?X͞lbc>ٕ�t6�{4��$?$@e����S�#�c�����d�1�����ԁm<�EK����Eɗ<�ts��Y���좖�����,��E�e4i��m>��w�|fE�[���oY�3g�Sϛ-�yz�J����3M�Ώ����g��l�YQ��_� ��O�~Ny�i��Md�>��!�l=]�s ������:ݢdi�&����:��e~��y�:����q+M�h�a<M�-4+a��������8�x���p��A���S����a�*��K����H�qE�QOH��umD���@ �ѐ��b%���+Q�@7!���!���H�6d\S��(Tmp�VDMh�N����qEI)�q����2� qW���:�WJ�,A�
�����\���[���3���qHmtVV'��e��M�A�1�K54���~>Տ�D��x1g[T�8k��<�՟���߳<�;����h��
�^��>�)k3���+�{�FR�(�[�n�*K�x�)+H�ҳW�vu4��'}�>��u����}�-'��
����s��<�
�>޼y��͛7o޼y��͛7o޼y��[�D����3���2Cy�޽8C����DS��W���e���|c�������w��)����}�V��д�ф6_Dϣm��y�k��i�	j���
i8�Z�*���H{'�L�{��}s�$ ���.EU@!�ꤏ(�Զ��sr"3�-DY��4Y�,/j�Y%:�QjO'<2�c5`p X��QQ3�Q>I�$����Efm{�6Nn9��5�����y���3D����П}��F����b��!%5�fW�D�z`�>T�N+�fX����F��M<a����\E{�a$혽�@<\�ڨ@�bjD�c4�D+0r��(���O�'�Qc��r6���5hi��yY��4FW���w��W��>鷊�b���P�%��%x4� �����r aG+��Q�]2l �N�BPoH�1��Cz�֠�������u9?5^v��z�Dv�	��V��X~uDw���-���B��|��RS�$a�?0Q�T����%��˒�[J���i�o~?�h^��o��K��UԣF��=��O�H5�����R�E����je�����#q���o�h�)�_,�8x$G�,��ԛRN��a���]�sp.�����o��6�(q��Q��B!�EVe|vKi��#��s�x�fm�E��'śd��w��Y��˞��8��%�.��[Բȍ�(�)���.��E3��b��&L#��j6�xr���������G?�"w<�x;E}�{��w�8s�GR��}�ǁȇ!ᕸ��E^�$ �E�;�}�yYV�Ԡ��Z����1��g��l=c)���S#��v���m��	V�q����2�7�9N�<��@Z�+��w�c_�������v���g9��a^�J)��#�������^m�I}�@:2Z~�}��8��P^$�Hx2�0�D��)VD�J@���J.�l��nώ��?��e���~��63;�J���8�[�8�;=oރZ�\!����Z�f԰�s���Xg4^���ѧ1^e,�.㻿�z�D=_A=-��;	Q�O�|ؓ�3j����﹒j>J�bs)reP��*��$�r�D�7o޼y��͛7o޼y��͛7o��=7�g<ϊ�!13���?Bɽ]�2���}�8]k1Ra&�-�mS�{M�K�/���d��ۏ�t	$T� ����G��kW�: ��@K��5֍��ꀄ(��5a�S7j*g���Ӑ%�|S��<��զ䳇������g%(��p=���<���C6Iy��Ԋ��H�A��K��H�\�IXOZ�`kqY��KO�T���q=I$�H�����͍�f]"�e�¥��֍[q���������$� ����ߏ�>���mwe5�폞8�W41��[,�D����������z�5!����qZ�G���(ɤZ�7�y&SF�O� ���ᬀ8��
�Wӳ6�s����5F7O(7����£{�!�YO*�j�F �������(~x�!��w� �lIr��"=i�a�zTLP�8)��N�f�g�4�W$�X�-h2��p��u�?����e+mٯ�o뎔_w*z($d�g�mh�e��=BهF�d���Ӳ�P���h���h��d��j ⽄�E��m���0=�3C�cY߬N3m'�
��������M�m����$Kh���j�zry4���v_j02�j�&�I�_���b�l_���"a&�r�eݿ�d�|Oz���E���PT09vV��Ek0�W;�H�<�ƒj�f{Ě��}V���Y��ޏnX0?�V�`���9����Z2�P��%���D{�$߂fo��g�}���)��kN��x�����ֻ�bm穬��Mdܵ��.3j+������:�F/���Pq~�SSyؗ�+eF��?W�L����+WX0��Q˹��H�a�P��c�;5�H2��X	8��1���	�7ǭ���N���ܥ��6�v�~(��?���~7k}����( ��<��P�}�j2��F ��͸�ߙ�;W
�4Ҩ��=���`�q�X\��_��Wq:$�W�u�߭Q��Z�S3^�x	�_�B$w�X��hʉf��z61,X����+�ynUdE�%�7W��lI>N�A�{,�i���E����\��ʘ��	I����D�7o޼y��͛7o޼y��͛7o��-=�73цH��X[���W�D*N@!�^���D�H@c��H�>� ?��4�����;��>̓K�&�nI>�@2PQVZ �&=!|���}��fn�_��������b�&fr/�I�߻�2c;�X*��g�\���\ʣ�`W�Z���E�X^]�Eg�OtLI����saЍKB�%����gy�aH&�Ɇ6�����M���D�U��h���;ӟ-�����G�[W��������Za�q=�w�_{������7���O~��o���� �5��Aҋ���-����($�}F��9�v���a3zа?���7��C�O�a�s5P��h'$�@j��ǆ�u5jC�G�Nzz4|��/��H������kc;����ҞO��i}�/�	<~ͺlk������1���P�)�:C��LM)�������Q��'��|4�#j���\Hd�3Ws��|�=B����qZ�F���ޑ������3�x�����0��)U$�/�c`��fjz�Ϊ-�eE���t�%D�bTc��4M2EdZ3�i�6W�/�HH[m����_�%Q�%��3�p�L?�r����r�ӳ�����	4�t� ����'�óN�v����-*��>�$�g�}��X�&�����;��i��[FhI�D��s|^y�E)^X�xA4*K�'��g�M�l;��dE��"��v�Ϫ�yfO��)2��Ek㝙 ��b\��wV�����<m�<�Ӭ�,����-F��$��@���I��a�S�a�{�}?NU���a�d�Vd�UD>8�+a%���j�}rwŊ���{+�6#�$��{�?����~�$���;��b����ue�Xq�N1�
���idV��R��>'��$2�Ps�7��9>&I61��o��{���o $jV6�h	�-!��}X�jGg�7]�>+��>�����~��~���?��8=*��.���>\��L]Y����_|ΦM-��{O�;�s�TѰh�-����|/7�/$+��:�o�!��֣F�%�'��D�7o޼y��͛7o޼y��͛7o��-=�G�>�5�0þ�^i��5D�mb�2c&$�`,���$+\��3���\�$k�{}�(p��Q$��D��hڇf�+B޴��I�
ȋ��O'�O�\Y[�L�̬!?������3ę��=!\��.�j���Q^ZuGMD��tF�s),c渚G�!Πs���k� 6�jcS4��-�?{;�\������5��8s}�4�KM��3�3	�r������?�F%�ަt����̺Kȅ��K��AG��7��ߊ�_z�;q��H4�����qU9��Cр+Q�}W7����������������_�鿏��:�k����͐�VÐ�nsK����'Ҟ�3�k�4��F��hR�m�v���A�h��;��]-�2�o!î�h�Zji����%FG��_`��֨�)�G�nǡ�o������_X���t�ݗ�r?�64$�J�M�
�D�2���4$x�K�K� ��>�Ix��}W3��)�c9 y��[o�i]IKԟ�d��i��x���D�E�{��6�m8�U��S���K2s�ȐJ������cTf��Yb%��;+Jt2*�Z���2jSMH�+Ige�����1E��JIR�R��ᾐK����=igk�?,�m[{[J^��!w�<��-��=�c6�uCDS���SF�{��)�c�xB�."5�N��t��킋����^U�*�<��e��`�u�����,� |Q�+�@�z��ɘ$�O��xӿ)����.���$K����`W��1�<<�(��:���d�X�v]+n8�X_�D>A��]N����ŕRJ��
��KnjR�"5��,h��\����o�<	>�p�V;�� sYϗ�c\��P	+����.��i)�;Ǖ[�<����8~7��F9YC�UL���;ɱJ��r.����?�[������u2�a�3���i`�l�'�튂t���	k�a�v�D9v�_�#�+�=�<�z2E+��3i���(��M<_j��H����)�aT���2?�*Is�-�����͛7o޼y��͛7o޼y����܉��LX��1ƌ�ɱ#îO�Eȏ�64�F2�VҊj�o�'F��R�%W&�w�qJb���{q��;B2���?}"���{��P�Ĵ�,z�#̜_�,Q{#�?!�����RIQIQNS3S�)�[�,���~A��F��ܚE")�2R�p�׎H̝�N֬�dy�����<"�Q���Ѿ��G{�{R��ZB��N�I���U����W��xԷ��g�ܵ��n��[�A�����1��x	���ܔ=J�!x¾��o��w��O�����ߍ�?���[j@3�� A�0=z,��
��U!�~��B�{?'�}�������D��U*��U�,6� ['�%��� �X^]h���SMFE�!iVTH(<w�e�k�h�m����Qt��Ք#r�0v;�o��P�6�g�d�P�~}FՆ'�,岲&�\j�2�Ɩ�cD+.S����Z��&�߻�%Dsbo6�&��7�ڮ@󎚇$ iͶ?0$_я��z����ξ��I*B�R��6�7Z���Sor�r��H�]��j��h�F�/<s���9D����K�)�13Z#XL<�_�je�C�����ϲ\5}��JR;��ߏ���~FF��`i8磱޲]_G9��>���������~QB{�
�E/N��b?K�50�i���_�槽�JKʗQgv����>�Ym��*�eɩe���I������g�$j���\6�p���Ӗ%�lYM>���e6��^'7�}��E�������7@lE�x��)�߮@����ɱ�,����t��%���,��z�Wx�{o8������"�oa&�u�-����ZxvŁ[0E��I��Bj9�8r��L�+|0NN4���QB3V4d�W���9�X��v3�Lׯ���$˸ e��\$����\Ɇ�VC�`���
�PR�D�c{���|�lW��3�c4�#���jV&�>ܿ�����̃
2��v��Y�,'���<��&�ȴ/�IEUW�g�=�_��c=��������y�;Q3D�3�w"5���^7ןbJo2�Z�����͛7o޼y��͛7o޼y�����D_�3�k�c)��Ɗ�+�Ȝ��B�y.��CT#F�!)��.��AS<W�\u�A���D�&��Д���(>�GB�4"9�y�2���*P3��T�3���\��wW4���l��}�7�ɝr�Zo\���y$_�e�fF����3�T�
Y�l�S!�e6A� z��x�zȬFAH=�.�FZ� j�œV���oܒ蟌��^�\� D홢����[�rN�?��QR��*�)<?���7�tg(�_��/㴼R�R�Z!�}��ãT+���O���>�Q�����r�������o>z?N+��3���D���C�4��3�����#q�PS��c�xϥ�s�X��GB�l�)���y��m����'��F�b���mJ?E������+rw<���-�#�N����|'ڐn9'�����A��A6уC��h�Dy=��r%qI��	-��Cmj��\����Z��<<�v�����K�V�x��ٽGr^h��ZҾ��\�����G""�~��Ly���I���ډ$��e�|gFkw=�J�[�tr���i��c9EK�v�t𦂝�T=�J
���'G 0��D�����$�����E�kA�h6��^�*<�!��"��1�K�͌���fY��(�d��&�|5��je�q$��tsC��CDϞm�e��QD/����Y�m
Y��b���Z~�:!�w�E�n������gg��{�������5��Y���hة�zA폥J���}�n�ԇ���Z�'Ъ_���>�gK%�o�9tп�zЪ�Rc�^i��cG��T|G�F5��3�!!�I`��d�@ ''[��O���|�����R�������3�6�̜?��|T2�8�%�$cv�c�{���J/�3&X�DԠ�9��v7���75����X�|�]�1�������}�� tv��L�S3��]�m��(����w���X.5q_Ԥ4d���3�>%Xq���c��Wv5��޹Ґ���U��*\�WX�L�e�'�^��v��2f�G�s�J~'sel��ƾ�y<��͛7o޼y��͛7o޼y����+`��>jr� gB'XK�(�ux��5�܂ā�",���p�.F�a�J�p3*+����#̴���"�5�ۏ����n�%[��ft�*��QiB��[Jp�6g�1��AP����ߜ!fi���;q�ᶐU��C�Hg�Q�����b�/c��Tt����~\ZS��H�{�V�����!�g�_I��οc>�JUʹR+:��m :)���CFɒ�+��r<2}h�a��F�T���$eT����+���x 1�z�AZ�Ģ�CӍ2��UA�8i7F�z��W����u�V3,�kA;���><j��P�Q2I>����.5E�cj[#�i�gK5/A�Qˏ�ԏ��w���hF�rE��Z*yѫ�y!�Bji����I�C�Z�c��|#N�W3��:�FF����p��:	�Cx$i|Ԍ���I���(�М��C���?�B��kB� �� iz:��x�;qz���#<'��Zg4]�Wj^�<�J����V����~�薸c��	�'lOM�m����H�N���PT�Q���©�0(e���qKzs=����܂!^2=��|3�U�ѼG��]'�s_\��U�q���L�ZW�o<���d�h���F΋�{^�kQm-K����mc|D�Pj�Yr/�������Z���
���C��F/>_y�U#���c�E��󒬖�*�~9k�/����ĳ��쨻��g%��k�%�R��v��F#�D��=t�n�w5z*����N4�d9�;9�EV��b@U����8��x�$_�'�ٿ��w0��A	Z��:������3�/����74��MeW��q>�JF{_�ϔ(�ߎ
�:e�~�f����@A˗1	�̵&J�U�d��F��YD��1�?aF?��H�����j$�^㻂ϑ�|��K~�;	U�[%J͓�wYP�����F���cHΕK�������Wl�h}ە.�ǕZe]X�V �7q��q��3���u��a|����A}�B�����^�,�����yo޼y��͛7o޼y��͛7o޼}魜�9��Ud�r҃�:�1�!��Gx�ZY����)SͲ����7o�6�3�'�D�[)̸�A[���ZS�#qS�����^�d	�7�Xi��������#�A�F����9��Z��ߺ|�%����⩦�|�K���Ad�K���dsMʣ�����3�~���	i��4�F¨�D-7D{.��!D�4�������� ����e���s�n�:�.���[�jC9U&�U���WChU�A���?�������=* ���)�O��G��[=�tP�8��"�&C���`��P���'�9����;B�iV�Um�ㅨ���~=N��E���`�$O��*y^�$5��2NH�����iVo
���6�8�q���z /���~G��+�\%Z0�]5Ou�ͽZ�:��lZ�=�?$
�4c4݃}�RNR�M/�TI�[I;]���_F]�"j��Op�8S{�#d�{���8ݾ'�}�M��@MBh�L�a�~�a�K=��|���V�����f4>����VC=�G�҆hp��:8�zȨqV�E�a������|���؜�:t�qٱ�Vʃ��l�g)��E.Bh��0K4yC��Q�kóNr�Q�َZ-�<�����v8p�&���amQ��$KW0�"�G��Dc��ޱ�<c�Q�oh��Eɠ�j���l:k~�E	�/�-���yi*.m5�l;+���7Zm��^�x��d��ϲva�5�GIy���b��^� ��V�e�,#����KX1TCztx/N�w��)W�I�c��nC�㭈�w#w�,��񡨀�-W��h�`~�s�G"��P]q1u��r\>5�C�r�,��e�EdS��f������u��>�+YO8^)���Zz7j���bMS���ҩǅ��$��ȨE�+�ٟ+v�{�Է���߁C<׃Y����!�����c��㉖|ϭ��;���vS�Mh_�|j�������s���ѿ�q�[nq��Dj���#�2�/ʽ�V`�;k:�V̄tg�"��y5��F۵�L��ߟE%;qLB��͛7o޼y��͛7o޼y��͛�/�͙�N���i���N]�@�A�h4����� a�.Ȼ	HjQ�?B�2���Q=1z�����Zg�Z\~����kg�u��3��Y��qƲ�k��><6[��К�#4�H>��J�G5xr��)7ײf��=���e;N^�Ǜ�\���������ߋ������8���?NIL�B;h�h�$l��B#��$J���D�zD(���x �1X'���R�/k�~B����|����������߈�Z ���� �}G4�n�%���M��ww=���Q`����ǵk��/RS���pcr���xl���D-F�"iF���r��K�S�+��ޮ��g�B޼}'N�}G���
aF��G�E��Zio��Z�%�M�C���=�s~5�A�g���iT,`'�c�Wʇ��KW/�)�:o?��E��$p?D�\z��muM<`�Ֆ��՛��tO����@��P�ǒ�4�Xn���|�]F�En_E�H-�Iѝ��E�#y�%�������R{,o��*MZr�=z��ٚ��JĖ]b�$`�hh�ެ�ĥ�dч� J�j� v���	��jFO�Ѡ���D���W�9+��7�3o=�y�6䖨I�o����M�""eY�-�c��v���hK�|�7��h����Z7x�ch�p;WL�Qҳl���o�}������c���g�E��*����ɱ�jѬ'���Ec���  ��IDATP����˲/�}���>��}_/*Z�E_�E���O��~Q��~��@����Uj)Og��HDI?X�P�ԍ��nK�<�8��ç8�|�c�����J��E�;%�֙��H�S4�W����ҞE�Ӂ;�qO�Z��
����W�Ԟ�y����]�l3d�~���"��롫	G�8�3�����{\�E->W��*�3�V;�I�&]�`�-��.����$ǣc��������L�Vd�?�8E���w(�gSk~6s��<�+&�X�6f9s�e�5WӯT�O�ђ���ܿs�*�!�%���������9$_��g�L�4�|��\�����~�̀'��y��͛7o޼y��͛7o޼y{�'�8�k~c��Z��Um#3���.����W0��l'N�M�l0z�x�{�n�Y�
�M��Y3�(I�XR��u���w��A���s<׼3jJDcX����}�j(o�s_r5�
��h��x�J9^���+&��df�1c~疐k�X~O���rY�j[��w�F
�P�@EL>Y_�1 	řr�n�G�/z䲌�9�j�! ���$�����q���࿋ӟ|�I��v�V�6
 �F��'��:�J��~�����_��e���U�۬ �n�
a�}h�$�uf<m8"��F���W������!�n߸�G�ں��o��?���;O%ߗ�_s�φ�D�F�j�-G�@�P���č:����<�V���1�k�Թ�h}� �y�s=Fa>�ҏ��M�{$��SVC������\��U��Ctt}Sj���^]�y��'�ڂ�
��6@+�~D՚��z]�d��%�W�dQ+�8�F�=��2��l��>Qɒs\d�A4dxV�.I9�K}$�}��<���<�4t�̱<��̮F�EX�'��q��9K#m����̛O|E��e�d�4��ɗFg}-iyŖ��V��+55��<5�g��(M���}R���cb�	g����,�u�~��2�ﱳj����/JP}��/�-���w�E��H���(����h��i/^4ٗu�^_7��q�������7�%�B�o?����_Q�u:&�����'�vے��>׼~�bbV����!��������7��>gWK.�W�s��R%�іZ�`V e]7�ts߯%��Uˍ���v�{Ғy$�JVr%���H��WR���#)Ȩ��3��Q���,��HVH��}]�v��sv3���Sw%�,t�Wm?�]^�����p$�Q�
� �ҘQ�e|��F1�V{F��r�d�j���6�;���|[���kj���f��5��}޼y��͛7o޼y��͛7o޼���D��h�k����$�8s��$�4zf�Q�dF��B�R��jQ$���m][�#\���d
5��tscù?��4΀�z��H����!���o�+ d�2��'(D�\iyI�,�,�ϵ�ڌ���~E9\Ÿ/��{�����y^����OH>�s�\���J�WDM/xV=���L]R��D�k4���̏�J���RA�������������8��Wޕ����g�{,�peE����?�/q��Lz��a�����+��<,>x��	I)��8u��&.<����h?$hIH1�n��
����H�%�F��kw�����'�ل�	���X��`$��]��oQ��T�'	�*�<؏%���X�牞3��ݧB���%K/�zɨp��⡫C{�Ү�(�m�o$��wQ�����`<�4	����D��6��V��lWu��i2�ǹ�3-X�,
������ձ���D_��Xx^U#�C-��K�J��b`��'��s��]B��Z�[�|i����3�fh��]?���=�$�":�)}�z5� _��Kj��|��
��"�۶Qt5Z\�wV�q40���G4p�s�~_ѵ(�w��v���:�E�g�g��������_4i�}�eii.z��T�[�_����LK�o	4�D�`�1+P�L��Ή��z ��=υ:^���j\����Fh��P:(�J��K�6���bd�5u׎?���n�}o��2��(��O���̾�2cQK}�f����h��S�R���Y5�Di-��Ն�8��3k��R�O���d�����W6�=��0B��C�Ty��q��2��`�"r��~/�*�}��D蟶.Mq	�J��sh��{��qĬ�~/E�����3���2Ғz,��H������~��>���G����x�q�;;��VrH�,�:�Ҧ����z�ϛ7o޼y��͛7o޼y��͛�W��FiNt����UD-<ܖ��=�ƻqC��Fm�9=Q2�a�mG��2�\�ZwxV�q�uV��3���Ԭ:�|EJx�D�f|�|E��lc&��%E��������Z�,(j��&r|Ț�Z}�6�wSˌ~�1ӛL4G���L���S�y?�%�� ���'R�o�.�u]��1<g��n���z�"d}�:����k�%7ڡ��cɅ�B�v:���f����K�����r?��K�nn�������8��?��R7_����(�$���!���p~�������㴌�����rxZV��&��"�HFF�b�"�h�
��c�2GRԊ�u�������Hh��#�4ECI�@������V�Jy�@*{r�)�9	*E��!��zN�%��n�|�ֆ6C>��$��_$Y�
I�	4)��T1��O+i��8��@{������U\_��h��e�*:E2@]�l+����'j���.�GM�*��v���)�� �*�=�$��~n"
�����B���+��;��B� Y߫�읹��(S����y5�r�9�M�4��$��?X0���2��z�ױ���ni2ǲ���qE�e	>�~T��%Phg%�x>�{�Nd��\�`I�e�!k/�l�&��5ٖ���>=+��,��e��[�.��<o;���}o,Y�Қ�L�~Ҟ�5�'��*��|�-���hc�0ʸ�-��%~oθBƐ6����x-�d�sj5���|^|�f���}���;%������N%u��U?���CC�g�|��i4Z+�?j�a�*ޗUj�+�2r2snK��ϕ$_�+ߝ'����y"+�>|�����7�I���g�\G>�^7��\�J�>c��ήhP�F�=6K>P,�fK��ļF�8i�-o`�6V:Ҹb�N�nF�m)?�M1b���I=��p���=�;�z�F���F��2�ǖk���'��y��͛7o޼y��͛7o޼y{,=�g��9�H�gLR��j
�ߏ@���*4�� ��=5�v��[�uK�K�d��v��gq��o�~��%�wQ;�2!P�A��e�f���Wdѵ�BX�@j�����r_��ǹT�׾j��P. Ѩ-P8����e�}����e=xa�#�(V��d��ܸ.���n�����K����%�h ��r��A�M'Ԑ`4Xj�9�Qm-�Ds˝��4��/��o]E�ۑ���nY�l}K�G�)�k�1Q���9�o�C����u��Г4�������J��Ӈ�dׯ�Ư���@<?���?�����P����'+>���Z*�1զ���+���hM����^Q�����N��\�ѹy�Α�_��h�V�@=������9<�p	��\3������ի���0j�
H�)<WCD�ըȌfk�����5w���� �|���}�We?F���GlwP�~[�@m���U��Lt6j�$�Eٹn	Q�TKG���h���9@�Nr2���
M��D�3�G��-�Ǩ¨i��������x�g$LrɈ��)�ϒ�����RJ���u���G/�0YV2��ig�^��ֻ���u������Z�/0��EVe_T����}�b��������S??_�ba��տe�ų��j�����z}\����~��]�q����ߗq��tḶ��?	>�37�g r(�&�o|�SK��)VX�ge^t���L�Dj]�&3��<�9��E�|r.�4��񇓭d�����#t�h>ї&�J��|�t�3<���e%�\❚�I9��Es}���x����da���8�������8w���VS��o��N����W�R���F}�#�K2u2��C����=�ɟȊ��?������� �++��M��+����l#�/�X^,g�~?T*�6�jp�{���$��bi����©���#�<8>�.A>�UO�D�TJ*v��&�� lO$�h�K]�}޼y��͛7o޼y��͛7o޼�VNjpf�D�53��8����;x��ߋ�[�o��\��j�F�a�Z��("*�FS�5�@�*��ܽ]�P��-�!����g~8�˵���h�nάo :&5kx=��ł;�� J�̰Kf�5������L�	g�Qc������a���$@A���X}����(�$f�f�V���
F��h)F'ZG��RY�wt$��Z{hq�D�N�~L YU�J������8��o}]�c
�n�tw���+M�����I}����qz���pr�D��?���l�c�t5�H`�cE #�������ڛ�Ax�]�.��&�V�%�x~�T�VU,�'�؞/L;�ŔU,����4�z�p=iG�)K<��?z3N�����lgh�R�9��I,����������QB5�����@�iů�ħ��f^O����A��C^+I?�h�㾼?��ݍ���[_�g�$d�5����|+�d�s'�%��[�u�}wY�O�-O'6,y�wޔ�\���fi�\��hm={�5}-I�-klol��&��0���j�0�X|��E#�����w�Z�@_�@��@lQm�u8�$��=/�u����P�w�2.�⊂
V$��/��ha<����))W*M�wqB�����'��\�M��㌬(���_�-[oR{�ax���G&$�#C�ao~��;��ߣ$���G�r)����H����@��B�=�� N{'��彼Ҕ��b�쫢m�ޒ�24�k�&�G�;<D,��1��#h�_ڔ��w�yO�7D����H�H�vO�����i��<�'��dW�mH>[m���c�B�+~��?����BF�<8?���b�L��?Ew��^�ߙ���)�v���F_^��L��h�D�7o޼y��͛7o޼y��͛7o��͙��L$g���Ho޺��U���d�����m�0�2cZ�����it#DW�Z�nWf�9�N����R3�ͥ0tgx91��uh0Q��z&��B3�k�u��5�|�D3�fߓ'2�>���k�+u)�KW6����?K̼|�W��.w���x�:s�$�4��u��F߻?�Wt��$�q�oaF�{2�q\�?_��F$���ǟ�i�+�фQwA����Pd��r���m�����������H�A�=ױ���B3i|$���ץ|���}/N�|�-��#�����/��(��Km!q�5j(
���(�[��X�u��O�Y���@���Z��Q�G�*�!R0�6��c�[�7jՑ�Z�f����ǔg�z�K0�B�a�2V��s�f�DםOD�����F�SA�������f�f[l���8�J{L$��{��|�D)k�I���-Z'o|OȾD�g{N���f��G0����P��V,�ԣ^Q솏��3G#+Z챥��^�^ּ���t� ��/8���e��;�-KF��ǜd�?u������n6:&��"B^M��)��%��.z=kg����X��_��,��4�����I��\WQ+���I��"`Е��X�S��eV�&X��5�'%�Ǖv�A|�8?��K�ڳ�e�+��/���j�f���;*�v�O�qޢj�Ú~;4�"��b��>H�Ή|�lߕy��{2>-ER߮"FB��kU�� �n�G��"��h�_�z=NI�v����ۣ'O�~���~C�3+��}�X��;�#�B�2�>ړ��3��@��������A0n\�om*�Guh�{��9��>�*D-���.r^K�[�4TQ�ese�;��~� �%������ڢ5�ٟ�<��͛7o޼y��͛7o޼y����+`�L�ex>
�)nܐh�ב~�D���чqz���8}��7�t֗���H.}|(3�h�p�T�*le�Kv��"\�*������]3��K-����~�Xf���kj�p�d�ꪐF�O⏚g�H\>� '!�<ZO�$�j$}N��eMI�����y��ٗ��c��mY�젝{�<���z��{U�����Ճ��l�lc��@B	�0F���� 	���@X�n�ո��tW����՛�;�{��!�v~kE��r�����3�S�~8q2wfDdddLߊ����O�r��izʦ6q�b��B���jhK���`�R������zϐ��� $sP���0�2P5���������������.����[�������p��vRC��L�d
Y���1j�$��djcV*r��%�|�;w��ໝL��������M��Ih{3�١UBƮ�q]�u�Y��uC�S��d@%�R���<h>�y&L;�bt��,q#��$�\�=�B�Uv�`Γ��_���Kv^���#i��.�����J|mX(����~'�����vdz�R��b�;�)H�4Γ��G����m������7��ʫ�A���:R~�����eG�Q�C�\����ϫ���?/�>W��AF=I_?3I�˃�.�*�mLm�2���]�{\,�+��T3e��w��d:o���f������|�p�|g�����W�o�|��?g�T3|`��8ݞ0�Z[��}[������0s�;L9d���a�o�,�a?��u���e �݆ ;�	h�5�pA#S罓�q~�d�c+Mj�?f>I�����1>	��xW���;Qe��@捅���s��j.5E3�#�T�~aЗx��ѽ����w~(�1����G�*L��*}H�1B;�c�T�4$�*�5�zI����U,H~���[,`�Г��t�p8��e���/�'WCy�֊䓚�\���~H/���ӫu��+�	�/�:N�*�8��S��?whb����)�������]�FV;�b����3�<<<<<<<<<<<<<<<<<<���p�Y'���bi�F�{�?+�3�����g�|��8|㕟��e�D�ʒ.Wd�`���V���<8�w�:�t������>��s8��EX�����CXfj𚴱!{�ŋ��ڲm/j/0}zw��3-�c�[�++���0�T'���`A�Ĕ�SC1�������
3�6�������jSVؿ�K¬����:2:5�#�wC�ħ-3���~�\Ƣ0���hJ���B؁�hZJ0�xl���4���$8x$������8��_�W%�����O��8���Ϳͻ��PnJ�C�͋L��! �B3�0�F� S��1���lp��-��2�<z`���٫�f���Z��u1������k�W��Lbڬ��������s�Cbr0	�wTW���^r���0ti��¥�B9��9>��C����/�b��[�wڶ�u2�G��¢����,|F{GSL����O].�1���.�/z?�Z3�~�`�f"5J���%��v�i�%��!4:'l�H���Ejp�4�-�OȘ5LF2*�֌�ߢ��沄�E��̚f`dp�����g��1��b�ivf�wy{#f���,�Kj����#W�b e}g.�e�ͫ�vU4�fmW.JS/��ެx.��ޠ��ޚAS���#a��w���ơ��φ�g�1��QZ��睘o�����&dx�<*�Ζ��6_�4V���:������9Ta�1g��������@�����z.��'ǘ��#�{�SqЖ�E�����B����Douu٨#~���+�
�/��r��a�UP_ז���x�����:���~���a'#��K�uI���jM�-�fhԅ9�Ԓy��ޞ<(}����<y �C0��O���61�k�����@�c��'d�a#WA;�>����_�O��S�L�*aG��!����N
ӑ���^zF�������������������5�s�>�0�i�0�l�����'_/�{{�-a��r���%a�M�Ň=ܔ�"Yz��>�7P,��=�D�ro<����W��o܈Cj�FF�\d����Lzc�t$���V���Z�����eYK�6����g� r!����ڻ�F�
���/�N<���w�y;�o,�B;�!�����EƝ��l����1,30Hi� ������ށ�G-�	��@�-�$���ÿ�_��o�៾��8��?��8|����ʭM��h@HHm%�s~���P�4�4�\|qì���Q�#����+]�;0��͑���C�;[V�n�%vA8//��C'8��y�_������/Mm8���?xW~��d��͵e;b�7�ű���?_��z
c�sX��}Rt��NG��^�%��=0Ij��-ȣ~�4��G��h�Rˤd?�z��x#���1�z�-����}�u����Z��f�����Ee�-��p1"�їx�����^�^^��,�8��a��=0"f�Y�颵�R��/(�E���.�g����;/���{��|
�7��Mx�κ���H�w��J���O�-��~�[V���?���̗�1��΅h�j�W���X R�7'��?hmC���� 	���c�����P�ג�P$s��d���`>"j�M�`�a�7�BS��| �5a��ڼ�[��3�Vm!5hFd�I:��[�8���<��+w@6��`.�dG�3:`��aݣ3��z��0�lb��
v�q�YF�=y,���;;>o��ǲc�}�q��\w�d~����u���Z�qg�{�����vt֤�8���s���D{�:����y�@�w�������>�Ч�}��B�Cb����n�گ�j�������`L|g��q��,L����Lo���f�XVx{�ʒ�� W��� ��\��߹B݄Wē�[��!L��W˫�R��ʊ4�P�2]�J=��}�F�M+�#h�a彏���O�p�4�rL�/��wN�����,���N����ۢ���XV�����F�������6�WPz����$,U2^�IG��%���m�睎�3z�-A;��L8�%����/�n�q�qH�Ϳ����8��?��8\�!ڒ_��W�p-(#0�"��K�7]�e�Z���;���:|t$L�#0�8O�ff���\i�\�� �Pk5��wQp�j���+������������y?i��p��5s��R֫��rE�2�J�����85�a�:I:�4���Oj�ta�$� ��3��Ӗm�{R�qj�L��G����zZ���n2��6���=��Nk��u�5HK{�P)%0w\���k�ټ^k�+�6�)A�;5i�x�׻Lo��gSI���f0�w}`���[[]��������K��c�8��`�x⺴YZ}��̡�
�w�Fc���NFk�G���vc�H]c>V$�K1�
����"�Qj�-��K�,�>�<M����H��"����>���t���C�a��1�ܑ`�%�<�{����%Y'�<���^�-�V�e�Wo���'8�A���:����m����'�c-��T*��4��w��[���]�SE���x����a0W[2�^]��om�ά�_����^>�}���J����nr���w4�1O��r����w���+І3��W�i�.��ԡ-X�:�YV����LD6�%SWk;��]�	�0������	{��}� ��>��������&��~�S��k���8��o�q�����!������6��Nd���#9j q�u�fP�{�ai�L�\y'�J��{�יW^�$�O��Z�J�+������!,��#c�̫.��U9F����Wk@C�H7�O�X__颵;/T�P�����a�h?~�f�Wv��;��R���qa^3�qi�:��S��,�ԩ�����a��3_��W��_����eXF������O���^�J��QW���
���V>��b]N����g[��7Җ<N�bѡ�Z�K���)hp���h,�=͠gk���^K�Ƣ��p(���GT����sF�	!2��e��ζ���(����g�v���-a��,,7_y%���Q^�VO���""���(fZd7��|��/�����,�u�?qzcW�u)d0u]g�����\i!G9&�c�y9B0'��m��K��pL/i�c��(��H6��h��B�iy7�U�Kk.���Q�Z�;��e|6@�O�iv�3�X��y�z�z~�-�^�=�)����.��=9>��ϫ�5#�K����0��������3�s.��w�L��9c�ס��&�u���
����E��PB{i��J�OK�&}�yw����g}�.{��IF�o�߻��;Z��������|I>9P��0LKü��Ǚ�f����e�Op�F��z�^8B�0�)c	f�VMv�
~u�t*��-�_"j#S�Rj73�H��m������윫`����>�9V�,�1�[�]4���>�qA�3u������&
��O�W��J�L<�;m���X�)p���wlkY7�[xn�'ɴ����޴�䫔�?-�>0O0���[�8�k/�M���ұ�LB=NΚ��k��}� ΅>�Ϭ��Kxw�J.�}��ۿ)�!��}��q�g�o�����V�W�F�~`Z��B�
6��Rc�8Q,�"<Ԏ�"Ya&�jm��٫^Ǌ�꺬ds/7����~��a��?��/|�q��g>-�ay�P�W��\��S�0�Zy�yW~#eɘ���C1R�p���/�c#����i�zU}�?�cǇ�_�c�Ո����9}u��_ې�R���JU��ܓ�Q�`��:]<�M���"����ߎ����ߐ�ń�Ϳ��f�Uh�F
B1��'�;�������H�gL�HY�ʇ^������g(�G��l���Җx�wN핸\���wޱ<P��E�g�,f���x��p�����ɗ<�V��<��Jd��3�e/1ّ� ړ.4(���|z>�O�G_��z^&�C-K\2e��L6e4�}�D&��D���Z�ƻ--�F��;9���}"����h�<�'�j�6���âݨB[-^�䪰���,��=��)���_���z���N�ޞ�����|�]NZ[�5�1���uy>k}0�|���Δ�c韹C��./Mg���\�vޢ��&��|���~�:��qQ󁋟w�&?�N��}��"����aD/��aw��Ś��ṕ�����q��xL�� <�bι���;�Zv�#o��/a�0��{}"a�Mg4RXm�x��.n7��;3�߻y�*_�>D�7��2��0�"�G��Kq���w����7����mo�A�r`(�QS���e�e��s��տW�S�艬�t{����d�52�d޷ܔ�߹)���mYw	Qn�%y���<v�A�0�����HO�=��<��Iko�S[>2�>yN�Ϗ�D��Z�!�:��%K<���Pͻ��N/5NW;d��3���<<�������������������� �B_z%�^��`E���Lzs���-�FU�����8��D��Ք,��0
�K
5�h �T�y��
]`\��
hh�4����o������8<:��\aj���x>z�%/��r��Y��ɊpԐ�.��7B�5�d3>�8N�����s"��L�=� ��}��+�sZ8q���3�
��O��~�&��G��՛q��^�ɰ���xL�E���<Ȥ��B�왟G��83�ӱ- d���-E� �2Z���?�In,I���D���t�7��*f_bb@9���@=��!5�vE
�3?�Ų����;�#��2N�Eô�EU1t��L���~�E!/�V}?�Kc�^��X���h,��K-ڑ�`[��U��!��Ѩ���0�:`��v����vn��ϻ�Q8��sƁa�Ả���e����g?�1��j�if�^��ݻ8�����A�*5��~��250��`W����H,�W��3�w�,�6� ���zj��]p3tf�Ջ�n�1��忶���9n�zK�h��8Ť�����b�-��z���Y�O������@1��w@F���'2^�d9�`'Y��Tzu����71�����ǘK��kg�=��@t��V�����-H�Tk:��֡���]/�`z��0���]�q��Qfc�2c�Y�\�	p^v�����h"��]o�òX�x��@�Mc�G?��I����ĺLL��Cّ����h�v�������+@#��@��a}csE�zw�E��6�M��;4L<	����z�+�㰁�~(����̿wۅ����>2�-�'S����c��P��
�%Ǎ���CF_�8] ���R������y�H�g�}� e�⭼%�6��xU�Z"Ʉ���%Y��տ�kqH���#Z}?~W4����.m���&�����93+�'cYa]��s2���nV���H,׏	s�����x`aI��,+��h�ln���˟Fߓ���W�H�����Xɍ�7�;��(,���p�)��E/;[X���:����o�����������5y�{�{qH��!�e,"Ej�@Zz\aJƢ����Y/��$}z��[���&��;)w��z��hP�����q�ekKQk����jFRB�C:`�~B,*�Ɗf�߶ �jG^C��a�2 aI+��Zf�T�sb���F�h_XK�%��PvöP'_���lZSNg���b��x1��� ��Xy�M1�24��7�����b����n��@�>���`�d0q���G�L��Ez�5��OFz4��o^MMv�N��G�p;uh V���W.-4}~&u�߳�ON�٪�yZ/gfhf���j>-��U�^�𩀡���b]w|$�HF?�s�����8��h���q�}���7������Kk��%.�[��v������=�͋tr̿����B2�j�����R-�h/��DٴWl��|]��n6��<lm2j�e%g� ��<�x�2Q����8zw�rz���t&��F��Ck�r�tR��<�6�����F����8�J#�l��x��P���.l&_r�bŊ��I�_|L9�߶7;G���*a�+���5h�Q���#a�Q�:���Y��f��6|�`'e�����͠]]�뷶d~���x�d��K��m����.0H>ڇ2�� 5��2w�I:5䏌M��߻�"����K����P��ي���LE��h*����x��e1��g�yxxxxxxxxxxxxxxxxx\��=�\�v1 �w�S�HiPˈ��ZK���W���^�����8�M����O�!����/��ZU��sAz�=ԑ�����b�ʕd>0��	3ke^bVeŗ+���党(w�܎��PV��뒟^�Fv�;)�y �-czrX&��"zV�Ǭ�W@ˏ�g��dT�zT�;/�	���kR�O�6��>'?��h-��Ͻw�G��Þ��Y݈�͖h�ԗ$����l��T�� �ք+��i逅�2�|�[$�=������h�11ay���}ޛ����@��g��iQ����p0J8����0X0ʴ�M���\���Φ�N�FVQ1����E�����o�ę��|��N�����c[tS�/��B]�z�N^��hz��%Y�c2��2^Ŝu�ׇ����K�Ο.F�*g��q]��J�	�:��m1�}�����o�E�N ��:�ldh&L?��H#Ȭ��т���}L�2�6V��wW�\�F�^��)?)�ch�t���Y�Ȝ������G����9���Q�S3�Z`0���$c�וc̈́��C2���X]Y��c~�������U'���� Û����7�+?�E[��ɘ-VP;�T-[��~��X���(7����C��sGǵ�0Q^cSڙJC�d�!���%2�
*_�q�>�f��?�{q|>FSψ�����q)��
f`���)&9��Aiv
�������.Q兯4e�X/˺C�+�p^�C3-�t�� ��^���&��_���[�u�nC�������K��О�L���m���|!�W�XY^�߫�9�l�s����a���Ԝ��(�Mh�>�7�;�e���;�I<�»�!;��d�=�v� ��a_�gЗ�,!���\��F� ,-~��1�m�_�CùՒ�*jø�;Y�6Q�t�+V+��Ei�9�}� e�E\1+��n�풩T�X��p/��B�+��+��������Kм�����O��Qq��!{����Z_�V�)+�Eh���W�xnE/M4�+�`���^�.zk��osSү`�}Ɋ��`&��G���N�WB�saL>�%<Z�Eթᡴ�&$��2��E�ͻ�������A~���"���P����Ӓ��O�+���E� ,����
�$���K��K/K�ex����������'�V�'(�ZR�����w��8��_��v ����Xp���A�����������%p%����❲Dˣ�*X��]�,����׌?�r204#�g�ŗ�����$�,u���˯��e���c�F�$T�W�\�}��egO?�~W�G���3�f?o��;gHm�����,���� +3j�qGC��c�ܡ6��R\0��x
�� s�	/�dP;HkW������қ.���Lt������n�GF��x���Ei���X�h&�U��;_�,O�&g�x\������F`w3)�D[��#,�ǚ���=��C��if׌���Ɛ��ȡ!��X��f}}���2���U_���u^k�q�kYMg�^��C��l��$�� �3��C%�8�zE8�1摅H��
v��^������<R��!�c��%<8<��k����>���4i'��/ݹ���0魶��.4c�䣎��?�x�S��~�w���x$���ɞ��JQ����G�?C+���:�2���"��e�#��Y�#���r�#�ٔ���]*���	��M�E�ѧ���|�5�qn�8?-V��������������������p.����a�+��h@&Bd�%rŹT���q����qx�Ծ���qx���8| m��;7�p�Y֠Y��$+�ej�1?�@��yz�;F:�[n��=h64�e"��"��a~B��|nj ����B��ޤ�rM�.V$���7�[{�b\�*|�0��+^x�%��q��뤾|�W^EB����}ɮ�F[!�!���� �r�NG�?��:KE�|w�����q������/�q8���h(KT4��Y������[r���Q�(K�9�ϢL\9&�����/W�煅i�S����i����lN��=�t�}Y���2̟nw1�4Sۭ�4{#��)�B���<ǋ�a���+3B���:4e�d�a���%h���`?�<a�,�|�e克�t^�!��++2��7iz���\kF�[����4�4�{����ӻn�Ѱ�5ZH`,���pԃb�������Թb��U��sἽ���}w��S��~<�G�W0���֐�|������t�3�xAE�MM���+�D;�ϲ�-f�٬���{ty�]8�΂��]W���9��6�~N��0;�����w����3�"s=�g�u�Z���Bj����)����{���<��:��
��<�u��?�P�-�t�`�|���h���'$�a�=}"�5���Y�|(�X�<��r��n��<����c�#�w1�~�o�����@�##��c�*�r��j�Z}�z��(�wƝ%`�Q�C�O��J�����`3~��<�R�u��Zj�*%B�v�pǋ�Qc�:a��������������������ȽЧW�Ʉ
"{�ќ/��l"���C�.Ck��]a6ݸ%Zl��C�����&�g?��JHK,5o�%�J/x.&;\�-嫈�^�x�X\'`����o&�+�d���R<1��6�Iq���p�g��!A	Ȉ!��ha�#�i�kU:����!���X[��&&�/���A{[J껄�����&,/)ͣ��+��U`�{��Gq��'��X��mV�T�H.��w��+��|�l	�ޒ��E1������m�^.ْ?s��6ѫ���f<?o:���K4mNg����7�:m9O3� 2ۂ�S��C��gk5Ѳ<o|��\�y���6]�u��0+V�8�n�����!ǓG�~����#�N�/��ӚQ��n����Gf�``38�uF	�m��<}�����Ue�q�H��9���� ��Y��.�~�y���F�ߗfޕ*�9F�����+����o�dD%�8��M0���줲�)�2g�k���<��eu�J��h(��G/�(���^�Sߛ:������z�?!��sKX����1��9���;5Xu{�5�L��䗽��8܅��F�i]7�q��䧃�h��Z|�;ܶ�w��9�����#n��tL�1�mcUv�}��O��ʲ��TP.�v����.;��m��O����H�䛌�A�Z}r� F�~�dx0���d�/5D˟��פ��;��������������y�c�g�yxxxxxxxxxxxxxxxxx\̼Ч-`��gV4q6��}XЬ��	6�s�<�Po����ƶ��:�B&+��������{�M�T���@ov͆���+�N�B&��c\��\I/
��������0�Bm�8c|��Aʂ��AK�rF�5�E61��2ޗT7���dr��	�;-Z���۩�`��S{�<H�T�~3c�B���x��R���S��,�|��}����Q�}R�
��^5m�+��s¼��jD���L>��]��Gy��0ͨ�ȨbD�h�!mS(M������U�>/�ˤ;/d1���[[]��k��#c���&�}j�YGf^�+�S2�=z�.m>z�e�̟��#�����^,��;w��!���.��_4,�ٷh�I�/��������{ѽ麐��L>���rɰ��u2�8�O�2�l�z��y�-\���>�w�%���Bǎ�h�~-S�75Q�3���w�q�n�É�Y�]x?���_Li�1�0���&b50�*%x�3��pa�N�Wh���n�y����s�:�����ҏ��Ӏ^oQ_y�u�.��߈�#���u
F`��w�ߥeف��)��-�$[j	no��&�x<�f��O�X����=�#��RC��0�`�	c�׆��
w�B#�*���ܓ���Z��ch������*$Þ�*�� w&Xlmą���پ��Э�g�yxxxxxxxxxxxxxxxxx\̰�g��+�F���-c���#)�ő@cY҆��V�2[kʊt��L\��^l��b@��N���1W���b��#���Q,�
�@�`���/1�b�����P����g�4�RT<0��J�t�$�wg�/�<��q:���{��i�V��L;XFVVłQ��E%(���ޜ�,X@�QX�Ea -�,Dcx'����pn��EQ�fd�1����.��ꊧpA8_��ǋ�O�z�u3��2��5��1=�͇���rd,�&��U�ue�\5P��ZW���0hA{�T�>�"CN������>�3荏^x��7\2���t��C����X`� c�L���+��%a2����[Y^����N���}���|�Y�y��/�b^D�<�&�!l&����Zl.o�ZÏ�T��Ѿx1���M��LOm��ɼ��'ށ��ɬ/���rp��9��,'U~A0}~Ɲ�A��@QgĞ�'��vh��;�4��1�LN�dj�B�� �<����y#��
�o2�t����(z��Yj�J���8$3M�CL��ea����/��y2�ƨW#�350W��_ïV%�Q"����'��q_�V2��77�R�xc]�;O��Ư�`L���Ն�_�C��G��<?��j͞�3d��{3��!��:5�8�P;�\p9���3�<<<<<<<<<<<<<<<<<<��X�S8j��0�Z8
�aD�39MxLM��B����%�5
9	pQ`[�p�+�ƒ�o��vq�y1��u�b��
m?I��k_8��,_j;��`�X�-=��hK�T���c��L��:�ȫ�#�!��7���@���ϩ�3�U�υf�{~���������=0��Œ@���F���C��y�x�~��qxԕ�Ϟ�{�Z��|�����!�L�_�Fܙ�r��=�$�և�5���=f��U��i��u��E�p-��a�n#�\/r]�O�*��/:�*3q����8$ÍL|È����	� �|���:j�1��L^�#^t�̣��讯#�L拚dd(jF����-����p����kGCV:WU���p�����Ი|�Ү����`����ң�g[��\�v���J5TL6j�71��W�_�_L���=�|S�l7�&h��`��v p�w��q�q���=ɼ_���m�sH���
����/�����Fc{݁�yex{6ځLH����8�B���{���7 ��0�.��@����\�Wf?��)ZOM�jy��w��Wd�r�K��/ǆ�)������9�ãc��nm���}�[��|���nO}��;�oЃF_C������R�]��^x}�O�x���{��if��0�=����������������������})˹��M�$���	"j��m		C��왧Ɓ2݇)т��y��jˇ�00Z}��g�]��Iy�����Ɨh��g���2�02ܶ$�B�U�:]��h2(FgJ*!��Mχ�/�"��x2��D��ѢW<�Ч4~T9�1c�J���~+�5���w�������ܓ���e�DF⽹)^����ߋ�Z ������R�"_���jo���)�ĕ(���L��*δ�?�=��2��-qN���vjj:~���죳�wF���;n������M��k�n�P���J��bHeg���)M*G��I��i���cte!�� C��3�f�K��wvv��Gh��0���7�7��Lj �d��>x#�7@�gH�]�pɬ��'V���3+?Loks�ʇfظ@&b�a{߽(����h&�U�����b������$����?���f#�s��;g3*���k+s=7_1�^�N0�_��~0��Vk��Z�6�p �Ћh1�-���1�1��8�<���C�E�wqa�h�������we�!�z�#�����w�i�>�o�v<Y���O�s�(�TJӯ���M7,�15��(o�NR+���߇Gү�t����=a���7����2&�D��v�{�ݶ3F`�ٰ�引�%��Sˎץ�m�5t酷f#+�Y�`z��VW�/��ߺ�|O�{����<�Z|=)�QS��y#���1���K��e>�����2l�˪���K���^��������������������Å��Җ���,"zE;T+��"�l��NH<2�<���x���x�B�d��cC��r/vbi@�)F�lL��Ж��I�tM�EC3��y��-U\!���t��+�����A`_�������H�&+�����bzNPa{���	��\������������8�[�o���w��8��K��Z�j��ـ����C0������㰲F������@1�J�{���X
N�~��� F�����{�b��a0���}���f����D���,�}t���O��fĨ�s��ӵz�y��f(g�0��x
!�#|WԸ������2�ݳ�G������������G�i`����ro���;Ж��v+�wj��N!���q�W�o^m��Ƭ�y��P���co����A/������{�q�i���n����u�� s��=����Ҳu=ˏ�
�ɗ���f�pp`�Ы���d���e�p��o-
.��y��y1�R�+�}x��<7�zF����/Z�4�&_V�����+|�h�>�c��2L%6s��#����{x_��a$5�d�F$?�ӣf<��5�-4^w�8�Z��C�bjr]cU�[Zf�/�ƯZ�8��h����G�+�-5�Ұ�=ABͳ�5W+�C����L0����������T�.f���hS`��k� ���~j�I�u�v�����H�;w�;����0�v��9���;���F\����[qH���������e>J�=�?F+���3<�a�!�m��!γ��`�G�1g��Ը���H�[�/�É<	;�^��q��-��*ҏ�e�۠�]�kA������������f��������aꂇ��������������������q���7��$��-���O�-F)�$6�'��I�Y��Hy�5��딅'��`[�]��EY�"춐,�)��+�kW����rh�E�Im�M3���d"�������7=Z�'d��@�=�Z�_^�}������{bQ�쫟�ß�����,8u��t�m�x�Q��7� ���]��7�Ē3�%�<�b�F�CR��;�����_8b��LExq1��J S�\�19T��T��� ��l93ǡ��<_y\�jvFB��>�^m���l	Ө�"L��X,���x-��=����=��?�Ѝ��&I=�͘vJf�C��o�w���|�亳1O���(�hQ�o2~��YL>ji�w�>2����m�g2��v���Q�Cń�^�� !3��M��+��[Y^��3�>0������gm_��}�yj/�d���sy��E�.�I��C��/K���?+��o��0ץ���{�^T�Q��D�0xa���Ô�oF߄Z�`��{*w�Q�0�sGb+��x��l����A댄���E���^��z�j��H�q�w �0)���<�������C��f_h������٠�>�`�3TA��&�Ymh��K쓧O�p���w�h�w;R&xϛ���ƍm���	�a!�U��Zk��a��y����kI��c~�rZB?K�=wRF�	2���`�s�f�Z�JӐ���T�6�w���rY���Z�Io���[�V�a���%�	�v��t=Dv��~��gjx�π��� �v�c~�0C#+]�z���<�����������������������'g�^g�M�R[,��k��tY^m�$>G��J�Z���������[ԝ�y�)��A��p_�&c���ċ����`�͡��<9���Sa|�╗ނZT
��Zb!*�����;cY�[ۍ�Lo�� Z#��2,2Z��Ж��	�T.���y�nҲv�-J��ҋ�̐"���O|Qxz��Ki�+���m�m�2��ә�QN�I���3�ѧ��^�@¸s�C`�JS6���͘��g���X͓`�������R.d8�{�� ���I1��j{Q��)� ���_o>������[T���ݺ� ��^f�Kkk~M������=jᱟ��;-d��~eI��;��89�5�f��-k�_-��Gf ���%3D��s��D��iqm\��c��OڶfVL}A�e:�ޟx���=�5,�c�g���s�{�L���?j$�K>Ʒ�τ�8=
�y�3!ѴE���g�{I���km���0��`r�F����|0�B�I�Om��ug��"���/�Z^���̨]Z�aMUJ��I~T����j���h�)mp��1wұ}�H�e��,Ԍ��P� L=��Uy���N�L�-a��,;�`����������0�v���i[v^�Ou�ê��YY������C�� #�-t=�b����:_��ތmMzSڷ|�aR������:��F]��&��v���'<�0 �{B:+��_o��}�+�H��d
v��W�m7�s/���ǜ3��w=O5_�b��z�w���9�=����}� Wg�ϱ�F�P�+��x�2PNOwV��lV�|xI��E��-�6���\œ�=;^�xlk_�'�z�=�r���K�^�7�����R�����S��I��0����'*��d@��Qߕ����̵��d��`�1�:�0l��t�틂[/�6	�!]�+`��t�7��N�nw��Һp!K�mV&]�8C
/�?ZpS��`5]k#��q9~�,(	��޼�\��o�#h���l.�Et	aU0���-��o��!�Z譯R��"�c0X5R^~#���T��;��h=F��5s}:s�py%͛���_0κ�#�BK����?�|�mH�wj�-�^k��H���a\�1���>���Z�1~��x=T鬬H���#���G.C�fx�l���)ƪf�D&SxAXT���ü���x0���L���/�9����&f'�.��(�.(�̳JUڗ�h��k���e4�#�>&h/F'��Q��O�a~�ޚ~�o��$v�a�f RC͔C�QO2��|�f��aڧ�ܫ�H���>���8L�_�>��{)$��ҿ�;M��]�H����?/뻇����J�z� ;*�&��&�1c YDX�c|V��*��x�~����P>�7Y�dı|��K}�y���,'���s��lb���&;I6�%\�f����Ul���\��
d���Kk�q8Ay���uU�^�8W���6��C+$��t�z�c^�������}�L3��Wg��������������������cn���s�0gYL������/iM�.����F�Z9v>\���ޝ�� f��#Z�͉L���]JZO3��kfK��ri���`�鵅i@&A��d�Ta�ܾy#o޹��nH���Xx�o��aJ���OD��̇FK��E��^�.
�����%,xE�o����mͰ̤"eR����w��=;/-�Y5u�vEz����	�]rE��`!][�f�X��|'Fs�!��օw=~g'GrߣG��2����͔Ϟ�a�,Ͽ�!�W2�f�f����ת�|�tK虑����|z�G�1y�5{]L�d�7]#rVP��Z��a` �N��7�;�ֺ�}��7A[�ՕU~ҏ����L���-��|h��4������L�u0f��7�Q�а΍3ֿ�C�ȅ��̻�8���ge�e2	y�#3���E!0��@l�t;_��#��T�=6�3� 4�"5!����=�f{o�A��e2~�Ԣ��@���l�\pշ����Hr^M'f�v@M�p��!��P��]���Y����G��EW�������Z���{�W�6��t�:2�J�MP�#h�q~��_v�d�6�</(�^`�1�d?�~�ە�����Џ��59�y~����x�P���0�����8���͆����KM?�G�lP�O��-��x|�YZ�E����SL�V�T3_��"����&h��υtMQ5H[y�4��~7��������������������q`��+��hP��4R�9��c.�'�ܑ��RȈ��G>dV�����+�	mZV��t��cb+�+�ɖ�eլ��+��Rg��)h�Hf��"��
�UXP��AbskS�/���f�ba)�����}��^�������©@�w�=�a05<%��g[`�Y�J�`���s���-�7������J���q�~�"8��L4l����#���Ev��T=0"�X�����Q��^p�w�zU>d�QU�����>)�q��O~,�9��w}r 20�&����L -���M�	�/��|����o���Ɠ����m�\�<�K�+�q0���<6ڼ[�Z���x�x����oݼe�G�>&�ED�9�d8h�>j�ѧ�� ��kiY�;<���)F��h��y3��2�^t�`^-���]P������K�*|)�:�w�}ל�@9�uQ��֝!��&'F��u��K�� }�����Qi{�^�����	�.V��䵵Kgż��Z�l'Yn�?V�&ڀ�u���/0ڊ,��Ǘ<.c�D�:�hV�/��]0��Аe>��#�n-u2�Z`�1]CT��d�/�$;����@�mO���	�%�u��qb����ǜGR�B����S�_ڂ�<�DiX�=���˘ב�ǝ=.ﺚQ���@��g
����t$�Ya�ui-rǼ2���d���|��w��������������������qpa}�V�鈦��/�H���^ �hʢ8�Om��NC��������:���7+��>/?bqE{ �+���f�j<�28���\N��b�bq!��MA2��P~_�F~G�>��ȴ(��4�%g�
�?j.����D���qzE��a9��+�^J����;�����*�t{��v�i��t�ioq�h�2�johY�f�3�M�E�b"j�LO�-�6�.��\��Se9WϷ�����G®2���o?���D4Tz����ʚX�_��kq8.H�<��#��`xmk��N`����F���|]���Y�w1���?��ڂpQ�_E��b�!����ϓ�G>˙�������uL������Y�/�Ь���:�L��2	�w�~����"���&��%}��{.�fN������^Ŕߓ������y�u֏�p��`�S��9�bG��~�Nz۞�m3�����������G~x�v�@/��/5ꐿ"�w�	��S������N&��I>���F���H���x;a�����=����g��HoЗq��Ɉ+�hn�]K��q��%wPmƒ���Ω���lCvD�y��8\[�q^�;���c?ׂ�[�o#h���J?GM�1�Qhӷ����cI-����=�P/Qߎ;����Xƙ�+2�쏤d��ҟ7��ߍ�M\/��&ӱ5�5��;|���Go���k>��Eh�p���B�e� ]�U�<���������������������<���\yT�)� Z�a9)N���FI�.�*�����9����D9�j>�Y-k��ìh絘)f�UǬL�,�M��h4�	��G��n��-/媭1�N��ț���JmX�_Z`N�Ds��2sZ��\�2�_�� :z9%���R��Ǚ�Y�O{-��UXj<��Jo���Q�R�{)FP�b9-��Z�h�Ӛ���N�	�`����扄Z3,pԓs��S���ư��Q��M�4�/E���dL���Ci�hɥ7�]0�h�o[i��#����3eQ��*=��Ǌ���1U]H���:��/eie��3���h�d���D2�H��G�=���\�k.�_��S�cjK�4r��c>]^u�<y��`�3_���1�wAf}�}Ыo�|R@'ma&�;����O����56�e yEp��vV�an�5W�H�fko�N���Ԍ���}�N�g�Փ���x��w�2������0��3��>3�&1�Z^d���j`����%SjI�1M�~No��Q����f���xM�Ⱥ����	i睹$^V��`�u�{�~��P�5}X��\n^�1g5�����C�w��<�C�#7n�Wۛ7$|��Q�)J�A�t�g=x�'#\�^����zկ���q��7�aj��4'J����h���o4�V��k0��R ��*v�t:��k6��G�>���t�L����iPT���\_*��\���C�wb���|����%<�������������������� s�Ok�Y��c"9�p��B� R,[#A3�c���{�5a�0d�yX���(fOb� cA]����g:�gH�ɽ��2ә7)KYEə�3s��f�&b}'sm��8<�-	��0c��Pti�i�����r���)=��؍���}j����Ew�0y�œ�&� v����ipq�33,,��bN�2HMPb;B���_���nI,J��������d�用�:TZ%3z��ןU#(R�<�;U�B��)K�y!�8��o��J-�@���S�bo�sʢn4zl2�I�|��̻_������ �Cz��TDSEՋ�#z��0 c�ǁ�9y�j�q���Ҽr^��:g�3+�}YL���P]YS�]�<]c������
��k��_2~*Za�+�jM��I�4��ś��qC�c��d�ݻ���ڲ���h���;��0��c�h�Y����Cx�g��u�9�,/����Aimq�_�w������sj1��[�¼g]dg��
s�g&�R������^ǅ��W�~�����c�{j<ȻC���<�'2�J*�l�k-�����`�eiкڳ�������������*�D�Ѩq�;��L+9�h��fr�	�F����a������G'үު���V_��D�+5�7C%+qg�䫁zpsG�+�O?Q�!���~ƒ��}0��]�\�p����V,���S�3@9�v|�f��7o��޽!�ӧ{ү>|"�D2�
��2�z��8�U�"��'mc�v`����95^�?���VͺD�;��kKzF�������������������5�Y�����G1��E�T�N}�]��$K�8��6���E{Ŵ/B�;�	�=�	3ɥL��������v��|����s'����|��fX���;�;>[�i�e]�Xςb���X���B��s���S^�4�/���T���_�)ā���`�����7T�5$��Vb�ٿ��_�c8��)o�����
r������DS����M�Y�Dg�/�	��S�pZ��/��rQ,��
3>�?ͤ5�e��`
������յ8<|�������`A-��e��ٯ`z�O�<kiY��1�����u}������|�(g���W�sY�x�b�Cږl�`#s�<K�Zΰ�~�&�� �AC3N�w���:f�̇�6<<b=9��c�d���#?9#�w�qN^S��q����5m�蚍��Y���u�B�����]���dLyEX���x,����ɶ�O���8~o�����=���y�̂��^��_j&����n��^���36��
E�5�+�����T}F����Ԛ�!��F�Oo�*��mhâ�77��:կv��|f�]x�jGb��u��yN��4��'���`Ws��K�c�j-������Fs̽1�xղ��ބ�^Z��蝌m���1��"�����8l4�8�T}����]<߱�|z'�����KЪ����Դ/f0:�	�s2���1�}� g^�sZ���Ma0Wo��Jz����cY�d%x�Z�ݶ�>���=����撬0�n��qs�1X�-�ɸ�W#�ؓ�B��*i��ȶ��VZ�3Z0�?T�]Py�,ND�d2f����g5Qi�`�*Z �wI�jN`aj�H���G��S��U��y��lg��bl)M.��m��\���X�T�|D������%\t�]J��Վ�Ȧ�	}8��O�h@#2���2�������_��N�+��ƖXx;�'V>��b�l�_i��j��ǅ�|��ϥea���Do��~o�44��.��4��қ~?����`��کY��9��S��A��K�=`�N2���z�x������8t���,�]0����֒f>N��3��=x#4ZP3j(���_�oQ^��|�ψ�y���'Z��u��9�QO2�f�4[}����lt}/�L���P[�Tz	s��{Ɵ�V�������yf��?B���i��d%Nqm&_�DƳ�_��f��.�_���9^���.,Xǉ�`�X�\���/V#���저�k�s� �_���j]B2�=9.����>��h���_2^j�ϗ^��G�ν�Z���-0¼p��^��ʭh�>FVh��`֝ =�C�������ļ�L��5Ikc3�ܾ�-�<[^�S���§���1�Ch˶��w,>ì�6��%[k��xu=th�R�����a����>�k�����.��k��� ���������:'`�����(�� �=0���ޖ�ݟxIV���]���O$����sKw_y)7o��ƶX��S3��7_[�����LB��|U-�W3�#�)���^�T�:ݩיu��gi�~�L��χv��u����Wc�t��f�ъ��ݓ㩷���&��O˚2ɥ4?i�Ԗ�ŀ^�B0�*�̍��1�#X�^��g���=�����t�$�7�v�shoJ�۞��\�J`-���D��ɣ����Z4s��p�wEH c�3�zS+�Q.��J��0T����%T�Ƕ%ҥ���W��:Y���ho��}��4��r�Ͱ��\7`�T��-���t1NT{���[,�K��p ?��h�,A�g	w�Mץ�7Q���^?W>赐�2!t|dR#p���T>�M����0����f�i��x<��騽��ʐ�����v^�Ŭ�F�>��7>_�6�q�xɰcF`� 
��L�y_ǭ�����e��Ձbͻ�̥�wV����Q�F�`�qǂ��+�����aa����}��E/��>Ѐ7]j�9Ϡ.�۝m١��Sc���qx|f4 �k�rH��Ԇ��_�l��Q-A;�����W�/s\Z�B����=a�.S^��r;)QO�a�/�-��F��o�y�Ǐ�s��8���	����N{���c��8&�����PN���j���*�W�i�?�6t:e+~�`xF�������������������5��5��-�+�Ը���DVz;'b��C�������~�����=��ߑ���W��7~�/����N޺){���F�p(�~�[��a�-+���H���#���#~��-	?��%�:,�E���J�8���z�V��R���Mv���+-uA�*�����j���m3������O&ʋ*�0&���*"����]��n���~�/��!�1�5jQ���6C�TsZ���al��2]�aQ�E��1-�#0%�@���
�Õ%ќ���wx��Lo�;���x��~ߢ��;������4b��})-��ᢘ}��C���=tv�;Z^Y��Q}&&�6s�L���₈[*���ߕ#�(gzE;|�k�?{9��\]T�f_��,��|�b2d2�&*�jCh���F"��e̅9�T��,��%���;�5p��F��hYy	~Q��.
��7�y7���ua���@31�ys�h�ύ�E����@���; c���\��A|g&Û���ܣ֘��*��)�v���S�5�6��w{�/�~�E��z��ě;WF����Rڈ`������u��u�V{�u�%h��؏B3�>̎IzgF��������A>�}j?'ߏ�f�X�Y�8��u�vl��WF��wjI��C̓�����\'Y���w_��7>�FnB۷/�̳C����o����AI���WaX��Kk�%Z|�6�i�fޙt���f}x�
�z��}� [��}D�,�՗�މX������}��qx�/{�'#0eF��_�����?��q��,�z\�n6`Q���Gq����r��qw �BI��#���~"�£=0�b��qW��V�e��V?z�I:ʲ�^n�Y��gq�p�1�&Ĝ�gr���ɨH{�o�ٛ\&����ia��kb��\ɶ�!�	-��\���\�¨��}���B�l�{'4����rE&`:?ә��WXj/hM;)KI\�1KK�U�_���+|��Z
`9��jX�zؖ\�|�1&�t�n�gL3�3�u���ꇔvj�B��e�d1�N?6^<�� ������ُ�e9Ҕ�0��"[e{�?��Q3O�K��eaV�a;��0Mg&�Mg$9��h^揋yjk�\����oЗq
ۇ�Uy��hBS��ў�`ϙ1u�3�zZ;��#C@�����ә�l�Fci/��	��n{����5��e1���x�~ёx�u����sR�\�w��|���7�kd���x<*̃�V�����C��ە��u0��B4}���'c0��R	��5o��J���;�FعX�z%���oa�W�z� ��O�-g�Jۏ�4z��@����\ULd�AR������x��p��?��܏�R�p�U0�^�d8�x5h��a��˯��/|�qH&_��	RSrzp L�rMʡ���������M��ǝ���_�v�Y~j�)f����b~����1�O�Ou�Ra��W�Q�3�<<<<<<<<<<<<<<<<<<�2��&^v���Y�}����᏿�f���?��AWV��}	��_��q���w�׿�q��)�u[%j��y�G�0�
�?��8|�t繫��H,޽���-�C�G�%ߑ�=|(L�O}��qx�x���d%��=�3-�6��p0i�wU�p�W����#08L+FV��ڟ������+�����D��e�7�9���"2RS�=�h�MB$�P��Z�d�m�+�'z��؂��az��^HӚ}�E��0��YL\��h�9E�4�BI��.����~F�Ti:���[-g��48�>7#J}�*�e��P^���3u�(/��D)�k0�:�9���ҊS�%36`*ڱ1DB�q$��FA�]�ǔs-�O2�s0�m�NS.��2�O�n�1-�+k�i���C�E1�F��0��Hŀ�������o��˰�/��ӭ�����)		2��� �ax����+`�=0S�m�7�B�x�`�RK��[�3��o�2mTo����u5�)��ypN��Y����z��Z.fG������S���^2�Q�w���-��/�^$��b߷���jS.��Z����q+wXL�/�΅�d8���Ԉc�/�� �{����D�&�ɉ0��6�@�Ƿ�+,fC2�q}�.���yʪ��knT���]����.�|wnߎCz��c�14��`���f��2?�}K#�2��K�3�g����ǃ�*�a�IX'����50��d�AD��7+�~�g�yxxxxxxxxxxxxxxxxx\̼��2y�ҝ6��'����G�ޟ��������8�Ud�zmE�z��������a{�Cl�.!܋�>V�����������|K�N�d�wͱ�HVh{`�,U�Kfs[,�k�Q_,�o��I�+��[����"h���W	\�w]0[��'ȴiM�Y��/��:];aV����!�QD!��#0�&H��hA�1�Иv�Ӊ7N�Y����D6�'�Ȑ��Dy�m�wGF-)���6�;5Y�@i�i&߹k2��!�F��z�X��]ڥ�W�����<3�UrT�>h�����E��S�̼>�H����{��w2C2TJ��h�g�[�f�r|>GV8�w��^2� �r�w30��&�91>	p�x�����[���ŲҸ1�O�c�a��
��}LM4j�̩u��3Y��`,��ݘ���DQFG���Ok���>ݾ�9�|\L�`�W���c^X�h/��o�V+�A��M��,�� d���t���l�2�?k�]��J=����./��4��c���>�6��`��]{����ç�Gf��^�ކM�����>����J1���dzt���Ҕ�`���4;��C�,�c�q���pz��;�;�|��y�5|��FJ��h��ߋ��f��x�M���3����λF�W��0�|�BͿR��|6�j���V.�u��ɺ���gq���|iaG������O�d�d3������(丶�q��	z�΄	�9�x�%�~�|��#��T��0���3�xKvX.QK�^w���U�R��w1;:_C�|yF�������������������5@9�	���b0�)�hв�J0�X����?��h�}�ߋÇ��]�"��}�sq��/|9�ܾ�0����8�uSV���DKo��0���a5����+���|J~Z����w���jU�[���FX)��h�2o��{"+�O�K����]�s~��Z�����"�S�\�l,)�+\�
x>�b,�-*[�*k�8�b;�� ���Zg:!]���Ѧ�a���dD�R���N�睆�f_�R��ͅ��͙���'`Ҡ^w���[�7�ݧ�s�[��u�9����r�,|&7%z[
y���,�A�[��b�
�	b�(K�j盰��k�����yQ�����b���2_"��}omZC��E�Ă�"�ܓpkS�����"�'&� v�Q��W���)v�W��a�+�-����K�m�dR%���ݼ^w��F���U�G:錸��|&��y��-�5��㺏��R��u��d�Ό32�>|����ɩ�ߺ)���߿�%Ì��O��rboo�
5��{R���y��9:�~h^��5/����]}�33�.X31z�5��3e������d���`���f�%���l�P����OL8�F�fc��0n���a�����く��n慻�N/�(U����;<o�%�0j��#���!� ������bG��Cy�1^0^�qY��p>8��1�G��I���-8��5��ͧ]Z����o��o�;2^�u�σ!2�ǒnw��s�����lA��7S. ����c��p��-;��W������-�?��"so/��n �oo?K�����߷ޓ������<w_�-e0�jMh"6%˫R~k2?��z�uW���6j�ՠ=���&���C�r{�Ÿ�;Pp뙋���n��aevl���}�e�2n�N+F�Z�7{�#+���9��<��w���qH/�����8\in��/��/��?��qx���qx�����D������`Ř�.�X�e%��c��ѐ��7���
�Q��̾���8�8�Ƀ펅�#+˫�b)?�����#��&�Ҫ�O�.+�\!�
&uK!a��3*�(�_�uNUN�/_�f�S,��F���f��b7��N�}�aR,�������z���k���������>wn�%�����ڿ����b�8�U��������M�A_��a��~pd��*��Kko0Ƌ.��H�(˶�T�-�4�$����B�&��.Iґ�t�GvFpiI�4��&�b��&�{�9Ny�:���̮��ʯa+�x���f���sV|zO��2D?U*��R���K6M�`�2:����j+FgR��t��#X^#坮��s3�\L8�>�N������|�����ml�v��,�l�jg��+/�C�*;���s2�.�-15���C�B��!�£#x�=�{˄ь>�s����)�E�Ɯ�~�g�]�8Zp��t�f�G�(m���)����~9�TF��`�WF�Y���N�1���U�/�_ͼ��z�&Q8]Kuq����*G����AƔ�)f�ѺU^g���y�"��/�%5�@y�x�\��� � Ԝ�Nj���-v��1�i`݃9���-�/8>��gg]�O��;�ߩxX���ף���WAu���WB�&����_����,C+�V��F�J�"�!8�&oʹ����]0�Q_����ￋ�J9`Z֛��ʆ0�V�%l-K����Z�\�)c�L�,�SC��}���(T=T��2v�遴�Ԩء�n���{�>�k �Зh)�LA�N-�ˉ�Ca��"��?�V��[ߗߟʊ�RC�x?�����W��U�����1��l�
m�4��X,>�'.�6��E2V��+�''���s�7-ޛ��sO��G⽅{����ֲ��ٗ��Y��Z�e�{o~���!Z4�<n��$��qH�ټ�>�6p��.�`/�<ak#�J��+�.��D��t�O'VXr��gh��iz�	�]@�@z:3�����0�5�}��Bh�T�l|:�MnBk�Rѩ�xY:�vg*:,�����*�h����ٮ0��5hT��ȗ���Ŗ�(���]��E��@��K���c���2��`�߇��cU��h��
s3mR���b���|Ȑ�	u>�2��u�������^��REuRe�]ZNa�7�/��HX8Ih��붥_@�s$L�,�{v��;y+�ŀ�+����F��?��e3�sb����QP�e{;��#�&���S;�&&5�0��駙MX�9��}��X9:��h@ٌ��N5�#�-��~䬚�/
�hQX���P��׼�Ӯ����?k��}7��gf^�w����)��Տ���ݼϦ�'��B{oMiu�A�N�q������L0�]�y��r<��q��&���@4��������ʡ���X�󥙉���Eu�f�% ���y���L�-��	����4�u�/�PkQ�coW�wc�G����q����G�1�g�^U��O�$;%��w�C���ٲ�Ӈ& �m�1w��s-/SnL|2'#�(�<�ĝ-�೙q�G�M�w��{x"���;?���?����qBkE��vܐz�
f_sIʿR�&���чy<���*|-`'L���q:wz��zq}�|�lG��E�D�Є�E1��9�}� f�/P���¶�����㑬L>�X��}��8<x
�'h|{���s�������w�V|���Hobo��q/z+�K�����ë��X"lM�:�l�U�ɓ'q�c�V#S�a���;�K咬�7"Y��\�5��]X�I��s��B~ؖ����
�E�x%�W����Zނ�t�U��QO��&rX�x�)Ƨ5Y�IZz�u͈u�
)˔�|�N3���P[�l��J͘Q�#�,�V5��a��t�e��'嵹)��Ԙ�F�`$���Xʗey-��+�j׌�^`���|��R�������Q�K̘bE��Gx@�dI�;�ی�$�L���r\��Ĩ7��7�Qna�� �w�1u����`����I�)(�H>#"�/wQ�В=�&	�i �Di<��IG�e�Џ�bK�jd��I�o.�Ev�h��3-�:�{r?�kk��^V�ev��X�c�b�AU�h����q�b�+��6���s1�X����ֱ��D������������d�9㟯�t��M�����.�}e�	JW��my,��c�jԇ,D�˩0�b���}J[p���2w�B�Pgs�$yMr�����x��]���;sCp�y�-W�Z�zGF��󓱭�7�8O]q~^�������ʫ14^|�3��	�b�qQ1�&Eh���#Sl"�\�riI�g��"��B-��R���n{�i�|.j������q��.[���q�G��I��ֻ\�t�d�a���0�d��&���a�l�}�4�"�{q��)Y��F�Pҩ#�L���~��Gq����/Fr}����&�x+��&~K�_Mi�Q{�L�&����0�8����}T�� KlFҞ@D�Ҋ,L����������������������F9�3�S.M��(+�\�}�D,�o�)^u���.��6W���eh�m��%;a�+��{��&+�d��W���j�R��_�j����#h
���K��E�0���O�9G���W�r����R������t����_�%����Z��J4�Vߋc ;'���WPϴe�P�pLm���ְp1[A�S1����m"_A1�1o���X��ʼ� ��&2��]�>-=2q[`�T������!���yMt���x����/��P�;��#h���H{VCj��A���̦&�:r���,�!�f\�DI�h� .˳N悎���[P��p�z�H��o�����Z�:�l��.����Z��]��O�5�VN���wN�Q�������dW���<��}�zcͥ�J*	�!@B �f
�lC�il��n"L8�a�nG8�� l�6v;n����n�	���)�B�jz��7�w�{�!M�����W�}3�p��ߏ�n��ܹs��̝k}�[жl5�0#s Hu�<3J�M�Z�	��h�S��)��@_}1��j�t�4����Z�(K��:�k�/q?jrFC��{� ��"�N�H3��h���Q30O;�o\&�I��q�?��nz��ў��k5u�I��#�kZ6�~*-\�M���v\Q��D����}hT����Qfi/�����j./�)��/�2��Y����������~Sˁ��N~?��y����6P�N�nGΰ��$++��&\�΀~�%�%\��P�d�y�dK���y|2�Vׄ�GF �;�<��ӱ}����x�띒+�����������
��g>�Ǳ]Y�q��׭�\� }���̂�����g����'v�
4��/��0�dYxѾ�_m^�_�"��9�FX\�v��!��`�UKr�s��P�qR1�5��f,��A�lb��s(c�>-<���������������������FG�\�q�0���k�^�헿�e�}S�oK��i���|}l��>� s�ģ�qW����*ZW�,1�
��{�z����B=0 ��y�x]�9�g��EѮy�a������ʺK�5��h���M�<�{C)i]"蕲x��RN}�Ά��0�>��&�?�t���])/�ifP:�r�#��:Җ	��"�FF�<�=�9���P�����'a��dt�S7t�X���t��D`���9�cmaՎ|�Ȉ�9E��kh=��ߒ�Xϓ:�LQϠ�~TG�;k&pZ�=��C-�bǒҬ�v�ъP,@3�4L�g��.�ݤ���cf��[O�v���Ȥ�2�o�^���>��w����@��=d/eV�""��#�9#�}h���J�Ed�o��vUD6�]dYS��cf��f*�,���ݖ�9�z)��{���6��-�{�;��_�Cy�R�}K�q5���c�9#�Z>��)�Qp⌧�=��|��=3�����!vZ4�ⴎÏ�)��r^8Qdet?���F�zO���p�s��D3��10�0^+�{��j�7�M��s��zSk���6�Ӄ���W_���fƹZ�NS����;*ŀ��ٝ�4�r�N-��Z���u�`��Ҕ��R�O��e�������rz��e��eW��.�g�eh<S��BC����LJ��t����g���h���������(��h���h�e|mF"Ǒ	��ޮ�qg�qsS�I�`�ݾ���_{�<_����%9��W�/]�����:���W)J;2�n�"�1��04M���>}�c�^�j��5-<���������������������t�O����@omID��^������a}�ɧb{���7���n7�s�A��NK"�{��{s��)5Z�3,��G�}d���5�b���������>pY<�Md��tȠ�=�}�Y�'Ydp�}��DJ��I��6<�Ձ�]��P�)����d�uVJ�7j�1rA-�MG�hL)m5�%ց$�f{�vC���bq4��ً��4"�����,�"F�� �a֠6�!�*�I���\��H٬��*�����v�:ho�>��߳v�]��vg(����U^�"�\����P�&N�~C�ް%v��dwB���{��b[)HD���PX��8s�w4z���4��9��_|E��}TE֩+O
c��,SŒ��Ƭ�s�|�>�q�y�~?*d>?�2�"p�~���㼁����~1�=0�/H$���y"�M0����h�Q+R�c�6�٨��~�Zl�C���~��&Z-mD�'�u��htB/��h���P.�|Y��{�1�&�`8ZÆ�ˀ��q2F��3�A�9d�-��P��;y��IC��z�L�Ya\ɪ�>�̾#��	i�M����K�������T#��L�DN�{�R�u��P��|857�����Ǫ,�|�3�)�aY��3L?0Ţ �G�2�H��;0�Q�9|���=���l�j
΄���ɱ}ֲ��d��f ��#{���Ǭ?ߗ�
�t`���k��NƷ�~l� ˾���І��Ō,��++����3��iU+6�/����^�vU�p޽>fRW���+����{wc{�ua�U��>����3�s���t�3�}�r��}������͗b�����ʺ�׍G��t񲌗/]Y�yI���f����\���rj����4�u��p!�`�_(��tL5�/Gn��b�{F�������������������9@��OG��d6�-̡~�yxZ��{�Qa����եZ�� ̘<���#���d�J�Ypk����&����fa��#��Ud�}�c;�/���^m�V��<��Z}���,���Ss�s��&�+]a6�PUh�I�%d�-��|�`J��l��8"�"X�j����.b���°<�F� �������%h�-�Hrn=\9�I�h��'QS��tj��M+���$�9���<�>ojEj4��Yg��Z�5���C �07/�����o|F41+�o����V=�"X�Ϊ���T+�������^y�yk�0p��ȽpM�d�-�u+CSΥEg�/)�}XA֩��e�x��_Aw��D�Ů��n;�})m��U�>.����[\��N�.�[Fy?�����rNř�=���b*&Yzy��{b��D���=�v�Ni�b=�Y���V�}��*�6���A��ݔ��zEd�.c�ו��64rY���ko�~�χ*B���\��b�����fv"�;������]>ۡ�:�2��m���}2�x_Q�poW����fn��p����h������AmA�d Sąi�I�vz�.��4��Mx�I}Z5�4�,L����aX��t8��l�!c67ߏ���'�-���K�|E�VpF\�h��H���z�����H���{	�
3o�R��س����</���р�:��9�̏�^�*F�^�3~3�/�>N�
�q��n��Laj��;��f8V�2�X����|sFC�)�� ΍�1��+�~O�_�zY��v�x�ͺ ��%���}g�lK9�?���v���2�M��f_���a��V��8�p�~�'��~�ӱ���>ۻwe|Y�������>�hl����*�ԡ�W�q���v���BjcFf
��-�{��R���߸ީ�˼=4C�t�|3�����N��}� �8�FS�����F��_FNss��T{�[��źxL��A����l#+��N�L���f��ݑ��ʃ���3]A�:�����?�0��goF��Pd����r�
�0V���9�s�A^Gv2�h���V.� G/=̌PF����G�$��ѕ^�"=����
�:����<�/��h<�!���ع��50,�E�H��<�H�2�����k��/��B	�釥
�b=hte;F��@���v��.��m��W�4'C�o�6��f�����~��ۋ�jG�Ϟ{���>��?{�a��h)&S�DX~��?�W^Fp�"d͆�2�U6��-ݮ*tb�S'Y?MC^����Z����2Y��0HY[k%9���}|��e�͕'�l̭4�EM35C0sj���Ͷ�#��g)�m�~����2���ػ���[�*���wb;������ϛ�٠m�;c7	n#2���/[���x�i�X�[EV��~���0 LVA͔�#ĉ��҆q\?���:��|�0ka4[���ϑ|�fVڑ��4\Y��.�Ү���iL��p �T�zU�odp�>na*��6~6���cR��<{�"��h�o��[�s���-&ͺ�*v�R���������7�P�����]��� dvaү]���`���e�/�K-ہ��J��9Ӏ��z�4�
!�s�MvY�#�-����{��qf'�ġ��@��m&�K{��Z37H�pF�����lg^�}�L����c=����҇�H�>0���2�[�]@���;��T)��k1��__ΏY��c�Qק��������G�KԔ+X���B+piQ���D�+�>�׹��keYơ��7�����(��6�M9k�eܴ�%�������~����k�ޔv(�~�H�������$_X��2�{p����9��<��u��=��}���{�&l��5���xDi�2�#��c�3�<<<<<<<<<<<<<<<<<<�2���;�H�Ζh�mn�����xZ�Vģ[A6�zE<���lg�T`PU*���J�@L���zO,�_#� ���ar��0dd{}�Rl7�&�L*2��)�"���z�s�c�'��덆Q�a�p 0#j�v�͈��ќ�J�,��6���{��l��9�u���d�aV��f����fP�_aN����\�Kׅ�Q[�~I����W+��P�oZ�� �rf.>�_�,��F"دs �X���Ǥ�x���а$^��rl?��ۿ�뿔rp�����9���ذ#Q`k�-D�^�뿊�
������5#3*H��ȉa�9"vZÄ}�x�j Ӑ�E��k�D&�K:��rs�.ض�!y�ڌ���P��*��b����G��7�C[�#��Ӏ�Ը�����0B��vK"��+�����Z6Y��>v��k�y�D���׭���N]�:���bohW �����B�3BQi��_�s��:Fn;ߴ�y�z���s�02��\�ge���F�>�w�x4�^�Vcp�@�Y�騈lg�!�fg���O�U��������M=�`�oޕ�O2��f�U�����MMj��(	Zs���0�'��h�j������8%<�	���82��&�ۼ��d2��*����f�ٿ��4��z�ۓ�i��x�Gܟ�O3C�į�׍���{���0ꗪd�a\������\���檨��kkSv�7�;�ƃ�V��X�	0M�bwOftnmI��^����Z�J��T�?��G}�o
��?�q�?��_}�˲{UN�����}��7d��rAڭT���gd���0�|E�d3��-��t���ߩ�-}=�C���.H��vK�|��0�4��������������������8x���z[ӆOf�ۃV�ì��gwy�h`��ӂV��B2�J�q�Qn�ۨ�W�c�����lm�fS�/Q; �Okua��,xa8��o<����q\����ē/ۓ��? ӱ+����p����QT8����#����E���dוvo5��ߓH��d}d�Aq:[##ge��]yX��F�0NM?CD*4���&A�A��f+�'�aQ����2�B�(Z��¤�yM"}��m�5�����vY���ǟ}��c��/~!��y����B3���틈��4wy��DHi]�w��a���,�*�0m��y�vl�D+��K�b4ZsvD/	��qE��F�֦.��d2Z���G�h��E�9��BED��m�Jwd)�1�̂6z}�#�9�P��j����T��b�ꈱʲ�l_d��~0q{�LT#��eJ�=򶯉�ⲭ���W��i�̬֜�a:+f�#o�:K��Ǜ������o�.�'F�9�p���0��&�[N_Jk38c�����*3&���F�Ok�/��?c����8���ٛ����;�H�'d�ȉF��!_�zm�hW����9>���7���.��r���Qd�/�v�?��Ilj�) dd�\0�-@���/��fK�wCΌN�~њ}z\�ј7�V�w]|�6�@2Ī�!�f�q| ��
r}�:��6�H��1���;���A/��ȡ|���9 �o2�6�	Sp3-/=pgv��0~~>����w��k2nx�qg���R2Y��?B��&�0��)���?����D�|/���ʫ����L��݈����j���#E�T�x�
�i����l?o���f���X��9�xݡ���o��皉�E�8�u�̹X��zF�������������������9@)����r����نb.�cj�[
mD����f�!���i��/̦�(�h�� @�m��0��P4���_�:w��\�rA����ʵ��_XO�Ғx���'s���}��.���c���lv<�<��苐�u(�%���0��1�>��ۺ/�jIi�yh7�_���a(̴."ɜw2Bʰ��K���(!kk�d��LDl��
fj��G�# Ȓ�~����`t��0a��u����7��-W�R7d�+�KD�3&��}������"����`�6��YС�,hi2t�����v�e�y�l�a)��3���q~&���Ugd���p\��"<���t����ܥ�<�lk��)��,#�hNDC�V=�:\L1�(��s/�~i��g�U���He����I~��p�5���m��4����Pi�{�7��{���
�l|�czOjF�z%��mY��1ޘ3Y��ζD�ww�����ګ�
Ӯ�Hd}iI"�Ԫɛ�����B^&t�7��z��r�;c��|�f���<��#̸�~?���N S.Ĕ�̭����N�}{�qD-�d8��ɗC���1S�l�}��G�:3uJ���Ec�֭[��{\kN�sU3�8>�Ơn�d�<-)�0@�hO2�Z�+C̸Q�	0f�n��G��\��������ڒaؕv1�p�!߇;[�ɷ�+�R�zT�b�]&��"��h�/��wv���w�ξ�S6�e&�5S� �u3�C?�[;���7���o~�7c��Ma�5zҞ<(٦�=.���Ŀt���W�̯j3������5���\P�%J}�qA��������ȅC��9��3)�1SK�gS���as�V��������������������q���GM!f�k �)�j��^�(YQBD4z`>5Z����x�k�:��X�2�a�ZS��_�f1߸���!��}�&WG�j�Q�fZDC�5ۊ��sN7#�}�_�"��|d�sO��u�҇p�2�a�܍K�:[�L�/��{�Nl��}s[��%h��6P��| ��e�1���Dp��jU���kXF��"�]d�"0S�fJ��{C�ɁtdGgc��o���>�,�����h|ⓟ��A_��a�2bV����v�V�11m�b�,
26SL7�$2�%1�@3y�~��D��3T&�ߴ���
g��b����8�9	R��}��G�aw�8.�ǄL�L�a�
4c0�42[����a�&����u�9K�]���<�
��h��>SYݴ�-AM2��w�{9PL�T�� �̶�5��1~����A���FGAv��hf������P�����baq��&2��Gͧη�lZ穙�.*�7\��b0zF��Ĺ�,���L��y��8���!_(���m|?����g�z mk3k�@gm�p�w�M�7���:�{b���}���4��D����ަ����>�w��4��������vd6`�!�5JF{�o���\4�8�A_�{�}y_�9���L��=�wW���J2^�xI��=3ުX�3�x'��<5��݂����컿#�o����l��Pʛ��gkK�����Tl����ɺ[^�q��~�=���0��>,�ċ`�qj\3(��'�:�J�8��LR\�莙0�0�+К|�����/�����q�`�ixF�������������������9@)���LOe�+f:F+`@]X���0���*�	#�X���x��E����1ehᐙ���r����.�1BOO}����߸~���0+/5��9o��e#��/��{�<�0�^�."�L3�i$��u�!8g�>�Ԩ #0_��c��w�+�ϼ���2���0��P��dHFZCJE$�%��E��P��٣�ݧZ�w�,S��>�D�
��"�Y�2����~6����������~�}l���nl�5$"��;����>�4��;Rd"T��t92I+���9ܧ$�5���)Bg�q�o�K-�Yo�H&��)����cI������X�{�rn7.#�m���7k�V'`��ҹ`��m.���tj���bp%�>>ӏL�$[0���yI��į�	�Ԯ����p���p��2>`F@a�~؁0��-.ښ�.H$�<��v�6k�p����!���w�5h�]����;�g�?��qgH̸�c�߆ �%���&���a���cu�\S/��Y�}qF���v�&�<�;��ֆ5ۙ�[�:yϐQt8�/��3������e�B�����E�0�Ȁ��x-�s�wHO�޷Z�O}7$�ɜY��}�Wh-�1���������i0h����ш��)�݋臐z�Q�/����(�7�"�7~�Uz��3��K��}C��>��A���[��������@�x�����Kk2N�v]�+���jloߑ�_y���އ��cO?ۯ�Z��_�JlVeVEV����_�㪈3��n��|��c\n��Y�.�a����HƠ��3���1�?��3�sK�&��������������������qPJy��k�]N�
� 0�3y'��a*+ �R�#�[��3�v(��~��7�J�V�D�f�-r���`W������8����#���Ng������z�ӎzQۭ�3=��t1G���\ �L1R8j*��@�#�}ZD�/K��� ��~��-�lQ4�� (�ֶ`䊑2O��w��c-�z4����]XB9C��a`,��6&�SLD�>�����H{O?�dl��u�p|衇c�cG�����`l���/������ے�Ld�nt�*�Z(��i#rIDKΗY<*�[�)gF�AZ�Om���L�$�J���@v3$�*Ҙ:����Ƭ��}<v�)��Of�=��Y��CM�uj��rt��<w
�1��X���&I/#��/P4M?4�?�[P�gX2
��0�9�񃊠S�.������}�l����S�0CD�w:[(�q�e��j���q̀��#����2c�3X>�{��WFd�LA2 5Ï�f���}h�0�����8���Gg3vec<�����f��!�efu�|�t��ӧ&�=���~���T9����톚9D�!���~?����PY۳4��
s�?p����N3�Ȏ�(�W�=V�����Hv�Ú��V�Fݢ|�����#����uh��d�Q�F�+�d$��mnJ�2 ��c���xbkG4����&�m0��1s�����/�ܓ���\���7��2�r|�T�Ì� ���W�f��&����s�g�|��� EX��L��LY��f����>P�zF�������������������9��>�J����ЪׅQ�=�i栘FS<���%� ͻ�u��6��7�,�����/��>�Xl���BlC��O,#������o5[�.��ل���n�vEU�
�{ǜ�n�'�lGD4L���f�\�(L˽}�T�%G�;hJd$����D��2b�6���t;�t���h�1�nf"���}�Zժ7Fv$�Y�R�@Y�h��"��VB��/���^�z!�4'���7���_�^�oGl����#��������)���1pDB�y&L5�0qw�R�Υ��`��b�:�$�$��_;�{B鲶�Y�t�ʴ{4���0�;�����ѸN�=N�3MLi���9e�����ݕV�~��0I��P�L���ˆ�B=p�h�$5X��ځ|�w�C��7i����;��K�}2� ?4Y�l_�%������ӵ�����-����ʊ���^elW9����r�J;�.�o"�u�pE�����u�(�s'o��:Kl�s���N�ޏ�<���w���u\ݎ�?~����L2̠Ƙ�&W3�m�Ȳ<!�(�`f��e�Hr=�X�+��ѵ���K�k�=!܌s�w����njƁz>�:�eG$'x���Af߂�I�d3�4P3�-_��Y������/�:f>e�a&s1�����\x`M����[2S�3'm���m�0�g.́���;e���)��U��|C�}��2���1s���d��������U�=5x��o��S��W�Y�O��ǌ�B����⸟�Y3�2�����"��������������������8H9�4��{2��"���#��>�=�ٯ�ģl�R�E�zq�	�Yw#%>��(L��a0P�!"����x�p/���J�{}�N�2&�ހfX�-֧F#edi5�ť%k}IkrQ�Z=�nD��(����@H�%?Ȋ��"K��}d0�!f@ͽb���&����װ?�|+82�-DVeH���Md+2o0򘭷dk"%L,0*п�M��N�� cp��i{YK`l-��n�Z�"����ݚ{�D��������_��SOJ��mO�}�k����?��������u�ze�0u !�8��#7Y?u:����
9�w�c�W�.I�5:BI��Pg�2��v�g�v��Y�3u[d"2�1,��d=��}�e1Af��7C�/u�c�߳v�H����2z�Ii�M��F;P3�M:��}�ezt�S�5��+#�����b�z�ڄ&L�4��2����p��]�B�K�����L=j�����,���7�Y���R�bD�Y"[`�q��dL9��K#4��V�O
�q&���煫��9����/{9��\�{ݣ���4�z�2�g�|8��S�Aw�`�a0��5��8Ci�'TZ�L��$����z��q��Zs2���r0�z���&��(d;��������߬6�d���԰��sj�6�웷74�}���PߢC����R�����!v�d\1�؏QcX���0crI�#h;��~�@4���Eïݕ�`�1K�ի����zl/\�K̾�E����R�L:�`0��Zc��a����`����g2gCs}��ŗB;����ifV��kL�\d����|?�8ƻd,zF�������������������9@��z�S����ٞ�Q8�-��l<��~Ѓ-�յU�޼yS�We��*f�e����h�@k��6;��m��_��o�,��d�����^�z�Z�hQ����ic}�֜�~FCS�\�Bs��p�4=.ӄ��ʲtrd~0�ioY�vQ��G��̣{`�U������#�SP?�^��gĄ�`dv{v�``B:���Xc�2U�7�?���?�Gz<��>,�#`��lH6����������c{��K���^ c�)i�b�e1���41�X_N&ݑE�3�N����4Ʊ���X3n\Y��բ�y�I��^�q9�y1�ّ������H���)u	cU����m7��Է5߇�û�#v�^f4p;���L���LYX�\��f���>LN��u�og�s1��eHfyg�ܹ�D�&9�%2���q�.��3�!��"�ј�a�����'�>_�j�1�v�7;N��C/�L�7���dt�}3��p)�EM=���b@kfj�^1��d�%3��D�a3�b���Zt}?�D�����\�&�Q6�\�!�ߧ�5043VBk{�ϩ�)��W�'��Yy�L�����~����(�B��HM�
����=���a�[�/��H�+�h�#��߫h��2��d�5(����^}Q΃�Z]�9�⏹pI�ߗWd�gZphY1��uI}`�~Y���R�q�0[r���i���O ��f�e}/��ӅÑ}��yE�)�;�ꥫ��\�}� iG��qI������ăK&���Ѯ/A��-�w{2G����V���w�duA�s�(_"����z�dq�ݑ8 �����:�<h��T6��r8���Ȼ�;��im�d�>Z�D����;*���J� �C��,���Y.�S��&=�`8޹{;�W���ud3:��0�
�:��X4Y��;G",�Jj��ؒ�#)�'��A�eh�u�R�O��?��{����2�.5��kUa�E��Nϼ������+��Գ���NC���GV�1 1�o�
\Ӆ��ϸN�
h&�x�i���]���!���0K�o��W�!��?R�Ù�b�ȩ���Ǫ
ܛ��E	WYy9N��̀mB����|�Yi%B])����߀VߴF����%DP8>s���{hfW�E��'c��cc�5#lV�9����ߞ��I3���љwf�KKRk��_��?]������|�	 6�(�x�g�GtԷ��g�UϙA��m6�k0 C�~ ~w����hG��=B�.�����xS���'�h�37B��@�lm?s��T�#���vz������B����6|3�zEe��A�����rW���|�lQ��������Ci�3�R�v�?�,�f����?�Q��'�1f&�;�f!4���}�٩%�S�����:z<)�ar��U�$[�}d��������������������8(T�>j��0#ל��5v�+Ƕ�(��ۑl��������v�n�[3g�gg]� Y[�M���#⽴*�W9w�s��/��yY�}��o{[l���O<�ȂCq�.����^�U�BY�2����^ �,T!�Kؑ]ƽ��	F׫c�>�i?D,x������s�t{�8j�=�O��t��t�<�H�d�(F'%R��Z� � �?��~F���?�{��u�fl7v$�Q�ͣ�������7��G�߉�7����?����؟Y{R��#�`��:�߇��ñ=@6����h4QRe���w�0���f��,�g��sV���L�YgŊ�V?Ni�8^��>?�yJ͚@i�=pM����<�֙MVp�^{5�Em�{!	�ڶ��D�V.���⹼�$�fI�5���V�G����������u��l>���9{s"�ʚG��uf?V���T�9��?j�����pZ�y�iO���ǟ4s�u_M��s1�rk֙������]^�D|�����L�t��\M�W�,�	�3���2YI��y��7T��R���V�P�tH�
q�F4��7h��ё�g$�������d�&!�9C�3&�{g ~�~@M�.�f�оP�2�!o ���CB!g�q���%{&�������k}*�������`h�����h�v��E�J�E�Ej	�Gw���ts�<9�����GΘ���M�P�3�<<<<<<<<<<<<<<<<<<���/+�ȹ��N���D�����{��0�n�y=��|�kqxH� �����9h���N�t�RA���������E��~Q}>�Pl�~7���/�qY�zȂs�0/_���lׅV��'��J�,�� kK�m��0W�$�p`���6i�E3����kt�����{�Ǉ��m"(���T�U��lW�Z*&��dY1SYs����d�B��H �A�b��09~���Il��6c���/b��ډm}LP2@���ے���=���3�����7c�!d���7	��/)��XY��7!��4w�y��~kl�x=�{�~�2V��BOY�0/\��c�E�g�Ӎ��;+_a,g��&�����t�5��	^�&:y�>�����@��d��i�,t��2�jn��0�O��a����EF\���T�(��}R;v�껊����=N��F��v��M�a���3��f�����^3��e�e1��e��fM��.&��8-̾��,fڴ����P�5�P3��� 2��{�ho�������.3�cG�+w��{2�����<;|j_`N\i�g��S2~Oi삑Ϭ�}�(Ԛ�&+3lq �v��RnX�?\�`�E��Ԃ@E�L�.� s�"ۭ��_�VB�
��X��̐ø��t��яa31iYokJ�{����\2f̹�˔�@mefЍf���3GD�8���h�=C2�|��9�}����7P���2�˕<���d���g�yxxxxxxxxxxxxxxxxx��}����g`Ͻ�|�Jl�*��7%2����4�]����`K��G�=�!����+e�,oޗ���\[Y��Ŋ_�(YI7�ܳ�%#��ggWTkX��\Ó[B�<�QG=[�k�A��~A<�s��4��!=�Y�|��i��fb��hO���xZB��4sx$[k&ܸ!�1jA%�vя*vD�%�w��窗��ms�����j4D�)b�URc@3(��۞|&�o��Hl���K��o�.�3��;����DQ��5a�|��7�㽱��o�Pl?�������8x��'c{��d��ޑ���?�<�Ñ"�Κ��bU�'�?u�LF�Ǎ���G#�r��&R��'s��iFLC�>��)2ޏa4�M6�ԁ͆(�>��0���fVs���x�ۖ�i�����xnn
z�2f���"��x^���X���h��-�LYψ���<���3np��{sb��ʹL"�ֲKcuR��Qi�M���}�QN��^���yJ1n��q�;)mKf�y��ǃ�DH� �����f�.&'��ۙ�un�ǽ�����\�#p,;���5Q����lw=��=�ЌS��=Y�D�-1�/���l�2>��)��0�T?�uE�Z�Y��N�[���kY3��!��.��i-F�~A�L5��9��*�f����>m�E��Zϼ���n��`h?؀�E�T�Q{������˂=n����3Y���g�yxxxxxxxxxxxxxxxxx�$}��@I´��ʊd�{�-����_��;wn��udٻ�*̿���w�#�u0߂
焋g�ѐ��8���֖h�ܹ-�y����p�g��l���"�պx�� �.��,�mXF�O*����@�p�C�?��@X[Z�q1�=�=���c<�)v��|�qx����Ï	����k#7gvg�	�G��aϭ%� 5Cd[����T�c��B���$��4nߓ�\���;(��t��flYl�+L�j&D(~D��ni<F��/=ۍWD�rwS2��b���ÎRH"{���'�FO	���0#���i�g��q��QФ��Y�>���f"֑Gf˝_��z]swn����<_�>@��yh�%�Tj��k�*���h�{�\��c}^��ٓ����Vl�|C�բf��G��=h�%ȧ���,|�f����\� bl�����ɪ��)5)�hZ��,ƚf�w;���nǼYuVL����N��^4�O����{.�ڤ�z8�b�f��c@��z�{"U����"�s��;|>��v��m�_��V�v���X�2���LڵW�X�s�3��w)g�;��9�q��V��7=�8��3�lM�������q{���}Υ|�7͔����F���LF#��9c�hߩ��$��+��v���=����}>I��`�M�fi��������������������̣4�rzC{�ͼy0�̾{�o�}�fl�!�bU|���xT[-����j�x������Ţ�K�d���e�s�[��wYw���q��\�/��_���O�5����#�:�,}`n�߁��5�ʡ�g֛�����zC}�:�tr�C�̍�߾Ƴ���+n0�H/=����л"���x'	ٿT����y�ђx}dw���$THjQ�s���#95b\�Ñ;��.�AC�]�ҋk���#{uyQ��d�-rwF&mM�&4�.�^�-5�Ca�޺u�:#}=-;�R[-�{0��G�p1+��o8b�<#�Asʨ	��(�7���rj��&:E�?���{��!�vz�<�����2�Q5�Zyed�m���Z�|!�/��f0��2����G�|Kl�}�~b���������C�����ϓٷCf_��Qȃ&�+;(��=F����(󽯝3*rvk����GL5<&g���¬�w�2���
Y�>�l��qT���}�A6.�ح�{�����	S��14��f-N�ɕb<9�;38���j �������������3~|��r�Ud9�5�f��JE��m�Yc{}�#0�\kɺ���>4�p3L�����/j���9sN�xs�+Ԍ���8��0�P>�5�?$�9�z&g!�q�d���+��C�;���=�-xxxxxxxxxxxxxxxxxxx�y��" ��H���F�;�-Zyw^�,���/��ڃ��{������v�d���C݁�<������Ɔ�w�0������h�	�]�̍��ˬ��K��ҋ/J}�=��Yj�1��U���	/b�2�a%�V�Ll6�9(���E)�� 4Cj��Yn#G$ș�hBL�MGAJe_Z뵦� ���Y��	)�d�FS�i��1�#�)& a$�+�^�GXM<#,�|q���(���G$��Sin��S�Q� �����>wW4�~�4�����ll�����Eh_�,��7h�>�{��n���߉�������^l����Ld@EtXs�L6=�'��M����l��BF��'����0���)c��e���������u���6E9�(G��]�Q�f�i��aJ㾬�V�f�*�|����Z�Z���u�xI��h�lߓ�I���}70���;[�%wwSq�*���LzZÔ����a�پY��bԲ��Áͬ[��qp��=�od8���~�q��޾�E�{X�gi��5UF�<Gs"םX��|����>+��ig��vm6S�hLN�h���L�Y!�p��b����K^M:��Z�f������c�O�4)�ZFV�@kҩ�j�x�`����z�Q؅����K� ��L;�r�d��ѿ��aƘ�}2)�gt���b���h�{�C��1��[�)|�����-���i���6���x�>~';'��z�h�r��%��������������������qn�d�͈��uG/f��J�1�V�0�w%+�g��LlW�Uy�a�5�=�y �r�YBA/�r�Y��4((&�wU0�n��zl�	�����|�6�^�k��7��ٖH=5�HO0�|e�w�+L�fGΣ�O����PmD"2Ռ-���d�鈃!N��YJy�ǎ���DrȌ��VE;v��dd�\�v�l7�$v�09Id`{Gd�,Tb�s��Zj�i�2�\�=Qk����\�ƁXg�� ۋ�S�~����O��?��O�?�������46�z�����[�����ۧy*�� k�~�We�9RY=�V��Lr��/*���04�v	�;�G�L3�\HEPN(��7����wT���q#cь�?���I��<&DtBD�,Fw�Ɇ�,��Y.�=z]���0R�>'�GjǶZ��}�rxj�Z�l��[��[\���@#��-<?�`�oܹ#ۿێD2��K�ٲ�/���(�קf�^g�g��̆�GM@�`W囧�z/y?���t3���fY��Ik�r]Yu5N�ђ�T:i��a�՞���w��S��N��da�~�����w�ftg�g4�FP���ٺ>G=�5���~�Q�ʲZ�9Pf��Kq�l��;gz1+n~�j���(�L�B�v��]�d��
��7!�&��<Վf���f��kD4a�f�|���8�Ƹ��9	�O�C����f�q;�}?�wz���3s㿞�������������������qPre�ʚ{o�k�]�����}�����֯�Vl������ul��6��k���-s����<z�u����]�%���޽ۇ��|}x��"�䢜�=��3�ealC;��n�hr��5a(����b_a�)gp0 �`	������"�o�!�F�����k*+��+_5�Sa�\p�>-�3�w2.\�6���Ԉ�q�=,L0M����T��!�w_�����_�{��&c�+ף�eE�m��3��v�P4d{jG5�����	m��0Z���쳟��{����>�֧c��g�ۏ}��C�:�ƶ�Ϗ���'y2�_y嫱����_Ķ����q���)&߀^G$��&X��nyHQ���13�z^��4'��e�wJY�>��N��m沎�������g�"�|�����y^�,�x�5М�{joG�`�1�M�<j���d-h�� VSd�����b-9��[j�4�����n�c4J����7�¢0��My~S��5��ltD�Ҋ|�F3��&y�M�Yk�e1��l8kL�������,�礼�	sG�Pp,;�˺
��_��v�L����"�g�c[�)��K����}D?E_���w���!g,��1�A�Ɵy��3�(yz{����CS�R�Oy�S߃�l��C? ��H�a2`�6�b�13G�zF�������������������9@����jd�JL$��ouu%����ۛ/ߌ��RYN�.���ʊd�[, {^S��u���q�������Qc�`O��-#K/#���E�����6�6��d���X�����r�����90�.	�b�d���S{�5j�)���.3R��餵��GV�i�D)O�����0K�WEqo[ڳ^�&�k���ſ�����E�/�y�Jl���dO���������.�A�*̍JE�#!"��\7�63�1�߶6�Ƕ�j�6�����a�dZ������_����_�vmE�,w�5H��	m����o�[�U�O?!��&�T�A+��,������55t�F3��������_^-��LS�	#���؋ME�Ni�w��Q���Ύ�o{��T��j�Zn��XA]�*�l�$�򝎼�j5��f<��R�/(�!g3�xR��Z}탦U�޻պ0��L� ��Ҋ<�v�����H��ޞ���ذ�+@v�墼7���ku����a�\25MJ�d.Lу?�(�$��+��<i��i�EG�mu��NZθ퐥��B^�ǳ�Ԍ�5�f��p�S�u8o3*2&V�#��O�X������﷓��'}�����;:��`�w�E�;����[�o��v%,�#{�D13�F_�����W�����jo��y��䈋?����v��=�D_�H}Ws&�0%6�4�3�ghm?{C��������������������8�t�eE���t�!p�������#��?�Rl��c���#��ׅ�u�eaD`��G=;+R�,U^����}0��&_ �*�d���z�rl76e������	ck_��rI�{�{+�m0��UX�,L�e�Ge������F�s����8-����EtB�x�Ԑ��ʍk����h!�����~�R�"���va�޻#��~�c��l���Py�%�^�Шk6傥��F���DfI��{����qi,������Z֥]no��d�)�Y��z/Bc�&O�/���~�/���_�L�&Þ��#�)�Y�p;�+}ZS���t�2+������R�`��?�5�X6�G����a���7#�ޘY���6ϣc#�|.��i��M�ms�>^�y2�Q#V�d��
��UѾ��^ ��u���F�,ch���gwC������}a��z@s�]2̺���:�Kڨ�ma(�ٕ�ߓ?.�~u0��Y���;�'7������r��4��j�y�c/�z⤙��'�t:m����ó�����=��7�6%�\ 8f&z�x�0�c>eC2�
X�x�0�lF�a�a�a�O& ��~o�o�5���K����o��_p>��فG�3�"k��}��ڌT1.$�1�UY������מ�������������������qP2�{�#���d<��,ғ�h�홷��ҥK���'?ۏ��o��#��k���?����v��h����0�K��"#'�d��G���췲$�;�ES�̬�%�ں'��&��ҳ:W&��]aF���+R�K����B�&���%aL�\��Ue� F�`�C�lF�aN���wt��b�Ho�(��j	���A�IT�=���gd�Y%B�zY�}��*�cg+
�Ǜ�}�qZ�m�l�`����|:�����KM+0���騬K����t�����[����_���~�w}_l/�Cv!fb� ��	fa�ۧ>�'�����X���L)m ��9	4��N+��D�KP���iN)����j��7�q6���Dƥ������N��6-���-�q��b�&��֞!Czn^��ղ0�=0�={�5a
S��bf����΃1��s`���=5�jخu`3���b_,�[�/-A�'5�4"��t&6������6Y���p�L���j���켡j�7��ߤ�/��5�u}�7+�,���&��G�q��g��4������R�~h�<��>a~s&�t�Jf�^o���c�Z��K�s���h�3�N
|�D*�С�����ad3�ʕ��]F9a�9	F���>��c�&{Ϙ�1��=�$���~<)�2�H~�Di&��<����������������������uWEH�:b��0=���~�D�C����Rc�c�G��㏋}ϻ��G|,����ĸ��R0�6Q�$��PՏ���9a��.�I�`�]�����=�����َڀ�ed��T����r<2ņ�hm>٤͝��l�Z�}h��<.&\� a�X��؞�>;;w+��� m+fyFhfon�E���������)�*��6^|5�?����ؾ����˛���ܳ��ĝפ�>��ӱ}�Ѩ��o�[���o�lĿ���Ul?�{�%�(LW&s_��_�6DN͖S/1��a|f��q �٧�6���u���i�>H����m��X��]�5�e82��d�R+�Z��Y}^��+��=������]�oi�MZf]h߶Pk�_پk5�.��P_��ڂ�����L���R�<�jF�}����-o��Y���|�Q����q6m�I��]�O�O��_���q��?�&��<��>q��|0�l�e�,"u�����zn��:뽞\�h�U���7�y�qO��qS�s���:��}�lų٭Nzf���_s�vM�Ϟ�������������������q�t��	�gL.3 ��9f�5�?ht�taQ���� �v�jl?�����ӟ�dlwv�����'b�ͽڼ�L�FL�wc{�	�j~Y�z��*��YSa�,w`8��@\� YK�`�u#�bv��K��7��&�����<���GdhX�_6���i� c�)`������u��F���f�t�-C�*H����H��?ԯ�^��l���#C����D~�#�K�Мlm���O��O����F�/����|�s�-בŹ�vB�>����6H�oy���������������#��g���^Is�B���WkF^V4���l��i�\ˎȟ
�D��S!՟B�Zgkz�!PZ(���ݳ�wngKvL7�FsS�fWG�l��!;�"48��-шm#{�ɺ�X�	Y�<?2�;x~u:�~�V�.���kk(GJ(�|f���j�&��a��)�qaI޷���g����f��R���8خ�穋��xݙ�A���A��=U�y���O&ejf1��2��j5�5d��jxF����u���}N��ٖu{fݯ��	��Gj�钪;�@�L���>WV�t9���Хd]�q��]���3
(���=�?��C�֐��:��h���
p��ϕ�f��2��{���.Sk�;�.�u�Y#�[:�|����>�s ���!2`N��-��0��+[z��`�G��,�su��?��[b{�0�>��O��ŗ���;�%��Ǆ�w��5�Q~�����,�hU�����<��� ̄ڢh��_� �--��?��,��*�!_0+p���nh����c;P�k�]�yϑͰ��%����E&���G����b���X�S}���P����p���@E��^��q{K��K��l�ߔ�*�t	"�uԗ������c����>��c[_�OD��H�߻���_�\ӑc�/}%��������OS��b��/~J�w���!�#�����QEv�F��06ÑY�����Fd�)�}ٺ��[�x����&�v��j)
R��䩇+���~^�� �����L�4�?��V���"��9yϐ�F��Y^�]�#�j��"�d�QU����<���� ���vÂ�%�h��޻-ڠ.^���\gV�����>~o4�����dm�WL?'����R�ϡ�cʉ�|�ɀ���h3\�E3��y��Y�����3�<�2�&������4sk\&���.F�aƨ������'�yv��32����3+K���0��@�@H�?����5c�xsh�+����S8]?�=T�;f��ۘ�E�&�J	�7V}��7|o���)-?�Բ�ϩ���}���f:�\����U�i�i�}gj��ğ�zw��������������������8(�]��������X��3럙���(�� �]��/_��7}P��n��Jlww�b{{S���0d����$���M����¸���Ԫ
c��,L��_��Kr܋�䛫K=�5P��A�-c"��#hhr ��|��	u@��6�i2s���C 3��"��ANf�훎2֧�3"v�@2g����Ű� �V���fj2<x�Fly}�9a��eUfH
�޹/��5�E����M7�������k��_���]�@W��UI�Y��g�12��Ŭ;���l&�����l�.�b�5�;��Sx�5َ�2�+����A#�00Sȸ�g3¬�4��ɫ�7�q�+
��'�5a��~��N�/x�![E6�Z}k�~��nd��8C�>/��VC�OF4��g�a$+��7&]�X^��q��3��z�-��پԴe��<�3�h�m�������5y����~6�i�~��d=�ce�02�h�x�p����n�iwF�z�l��ܼ=#��}��Y��j�,M�b�7����^��''�9����~�n7�L�{>i���F�:��P3��4���cٶ�i���j�M���+��l��Wif_�Z.h�_�./}������y2����E�wsLs���W�g�yxxxxxxxxxxxxxxxxx���~zx`�vvXbH�M�1eQ��������K�_�z�D�o}�����AC�I[�۱m��%�)���8 �fYwk�¨��	s`�ϕ˲��֪���`�E�F*�Q?a:�b��rJ-Bf��`4��m�Z}�M�T�ɥ3���G�U�PE��lB�1�d�>�8idE�H}����S�It��rj�(f'o�0����.2~�iy��-C� XJ"��k�nv8�ƕ-5i'��gy~�&.���:r��9SD6S��*rˬ�[�ލ��U�2�A+��� E�7���V�k�I롯�Z~߷8�7�{!����z� ��2������!�65�x�1�mL8^�����:Єd�q'�[gDG[XF��2�Lm���oo
c���tC����h��
r�{RN��rM~ow�D�㼑�g�s#�w_xM�Y��Dc�\�ɐ��y�E�g�I5�f��yOK�5N[�������<ӌȼ׋��Y�>���}��wҌ>'�������!tx}�}�͖��j`�s�G��	�q^���{��F[3r���q� r`l�j�8u��*�O3��b��N�֯a�a<S�R�G{��Dü��3�s!�9wO�+�aP8^���)~�Қ4�2����$�U~&�O�}� �їd��*F��6��F=�� �H� �T���ZwEd����L8z��Qv�h
�_Y�m�-�v:�贩�g{4��[.Wd��50�`RA�o_�,�}da�p>C�ݖ�=�]WY�xՄ�	��jƘ�g��D*����µvh8n$�WĜ�V�(GG��oJ�������ʭ�n����bM�_{a�D*`]���g����Ӈf\�(���[�7c{�5����z$��w��1�٥rc���̠;�,7��G����#��r]�q�Ț��֋/����/[�����}E0����c�л�������g�3�f�S��~?�V�S��>�I����v{?�E�.�r�.4b���낉�So��!vehʒ��������e�&ϐ*}����Z�
�l�{;�d���RsRGr��wqa�:�JE����^s�%�Mj�ݻ����o�0N#g��Ҹ��,��qec�;�8�Z~�)evE�q�_�Ξ���jf��?븧���4��=��n�̲���g1�ƅѬ�{/����9��U��v������<���=�=��#h��������F���1$���f��� �
ܧ�l�g�)�f� �ʏ45��$Y����3�+��������������������8H9���������h3� 8*9�x`�~�V�6Z�92���}�/�)�\����XM�F� @6�.w�>c/��4�`��b�m��a4���h�Y��-��Q��ӝ�J�ckc���V_v���6�q�Y���̦�#�s`��Se�
,�z�|k`��|��ؾ��0�����������ؾ�/̗��d�$���WԃFdSl-���ȿ�ò�|?���O�~�p���؏Q�Tkf���Xr��WE#��/뿺.�A� ~��0#���\����� :��Ay����0��e�?E0.ݧy�4�2#�cj��e�iD�F�]Z�5g���%h5���uf��w�:��Z��z���ߺ���lI���uɊ�3�̕ZM��=kG�|���&��}ԇF^�+��{�H��aa��Y��_��������A�l������b�)���X�MM�J]�{{V=���Ap�w��㤘_y5�\�&}Np\�3�h�i֌�����[~�4��E����
�}�c\���7+�j�L��Gu�Yg�u1��{�pi2f�/�e�E�o �xY��`3�U�����9x����-����h�sx��IAƞ��K1�f��=\~���>0/S���e�qA�����������������������80�>gćL
�JdD�lamO&�v\��+��n�|��a�{X`9Xf�YI�1������ċl-.�����l"�Ѷ�t��u6�4�R�_�'�qg�Ϋɥ��R�"�����[�������k`�lm�FUV�G	46j��~�ya
��_���'���������/�ll_~�b[_��a��׮߈�O��?����������/>��Ҹqj��GMa��DV$��>լ�ef;b��p���(6�L=f�_F�ޖh���l��1��l��",��NG$,7���`̌��L���$����z慄ߩ�I-Wc+bMo�����25�L���@&+�ۡ��j����!4`jua����,ϴ�Rh��:}�7��f�<����	[�.��9x��],�	�Pby]4u76�X�	���h ���\8�l�cJN��q���e�L�s7��#�8�jM[�Y3�\�������9��^Y��4����w\&��~R&ᤌ�q����1��R�LeK�v�и�˂�?�����Z���v��{L��'�U��Y�;��\�5s�gt:i-]2�ۛ�(g��2.��C�	8��L�ӖM>A`�H}���b��8��9��" g��g�yxxxxxxxxxxxxxxxxx�$���ȃ��1�Lt=۞����Ȕ�ba����+Z�drMdŎ���hF��"vdؠ̶j���/$�&c��.���Ψ~�ayX�X���+r���;�6�Ȓ�uW{�$�)M��������4�� Y4��W��?���~���獆0g���3���w|8��9N}��Q�^������7��7c������'�a�>����|�EXQaL3 Ro4���E!-�� ��cٵ�	$qH���۱ݼ)�6���^�,�מx4�K�=�ڤ��V�	h���8~N�ÌO|f]NFތ���"ŀPŅȾNF�ە�r̎���/�x�뢝W����������^|�D�2��fS�׹9a
�b���%�r�����ҿ�X^,[���]��[����#����z2��d�4wES�>?g՗�×��+�=ڥX�v!D�3��s���ؾ�G���v����u�\�SpN)��f��gL��wm?m�ü�{\z��f��v2̘�h&��Ëp��Y��Y���?\�i&�f�jﺾ��`b-����B�l朑�B�%��b�5�|ธ|���ͬ=�L]~�qn^���d�d�3�q��Ad�W�gy8��3c�)G��Q�B�:��15�Ew`{��������������������8(i�e��G#����L
�҇�Yi!4�ɡ}��^R�P/fUU���gu�x���e��KQ���c�gi����8z~By�*���
��Z�vd�d�Ekw�����P�a]�`�}a�����K��_]�m̙D��������Eт�� �>��w���<��ኔ�26�2K��1e䯱#����d��Y�%׫�DVݖ0/+`zuZ�Ȥ�Zl�y�8��2��6=�ǈ���A3�����pf������яa�A��0�B󞱙�F��d���~�{��aa�������k�0�Ȩ�}qI�{��y�PK/Z\Dy�&h�C�����f`��Z��e������{���F���l^F�����h��e�~�b�A���5:��>Y��ĴY=�)Y��Yi��ʝ�8��Pt2��k������T�j'}}43Q�>i��3S�փЌg�m�743�\�-Ըؘ��!�3���=�>��2>�}����FV�&?���<��^��\4��=3�qQ���oU��f���4Ug��Ӛ�Z{�Z�z�>�(��z�a��[�g�	x�b��<�����������������������1�`�$�t�a,��lO�K��h�q�Y|U$%���7V9v� C�+5Ŝ;� ۬<ޑjwf��ڪf���y����&�����nt18���v�{�	\�,�hfEEY^��n׀�W�l�pQ�<a��"٠W�ѳ_���}AE�M�c}�Fv�#�F��r���_#�pY0*9ѹaN����2{��>v����3o��ƫ��6@��b�d�VGQ�9a0C�>�tk�#�ʒ]�N�>�?��"�:��\���d�嬿+������PL
C&p �&��}2���y��2��Y�#����<�߱~��� d
(�0E�m�0���a��^���Jl�nyY4;`�����5Yx��X\Z����FlKe��W�z,�;����s/I{�!I��*�
�?�l�d�yE6�G��9�6r��V�������?���d�/��)0+m��j�I1��^_W^��9k�}���x�ߟ5���I��.W�-]P�+����Ζ[TL0��:o�#���Pt�?�,ݦ|����.^���M;�Պ��A_�|�U6k��nf�$b�<��׸��}��gf|��r<���&���fTk-�����Er��w��Q:�������<�l��{b���g�yxxxxxxxxxxxxxxxxx������D�s2m��p��hm�6��q����s�"�ٞ�qIGֲ����fU�=�Gyɫ���wټȫ9r����b�v�#5Z[@�P�c2�L�!S��ȂEvue�b{�Vq�H��AAh�c->��}�.W���Ԛ��;�
�����呵b��G��%aP�#�25�z=��R���C7b�l����׍Z|�G��뻷��`��Ky%0�旅iF1]�r�گ����)��^�{cʈn�B;"��_t�e� -;�`O��m0�Ȕ�YY��z�י�jU�o�;��"���$���5�z�}�G;��鷿��
���4!�]8B��ݒ�,�����<۝�*^����5a��|�9�?ԑ�,f�+i?G��¦N$��*%ǀ��2���h���z�ݬ�}��3Y����[���YkO�1���4�kVӼ�so�rȔ��[de�>��n8�ؤ(~z�n?��b��6�����Cc��w��	^��>�߃�c���ފ���ff�!�{������|N�����M��i��U�;)c���v�3i��io��4�ܜY�~��9c/r>T}F�g�����9p�'��g�yxxxxxxxxxxxxxxxxx�����fH�,�)�2��a{�ӑ���G�F�?��y�]��V8|�q��,=�LV���#r�#g:�6k͝4&�������5�u���+i�{#Tm�<-�I��b4#U�*��$=��O�`2eBgKJEZ�sJ�p6�5�T�����6�����U��%T3��l�ܟ�p��#���[;�r���P�#�*��4g$塚7�_{1/�o�o5�I�5����\j0F�F��ͺ�a;�>E�7��J�&̾vK�-����tI�ʵ�+�f;����jA�z�_��v�����r�%����e��}�c��%��}X�_Y�Ku9.������+da�x�N����\*[ڛ��`;.��d2�r�;��㎣�gY8��s�i������r19�I�fo�ӬpT���G�]y|�V>���'��f�M��ļ�|y׻������Fj�ф+��ߧ����w"�*��gj�gY�wx;�e���j硚	��q?���#e��I&�3GL�ѫ��8���2l��,��>�s���/�\�6W)��.Xg�LG�\�ռ�.z��$�)ЬG�Ug{�O*��h��6�7"����#�d��#���:�Q��~wgL��c��ͮ3�^�՟T�Ɉ:�!� ̚*F}hy95��f0�,`I���5sx�u�M}=����P���߸���[��V#i[w%�nͼbZg`"�-P�MЁ���իR.4�6o�.[����ދ�+�c[��z�Y�E=��P:"X��|�ٗ͜�0�^:�W�,\r}��vg���bӇ3��E��Z�l�u��i�����V��ن�c4��F#��Z\&�>���B__�,�d�{�c��V[�@o�~W�kb���u�E�GsO�y��/�vڑ�����g�"巤�>�C�dt�uR�Dg%O#�}:'��w�"��ѓW�/K�gV��7���I3=�2'�-G�+'eF��	}v_��`�w�^Tf��w�m�������y2��R߳fF��]�B&�}��QMo��)�q5��ЊK4�e�rIl�\��e����q��8NϜ͸�V�?/���"l��M1�\Z���V��=|�����ƿ�[xF�������������������9@��u0���e�@  ��IDATHɻ��}�XQԚhF���sz�'���͚�#������!ӑ��sճ�?��i�*��I���4Yt���߳�{2-,�)`3�y�u;�p�d���hl�8X�d�FKl���'|���&�e���ȃ����0�Z�`
p=��������6��۹��ض�����{�(˲�<��S�S��UYYswC����h1�ɶ�-Kb����-ɲ���x�v����2 i-l��j�,��t7=�S5�5WfUVfDd�o�3����ͳ�;q�{�u�q�w�s�=��s�����${i�j{�[aYD���5a��f��5=?�j�y�	����Ո����s�4'�y�g��#���a�R/�<�EdMf��<?��=��y�
`�2�.5�9��8��>�KKa��!�����}G|&k�"�2�nY����._��O&�۾�=a����\�@g�w7����E�ws#���/���q*��Һ0n6���=�)���I8���I�?*#�b⬈����T��~cR�>�WR�kB>(����{�A��N3Ѕ�侣�.&����̯
�����F�h�����J	�@0�)R �/�������D|����R>�i�~.�����%T/�e��㿕�sa��z�M��4�����/��y�	��s?{��������������������8��З.f?��.���6��ڈ3�]W(ϐ�.��h�~P<Lo5���hQ�Lf�b{�aH�NFk�e����� �<�v0�9�N�'�m-:��CJ�y �qks���еGÒ�VS4�n�-3�i8��k�J6�
�Yx��8���9|/���5�z��=9�cnE[A�l���N�q<&�酪}n�<���i�z�r�� ���W�'�h���WS��gmJ��~G���H�=���K��[햜��k��Ȫ�����e��(xzYv:��<w�JX��3���mk?2�\��轨���t��`�M�հ;�H������y�+��q�p��4�������l�i�=���H��ԙ������C}�����g��}�����h|�瘈��6{�����cV݈�W����92�>��H�O�e0+������|C�_��B�7p��[��x.M>2�]��}�k���K�ׇ3�]�#�9��T��!���nI�
�}�Zo?4�ul}�=��]�I;�Q��}g �(F�L����B�����-�qO�sq������d�^�?��TƮ��d1�%����曻���q{�'�=�y�<r'�X:&�FR{'1�\ٞ]���G�_D�If\SC���L%�Jc ���>����=!�l��Ag�p�0��pܞ�u����؁�ۗYK�f%+)����Y{[�嶰��EdO�"��Ԭ0��ua����+@�m@ޗ��y�����9!3㸐U#{���c�8(}����3+�]}_���+�ò۶��J%a��s�ͶZm#��ߩ��}nr|jkv�-��^�-L���f�E���֔��>�ߓ��_�~ڇ����,����迃V�:�~�"G=��X�W�Mb@'y�ORGL�R��I3�'Ղs}?.Cp\���4.t6ec�����.��t�̽{�r���j���P3�l�{s=ì���&�3��~O{�����5j�1"#��P6��r�Q��tkU��)#�|e���т�z�̻����Қ�͘���8��k�{�O3S9�h��4��<Z�<v۸�z���?�y*W���Y�q�I���ޯxߩyO�#?�|Yev�}3�7Qd֥��D�v��<	�/� ��fc�8m�G�-M�v�t��T5�@1�hi���`t)*c��Yy=Cu긘-�}Ϊ6��Ķ���v��[��<b���#����/_s%���Գ��;��hk�߼%�;��/�f����J�/��|	Y����4R�1.#�A�J�;�>| k*=T�	U���=0�����r�gd����Z�p1,7p:ͦu���h��.�~]'��M���8�1F�f\�v�/_2���X�����Tøl����;���0�U)��B�fK�e�O���7��	�`���^	��ר�����}y�_���7��)���8 ;�k�An֥O-�X��d��A�����]��d�w�����>�c�qTô��f��/M��jq%1�\pͧ&e�Mz��8�L��8Z��pV��&}ކ㎏)����8)�b���U�I1L�牏��n���#f�bb�?SpDn(�۬dVd��0���1r���h�Wc�Z�
�2"<�0�f�gq9�4�UĘ���z�tN�Fmq��~�:����x�un�	��p���ڥߕ�R����d�g��f�nOڍ�۫�3�Y{;4CAe9�����~�|/���u���b&b�:N��ubG��>�3��/�ew0�4O1�"-���ٿd����/����1�	7(�]پGK7�g=��Pc���gi��H�=ZX��x<O�IiV�8������v&Оݮ�h����������h�H����9���\�y�I��NO�e}o�ڎ�ݠO���%1T�14�D@Ř��|�)���h���8���Ҥ�u����j�aF�W0�8��C5���o�2�!�h���WC;�YU�'onI��n �+�C-�;����L��[mV�C�_��h������t�:�d���mʽ����m{����e�M��ScJ����&�K� $���,����mɲ\\�l�� w�ϙj�v���;��*A�e�6��F.W��g�O/�>�g4�nS��{R�<�|~��/�coC4%Mv8�E�+b*@����0?d&�����ԗ�.obFw��@���O1����Cp\ZvǭM�6���=<�u%1�4ck����j�%͛�~?i{�T���몧��������Hj�I�1=/>j;'1���=!�M3]��q���B�2T��nx��b�})�ke�6�4��{�j鄈2��Ua��G&�Q��㼳���প��դdV]λ��#]��g"+p�r�`}��|L���h+Sk�hM˼tw[։�?z�8jb>75-�Mh��q7��^���j�]� �?�uJ��o+r�l�J�b]�E�2��h��yf>lkۑy���BF��.3�-<h�mD���О?&���z����[WD�ڏ��b�d}5T���>�3�Bd0�6oe�L L���Π$��ζB�'-�Þ�%X�;`��#��Ζ0'��l�%5�8/{��+�ͦ�,+�aY�����5�m������L��gvԛ�nh��l�6&�Pz&� �Vaܣi����@�~�`����de�E'3�c�bĲ�*m�$l쏮�&���6��W$�&=9����㏆euf�>�:^�c�x�X{�����"��S:����v=G�����&����'���hȭݸ�ed[eV�NSƭ�K�2w����ˢ��q[��L,0�Z-�Mu��E��P�.m=���y>5ӁY�L�1���Bkz��c<�����u��C����l�<-�,�[r��𠮋��̢����z�P�װ��1�=N��/�̿�ܼ���ik�kW�̾2�d��G3��%xh�	7mzb����ԟXF����v\���>�ŤL�Ӫ5GF�~��|H�D�󞳮qxT�kM���%ݯ�~�9�4��d���9Q��=����Ȓ�Bv��Y�������d�5�PJ����b�"���F�������KEj�PĜ��	L����+��G&�\�F%���y���H�ψ�F]�$�]Y�u�2?ۃ]e��FX���Ze�%��y}��`��7�"z��X���X�uV�~E��A��rYڥZ���=@�J��N���92��j��E�ס%���>�;���AQ����<���)E&!5�X�G'���3�<<<<<<<<<<<<<<<<<<� 
Q���0&홒ɧ5���
����K��-a���k�ay���a��#1�]X��e���`╤��U!/kZJo]_��b�T.��t塰|�d��G��b��e[+)���מ90�{n�13�����8�j�if_t}����RaF�������ڬ0��c�}%h+4��x��xr�I�1�5�!Kix��T�h��<�9��z��f�b((��R����|��D���իaI;<]̶������χ%={Mxޖ/\˝M��Z}�2�L����:�����_��'Ò�Dj�[��.�+�O����V�c?�Z�.���{���N��9����x�v�[Ʃ�k?^7$�b��` ���8�y��y���r��2��٬�0d�����/�l^��`\�)�$��?��a��g>��G���v'��Dxl5��>f��#���j�-�l?�2�y�Y]ͬ�,�0)ceܬ�f��H�#��i��&e �/-�$L�47k���i�i��G�;&j��ZO1v&F�y��*}t��k� K�+{�֓C����c7����L>����ey������n0�
`�G�:2��5WDE�G~6A0����#G�Bͽ��>K$ɝUYO4�a�ir?ٮ���6֋mh�u:�22'B�X�7����O/^����|���qn�j΋��R��_�*ev�"c�d���r�2�;{���[�Oy��(_�����#Ά�oԎ�u�̺PϿ����)���j��s�~�6�>�3 c�K�p0�
y��SNJ��L�#�g?�|��_�՛`�����q7�(L��Y)ϝ��ՊX��e�hoѲˬ�}a��Ȣ����,ޯ��{�~.�E���°)L1�~�2}�G:;���WiK)-�q�����3ڣ���w��d�x.-2gV0zl� 2�j���u6���Bu�o����ρ������nY�##��[�'0Y�lM/��:�	��f̦��1ǡX�]�1A#Q�i���+y0��ٷ�ہ�ȽM񔑡I�j%�A��3o�
G�Q3M_W	Zd�mA����3�z�}xà�e���l7f!�֌a��ZL'��c=�Ѓ8��4� w��;�ݳ�?��uc0ӍV��;f}o��N��.���K��Ƿ6-�ŕ%�Y���RS��>2ߙ�y��Z�'ǧ&�ֆ0�V�=�t^xL���<�]h�L�cQ�61mP��x_��7C;�}d��^<ċ�=2�Q�����!�;��Ye
iĳ��߻>���C�|�u��f�=hH�l׼*���=#��YCz��Ĵ`S��	�}i5?M6L��M+���P�7���5�bD���89�2�]���S̳��̺"mď�*��Q?�͕eN1��{C]7|���=��\qM>d�ż��*0��<������XCfޝU��ܺ#����m�e[a�]eI�?7���ך��5�Rn2�L�FS�%���W���ܔϕ�h��l�|z��bX^z�~��W���|v�G�0�7E˺\�v����1���پ���̼��L�#����zD��z�_0���ʡ��c�&<Y�w2�̰�z���cwZ=��������������������`lC��bCc��L�<Nu�5Ѧ����hX~�ӟ�&,ЋK�Vy�0�.\�҂|?]�E�(���~T�����Z�bހ�z_,���X�_N���X�/=&����������?&���y�06����|����E�pB��#c\�����I�80;z�虲�����k"�nmJ8M��sW$[�a��f�Ó��J�lC�����|������Y���>��R�Zfܮ��q�(���lĤ�2�^�w��<�	����`7��sxL32�xJAO�9dٽ���aI�a�~s�K�]�2�n��2��$�r2H��K���U9�����C��GKj�e�������;�.i@E3�Ȅ]�{�������m��ڍ��6Svm��u��ov�SJ�� �^f	�M��(��d�����i��d����u���Q�3˜��4�5�њ}Á�\m��<����Tv�Ӛ}�����L�	�f�i�x�!�0U�9�xN;�3��.m���}���(2�d�C�COZ�Og�4�g����F� ��}���?��0;^��SRd�ac��<$i��|�_�3ң�,�L>0���Ps϶p}�������Y���z��'��AG���HDHyF�o�b�W�y1�}�3#P����?F��K�����ua�mo��r��M����4�Gλ��L���m|/���9�W��[Z�����>"V�4�d>��H;���4���σIIP��/��G�h��a���v�W��Q3�!j�����?S>z�g���3�<<<<<<<<<<<<<<<<<<�R�4�O3�rNǇ���K7��3M�O~�²��s�E���k�����riQ,��`�U�e%?Dl5�J�'�FPY#��O�tAR3Kr�fM,�;X�_��d4]y⑰����L����8��6����Ǹ<'C�<g3J���\�1�����q�x{�֙+�"��>���Ok�8�[�Y�w3Ъ<�۷����q�e�_�����m�ڢx`ؿ�`���.̢~��&�K,dGꀙf����`��9�T���Hu[�Zs�	��o���9����JX�0۪9�l���Ph�e���2����|��@���Λz<S�IG�c�՜�x:��+�ˇnGOg}����cv�A_�j�|������x奰�)�
�C�~������S�%���|��&�W��1��ɚ��t�s�O�C[[�Af\�ȸ0������Q�ǵ�+���QUg�sxZqڙ7��}���v]�q�K.��g�_�{}���q<piO������q�G��k=1�]r��yq���^�L��� �٧�e���tW$coOM>hrsɬ�d�i&牜�`��{�4X4���_������]�(v�j�6���K�R�V�{��f�R�C�L�\V����H��v[�7?�����8;�u�Ғh�mm�� ��w��Jd��o{*,gjr�����0Q5Z2���wWڡ�ui�������#s��c���XF�fq���hB�(u1�>E�K���M���<�k��������������������8(��X(�5�r�w��7_�X�OJ|���gò�X��E�z���a��â��0'���)��fz`�ud�,4�hQ7�0�TۂeUQ[2���Xpk�lWk����BVÛw�ݍ��xM4�斅yhb���0̪Ʈgl`z8L�Y����h�vZ�-��:�fn%�h饼�_����d̾��R���#�o�L>h ������������pEhs���Y�}�2����b��em���a��������7PL$��w���Ќ*�M4�)H��Og���@Rh�5���ed��u1ˮa n���l�����b�E�ߤZyZ�0�q��1_?����,����i��pws�ڞ���8����������^�q��83/�<��D���>����	ZA1ϟ����(��N�΢M��v[-ڷ[�&v~�&=�Uh��KR�vVڃ���F�%D%ew��{y����xI�r&�����j��U;$��FR{��>����f~�z�Nf�a���X;i��&<Lֿ'F�����~�9A0�)|�L>=Λl�؃�Q���~eD6i&#����cuUv]��c��u#"�¤;ؑ�C.��/̈��R�uB6��dy:���M�o����lͺ�ݖ�/�ad��>U��:�<s�h,`>��*9�%���C����o����ޅV�瞕�ۯJ�Sn(�)煙�)��Q�G9��d>�j	ïݙ���C����޿ Y��#��!i�f{�or���Ȗ��ċ�w�iT&·\Ve7�>�3��>�yd�|J��(��2��/>���ا������^����|[X~�;���/H�Й*�� �	�QҲ�3�IU)&F�����(��6��MB�t��=d)ܗ�ظ)ef ��ڼ�?_��?�C��+-1�\v�Ա�J���Y��<�_� 8_v�'X3�����}z8X��[�  �5��:�l�%d[�i�i->u���ӣ�`4������Z�|��>�ŇxxB���n���Zc1�Bs<VO6(�>�Z����<����1����yDgN�����rj�iFF�pF��4�p�M�ٶL�mh�u���Df=�)��_���'��"����K�u���	����z��﬏��
�z���9h����ZX�S,	������}EMK^���D���t뻒%w��L6f]��q4�.z����S�ǣ��dT��:��u�h<�������(�~9;��f2�zَ�WE�2��Dk�Eڿ9��i��֔:�8*���\ږ
z<�WYO�2��8�j'S�3bH����vV3?��̖R^f�.9\+g�I�3�����U���q_�l���k��z4���W�WU�SC��E��1>{�e�}���#k��R6�v�<�eY���r���,�'���e~ׄ6t��~���"Pxuj�ɉ�U��;Rd�}��*��4"/��<m��%��\�$���s����%������g?�[bOy��Dv�q�f]֩�2���v�#bjwO��M0 ��=8���1a^Z�:���4�ϸ/|�u)��aC�궘��d:�t,�\O���g��3�<<<<<<<<<<<<<<<<<<� b���2o37�Ƴn[8v��P)	��g����п��������o˯}�ׄ壗�r[+�%8kL��B��M�d0���e�0�6��O-ֵ���fuhh��e�B�aA,�K��E�\U�TAN,�SYdw��S���a��Uf��ٌ1��gM�9i��fx�����t��y�4�.2\�f�D'PLM՞�����Â�g�#�c0J�,����4��臙<=}k{+ok��X���<h�rU��<.]x.V�E���0j6��WF���8�C�0�V���Q�M��<��y���F}jǑaS���kw�ȱ���
���?��6�)��M��a4�0�?3����Z)�����qw�7�ߣ�K�C�Q�[Y��f�����%���h=��2꺒�M�&{�&�v˕�>l��[�k15'����Po�}A��j�{�㋁bȦ�>۟��h2k������7�j�x>����f_Y��=H���y��PD{MV^�z�%�n�a���h�v����^8'�3�;⡝��xR�f�&��q:q��$m��>��&�?��y\&_�z����Da�$n�1T��l�*�Fk���l�pF���3[�C�zbL��͎.�:Sk��4I���Y�ǵ��� 4��z�0�0_3�Q��!����؅]C�'A��@"#��^��:�Φ�?^�u��@2wY��u�����c��Dxq�֓�ZM�'N͊�c���%�g�s�� �h���+����ֳd�]yD"c�����?�����?���R��|�s��s-�S,���z��u+�Mwd~_,P�P����
v�1�X��˒����'��l�a5z���53Ͻ=#E����}g ���fFG��L&����3���~",_��+aY+�����O��׼�O��Ջ��Ҵ0�K�ϒQ�x�< c@1!
F�H�Ҷ�3;OLn�Clw�)���X�a!�T�b]�����BX�I���ѕ#v{b�.���o���Z�D0W��S��%��1�eh�,="vl{vt�JQ2����J%9� ���� L�"4�����oL��/��0����LF��|���ᖃ�}M3�+��,vk��a���?;%��fC6hlJ��=Z�N*H�E�mO�D�	l�~��h?`A��*h��@ݧD�����=�.����S�A�%#������592���P?�Gu���WyB�n���]���Y{���I�c��1��>��,#w޸%��';f<�:볋���!���ߍv���I{������rE��;�~j^�"���^�Ws9��G�x&��x~����j�q����= C�0�sv}�n�Ϫ5j���w��²�jg�"\YG5*�~�x����x�d�'i��Az�5�&�ZF�f2���L�Ӎ�����>&f͞p�i���_��V�WG�D��[�s�m��F��x��?�"\��Ԝ����<�aX?e�u�Y�|�� �-�����>�4���4`_��b]�d��z���#;-پ��
5����H}��?�Ӑm�ǩ�Ӯ-zn�̓�]�&�Wd?FJ���v��=YWw�@\Y�u���lX�Y��K��Q)K2_�~E0����͎4���fX挆�ỹ�EY3�)�741^6�oh�K����~r�jJ$�G��������������������q3��=�=ʴ���Fߧ?�Ga�ʗ�ˁ�ba��w�C4�� ��"���E0�^,"�Z�c�P���LB2h!2ڢ���,��U��F����=2��E�~n^�����̰bݻ`Xt�x��2X���P�KYvcI,P�~�\Id�Q��������}~��AY<4|�����Y�����)�Q�'��-+�;zp�q�2[�?4/=$�֧��DX�x�U9���	8�&_�Ma�\Y|Ժ>jEL��v��I��_���k�.xL�i�?W��d6��h�Uݗ�+km~��M͸pi�W���_���M�.��F�6i��7.=�HX.�;����U5��wL�j������Ѩ��5���痢ߔ�-v��x�\m���}[�e��[P���_3�d�L��(���M��{ЖcV��?��m��<�I����d?�ߗ~xgmUη%Y��x?����x܃'�P��!�o
�};����sf]#Cϭ�f_n4���eC��7+��Ez�!~'����t�}�_�⨌�Z�\��NZ�Z3�~3�����i�}�چǋ�2�b�'s�����=�*�"��OcW��mJ8^x����-���B0��Nd�Z>Gf�Q&��^f9�C��g�A[>����ە���ڗ�b�@�mD:�9���l�&n�3�Ku���Q@D%5�h_a�[	��9h��S�'/̉���uD�";��Kb�M�<)A��"��[]����e�[�KUeJ�S��~`�M͊�����F�<u�@�͌\�*{A�"�Q���a���?���	r�Gӭ�E�x:�p`�F3҈{����{c��Ű���m����+�ѷ�!L��y:,�z���|��n�ք	P���/�#��0
��&��1�`bQ�ZA���<���6�5FK���
���aRU+R�"b����]$�[sc{G,��@,���,��r���7�-�����q\�Q�����E��]8?4�X΃Qbꧨ-��a<+��%�,m�=���2<u�3�m�v����y��հ���P��������J����`�L Q����1,/L	����e���U�3<� �E�hD �0�����\X��x;P[���&�F�ϡ��L�����1iMu�HC.;r��[�Q"S�ى�}�6���RX�z��y]�F�S�;���/����1�"I�JK.P���I..nZd�:V�{��_�V��8�*�w��T�xu�B�4��D���,��a���C�8S��r��E�/���u�!����E�{�+&+��<��w���'s�����_M��5��lf��wC��
$x��!���w2KuV�{�#3�=����ׁI���������7.��m�zv��������2���w�p���f>G�����^�ִ�|�Z�9��횯i���i��H��j�[2��[{~�yM1��֓\w���ɶ��Ym�\̻��[�^cWʽM�_5�d}�n�d�?�	I�"�?�i�\r��+��M^lW�����7SА���\�D��:��wsK�Fu���Y�s�w��D~r~��K���IG&��2��R�iD�dq���O�[�ۘ�G��O���u1���ǩ(�Pkoj�����q=��������������������q����s�쵰d�튥���o����N��2;?+�v�y<,g�䫖��J�7OK˨���&��t�~5�ȼB�@2�z̪
���X����a��|���,2(˰lS[���TM,�ۛb�n6p�_Q��E�\�,�� ��<��j�OJͰØ�3�獞�^[�|��܏�Ma|�Z���/<�_��w�e�.��K_�rXR��p}U�&eh ����m�����[�-�o��o��e�������}�)S���yx�m��ƫ/��h��q���������'�:+���_��R��#�+�1Wʹ����
˥ea�=��_�64+���g�r�*�����/,/��vyV����ȲT�=�̖F3b�L4�%A��pC�ty�\Y�b]��W�ɩQÿ�:l7��	�hЕ�9�(�Y�J�/�?;w��L��#�>� 'j�B#ÀF�Ui{�����K���/>��q{G<�٢b2�Y�o��L<g�sX0i� #�֦��ޖz������"�y~��3��Q��L3;��o�W��kf_�d�=\�/o	��J�(��3�?��.����:&�e\yf��p����j�{��U�$����6�n��y�i����0�!;&%�y��!'�ɦ��&&k}&S���'�����Cv�gW�HGb�e���{R���`�r�>a{F�0P!��]���P��#K���;bgh RP1 E6��%�+���套^����̫��lC=�Ϙ�7�#�T�3B�����Fv����A�b��hF������I�M�9�ǔ�������v8۳Րuw���ԫ���(�k��\P�����x���д.�~e0�<�9�E��맡b��6xF�������������������@��g�6ӌ�e�w�œ�ګ�eoG,�s5Ѽ{�[�",���9Wɋ���#CKi}�t���ya�U�|��>�q�����V���{2���yS( +.��2�K����v;�C���}FU1��b�(L�~]4b�e[�k@��E�1ģ��}���c�O�=�1e�g{JV�M�_=�RX`�0��ʕGY,�7�q��ۑ��ss-,gf$����1��+������ΰܭ#F�)TsnY���)2L���;M\��je�3R@,�v��3��l��9����x��S Ӫ�+�
<�����W^f�o��o���^����<�W.Hu�	1�MVk`ڞ0���f{1b��G��;!%���u�d*�C��x��]�$�Mh�ƾ������~M�F�Ee�J�����{����1�U��l���``���0;mL���J��Zr.m��q!����p?�v��h�#�
���?{�U?>�mx~��W��3J&r���O�Sk�Q;�0Yo�������i��9dc��2�����3�֛��6nvݤz%��~��w��цJ`䜶�$N�A���NsScx\�q��^k��q�|Y5���iQz���%2��Nm>2�����h��f�%�+�u�+$'!+y�Y���sMt\�<�	���F]�ֶ+@s�v�u7kk��:4��Y��5d���&댭�����u�U��\}Ɒ|��'�r�6�t�+bw��G?����F�N��$�]Pj�e����Ԍ�o��4�#��`�Mj2s�G��]�?��c;0WQ?އ&���BF`���q��CV��^Ǔz��r���캸{��E=w����ɗ/�^�]�%�?F��s|.�8�n�e�m'<�yF��������������������!�>�1`�4Ģ�~k3,���"�Ăy~E� >��X�kE��3�eӳIKt^1ԯ�,2�2F�{e9��R���9\=�������+�ר�:���m�8S�\��V�b�}�&�ؕ�`����o��sQ>�����3������.��F{����{�׼#,�}�8/���;�_(� ��2+�~W�Q�V�L���x$
Ђ��~2E��Yh�!�͡�gq�
�Uv8�d�~��H�E�D@�-T�	Z�Q"����hl��IS.
#�	-�<<,KK�T��v�lAٌԻ�vȚ�B�Gp��e4	=0{�����s��Dh�Sv<&ٱ����e�� ���ԃ�X�g���r��_��{[о�u2�4����x^��쨢/	���d�>��=)�o��\쳃1�Q�ս�<��l��]j�Ę����G�xP�<�Y����0 ��5��1L񑒜�̺:5H1.FYL�$���O��G&k�ϩ�Ǭd���]�3C���fB���nn���q�p����
��Xri�e�%ݧq�`�b����{��̾�>����͊�>wN&_�~x��CV�W�ḌE��&!��C����劔hg3�i��o�Z�ejպB��
G(�����|�dZF�WF}����^�Q�=S��8�=/������IN����qK�h���;wd^�;JZ���D#c�_�ְ���d��:�	f[�&�֥�9�-��ma��?�ð�Ӿ��	���cl�غ>3z|���^�hIJ{��`2ҍ����C�/�d�~��c�H�4��~eN�.�;[;h�o��zU��7�Yz�2���>���|�:*efץ�����cn	밮�N��ř�aBxF�������������������@A)�9AC}_,�7^}=,w�x`�g�|:,g���C)���C`kx�aY�2i���<���b�����x�ŚYK��`�aէOK�-߯�m�F]�����e�*b��BSCLxYx��~o[,���H�ui�Vb�#�5��0<�2<���1�� bk0�"�o@���P��G��_F��7��`� �pf����a!3�������Y����`�Rz �) �
��;4��}��D>[�Γ��#�7���t��p��d����~9��63����]�d�a�R�Y:�Y��@�bf� mjo�hg��̀e?�{����d�5�$��7:ۨ�0�sθDcfR�ŜS����x�}j�֬ߧ0�Q�bw�{В���9�aS������z�E:���/��0����vQC�d��g����?.��03�{�o�_'���"��~cct=�t���~�Fh���l	�ڼW������м�{��kXǝ?'ڢ-0 �m�:m3�Oݗ���:�l�� j�&j����~55;u��G ����i���p���Zgi�;.R�q� �%1d�s�5��&�Yc�%�����}9.��Q���B}ϵ�+a�{���F̐ч,�%{��EdX�G�y�.�c��u�Y��DĞ��&�hҌ�!C\�Ơ�.��u����D��8�Ϟ�yt�~��2��q[ �O1���=|��Յ������6W%Bmg[%�[P#Ek��e��g�o���ZX�a���"�'�2�ρa��w�3,_}�հd�[F�Q��(�u[[�L����똂��4�]�w�XG�>�\/JD�Դ�>��������KYo�<v��n�1�ʰِ�Zu�ϖkb�j7�^�Z���Y��<����\>�%h�̼|�j�����ֳ�aR}N�8=.M{��������������������8(O�sZ���b��@F�ܜx���PX�i�fh�q=84��X e�Kf�YN�5��(+U0fTw�"�*��@�l!kk��Pk����˒�u{[��K`���W�GK/c�y������!V}��iS���@��_1�P�P�ȃ@���]3 �~d�1Kz��:��i�b���i��%A��55%�e�՗%�l�&��n��6'������1�<կ����0k3l�h�2������a,f��)�A���'��(�����d�P�0S�	@2�&�W�Ds�G�G��=ϼ]�	�64���PC�5ff�VF�w�hP�j��IF�esWڻ��� #�����Ѕ�r�`�FZRnA�n������={��U��ٹ�ݨ���l���bN'�p���Dр���硁�m��6�蹒�Ф�9Ѯ���-��ZS�L�>��������̢�����dH�L���&<b�����;�m�O����=�9fc��qazY�ڝ�U��f=��!���E(5oZ������q����Z��4���̀({���R\P�)�i!;�W��+Ò�|����d�Xf�e?�'��Ħ�)J-�2<���ԯ*-��7o��p���	�g�e��ݪ�6c�Yzy�<N����9�g2����m����VLFpc_�j��=�G1$ُ�Q_2������Gdt����n��4�"M�t�9)�����`B�y��2���邋���Ī�����pt��8�7�nҬ��u^�V�:Ob唌�C*�AE��q��w�:�F�m��g�l/CS�L�\�^o�n�{��gEs��FV.�ٰ$Cɬ۸������G{�Ȉ� #����_-^Fգ`�2��f;3����*ۑ�4�kf>��gj���d0re��2ŌF���s�/�y���ڙ�>D�h��X=ٞdVb]p�#�;�����k9]��_�KWD���#���in�.���	�}�˹��V��s�՗G;1[��]�W��c?��)�PB�f��nܸ!������9��b��zvF���9�u�چ�cV�d���H�Y���Yؗ�9����Ύhٷ�� 2�Yxy�8�e��&s�I���-̏��� ���24
���HC���y��n��W��>�3�dC=��P3�ގX�ia]Z���G���b���"��������� �xcIgVBd��Ź�K�B� �<��w ��,���0�aR�X����&�G,�3`V�`�.⼴���L�S�)�Yd�Y�t##�6<%h0�-�� ���1O�"i&����!b��c�աbBŤ��AK��L*!k��&�.S�	���c6�,�|��0O�g��W���V��,�pd
�)D��~���'2�:]9o�#��CY��aCOOW���0F��0�����<�(���������g��?���4,��=_���G�^r���\���D��ֶ��^yA�$�4ZJ;���`C<K���������췄e5��h��h�.�B�?Q?SZIZ+��14�5�.�5�s�b1��3����Pwd�N?n��x�hdt���lR�oO�K�f���5 �|�����D���ϭ�$1I|���p�9x�:z��fg����>.#{0����lG�<�='��׷�+�.����3=0q}50R��=����7���úچG�۷0�@�pYs��$nܑ��S��իRO��[�I��+ǩ/}�Ka��wH��ړ�X2|����x-�ú��zsU4a?�H�F�Ԣ��>��K��ܸ-�d6lv�6��hϖ�z��W���L�/�d@V������*��ZxΨM���=��Uh�p����T�,���y85$��u�͂q�C��q\Z3.Ƒ�]�YF�ꓶ}�6�Hj�������sa\ͺ�}��̓>>���O�]�Nr1����|*��~�ϜGf0/�7�=���gj9�5�C��p�=4YU�m�� �=�zw0��S��R�2�┓�/?%�·~�3ay�-O�^�:s;Ղ�L��]����Hbp��'���q;�5��V��Ϗ�7��a������x�Ȅ#��
�z���)�X$7���a��ߵ��\8`D拟��gq]�_�{=�_�1��|����3�����x��>���M��8�����mD�0Ҩ�I.��|_�z��ǹ���4��6�7��2)��l�>(2�	�����hoo-,Ƚ@L2	�H�B�^߳�t���vm�o;h�Jٶ+��7d��i^�c��g�yxxxxxxxxxxxxxxxxx��6�ђJ&-�4P� V|�
OA�C`���k������ 7��a␑%L�*�V��*d ������nYY`i���E=d�Yf�'�FK��L���P"CD3� ��r�i��3C2�����~d:�ds�8�ҋ�p&FxR��\֮_��5IL6��=��S�����!������	k��:3F�����3�,:`�ͺ>=;�Yh4�1����0V���D�
Y�6��xZ`r�̊ik=��<�>�kI��������������hI�ɟ�i��xR������a�����������|��W��f�yu F������z!�3+<�[r�+����ȏ�e	�<K����?��dl�Dn�G���>���2K޶�Q� fQn �.k3�b�Q�H^_5xt�����z �6�s)��+�t�G6O�����xa�̸D�v#s	0lI�J��-3���'��-ӳ����*�Y�q��S��9�C+fڹ�~��_��lMjyF�!]�R�c|ϰ��3�,M?�xq�d�Қ���e���/�dF����V��,�ЮC���:��"������*�_��[��~��	�������V�����mŭ�U̀.=�u�Gƭ�|� SC4�ƸDf��w�qHhf_�R���v��7�Mxʻ-j
�3_�{�&d*�HL�`7�f�ym���$�´��$&ᚿ$��I�}i�O����]�2����c��=Zf�Ks�>�g�!zb0���'{aE�X�4�\��HD.�uG0�<ڷ��2Rg|o֑Դ�x6ck��rМ7�R��>�_����s�'<:�+c�#�d�A�_i�g��nr`^�W�F3O��H�@��v�(�;#��^��0�猚�h&"�]�7#�e~� ��ۑ��/���!hߕ1]]��Dެޑy�_�t�c�%��X�zz�|����Y�������m�{C�O��12�� 2Ks&+�к����7;�p�:�Z|�o�����C���<��f;���O��_��N�7�	�q0�J2=q=�/����ثv��2v�5���3�E�NsDxF�������������������@Ak�(KbL�5�z� �� �'�D����j���' 1��`�;~&�*�n�
K�*���$'����t��E��������8`�9�����6%�J�Βi�+���k��V�ġ<A�DK0�l��e=g� ��b�ό���h�]�	M�i��**ZC�Z�����o��
���F���ʆC$���qF�����de���>&����0Q�q�Y���u����S�����\���O���@�S�&��_Y˗_�޿��o���}��O<zM�C�_����w��h屋��+`�
���| �������e�5�ҏ_��h����6�d^�ݪ`,ѓ��+О0ٲ��P�Lg������WYZ���=U50�����I�=a�\--I�S���>f�fV+2{5��Y�xv��ь�pQ��-hlL�9����6����12]M������2�&[=�v��(���֋�9���L1����h�f����ɦM�.E[8�&0�t=���\�m�P3����l��6K-#��������ΰ��.��χeeV�/z����v�FX*6'�����=d��_�G�Nm>�L�nm�ʒ�����w�t6�.�]0��9�o�v@W�C޿LJ�դY:O�!�8���yi�O��j�q�׽f��Vfڤ8jv]�3��8*3qRU����ߟ��僊��YOd������2?�4�3��-��5�C�� Bf�1�{�f���d�a]��R����/�?&�)���	���^��4�b�_�uj�_�xvd�+�l`}�u�a�f�12/jX��9����h�Bf���L��l���dlv3r��#�cYeKк{�՗��5d�����Z4�y0�`i#,�4���2���7Mq�U������%�捼~F6�f����ʹ�&����q�4�[-i���店�%[�+K�t�9ia���)��?s=5��
4'�]��P��ߗ�Ӳ׃��ນ�Ё���A{R��Z��!����>2��!��D��fG�s��=|�3)<�������������������� 2��dV��i��Ua̸X<��bl?,�h!�`��#/����a���j��R)���s��,�}��v�=���rQ�3dv\��2 �kH����i���5��>d
тM�<�:mh��m/���("���Ȩ	���0�=@`{F"��!!�r<해0L'\g�!����3[j{h[��y�1a3�e�PJG����|�Y�l���~�}Z{C�5��dlAC ���2K�
10�П�����eY�JKҏ
Ux��ц�������>��R�4���[[f���y�~��nj�?�	�[�R��H����d~�Y�2��?�r�����Vb�:4��v���ɘ��~���9��50��W�<��O�nmm�fR�����\��)�Y?2�+��̦EF��h���(�ј4�")=����1�nUh�m�98&��4����k���3O!��E�����իa���Ѕ���2���J �/ۓY͙��dU#sT��M��|�z��|�����7�7ò��k���M��,�S��m���C�la?/��ۿ[|_�g�>,Kx�:/��6n�e���9��׮��a�1�.��}���k�Q����G�V@��]��<%�2I���q�O*�G��~�a0���U���p8bY���i��4����qo�b��}J��s��ެ���|.��~��+۽bt�/����$��Xu0�2*�Jk�m�����4���DZ|��m�Y�����4̛�&�G���U�VS�!�YF���������ix��i�k?=6Yy�t�g�x�q�Y�+���ִ��R�k��Yu<2�ژ�P�����WZ�f~$�}lψ�4��H���L��)�W����7[�r���|��Þ24���gX����>{�x*m��3��Tk����mhFX2�kaV���WDs��l�m��y�n��i� ���#�ת��UYOp���|��p��>�G��Yo�̾[����Z���3�w����4�{�h�/��������������������8�����0Z[��0T��+�"K�&,�yX�+^���h���H #��H[�P����#+$����6-�5X��̲���������-�d���ϘozFh&�3��?�d$F�El7��m��{dn�bJ�m�i>����\;.1j��_�}2>�h�:4��S[,�?$��:�]�>��P2>������ӓ������-d��? c�5�,�&K����SG?����/|鹰����o�r�h��*�#�ne����Cٮ'׷�*����=,�x�d���?�ò4O/�s�d9z��a9;%����H}��؞+0u�����K>/l�A��0��O6,��aX=w]4 ���=���}�7���za:�?/�zv8���Q+�Ӗ�v�=
.2���l�h'j�QF�Y�@.�WS���dUC{nnJv�����D�+�=2�x]��k��Ɗ��w�՗��4:8��3G5fs(3�=�3���30��lw��Κ0'��qlԥ�[h��E����q�-j�f��ɘ��̰f���d;z�>��w�=�XXnn
��v�W���@�����M�&������R3fB{Q���?��0g?�SR������A[d:^�����ޕ)a��=t��G�^�_���F;�e�<��X��1;o���X2O�`�&)�Gf_��0��K����7�����V������7&NCe��0��u�a�i|�j��%.Ɨ���fǃ��v���q�/�ͺ캎�������컑6������3g�#K��2������`���c�������V�x�j�����4RS��#���q�ގ�X�5�mF���C��@�6e��Бp�NjA�o{S��� ��F+@�ߵ��'O��8~���Q�|,_�[�71/6�[Ӝ�@�a8��� ��{��5S빍r�,��D�Q��d4����z�E�+�7d����B�s�<`�a��H�r4t�6�O�e�����<ܞ�3�oj��S�oHH�_�h=�xF�������������������@d�ӆ}m���p�VJ�p K0-�%d�d�r��%0#f��fQ���z �ƶ0@Z��8��n4��Kq��r�`1�,�m0bf��;�"�)2����^�Z0F�:4=:;��jRL@Z�#"��G����7�gAiB���ž��<'��4�=d`�Xzƨ����U�����|�ڞ�f#c�MzgU_�Q3�5��ʲ��v��+��s�¤)��_t�v��ew��~�,�s�}`��C������oy⩰��_��aنcjI<dH�$?s59�O������I֢�y�����&��ci�I��O|�a��/<�+��0d6&�;�0�ь�}dî�Yv�����������@X~���y\��s�+��[7$�p�ɚ���F�ۭ��d]x��zh��w8�O���qpڃ&�xlO�;�*�(���j��_�-	����*]\r=K�7dX]Ȯ��z���
����I|h�uC1���\#�Z�C<WW/�T3By�˗��%5��;`�-/K�djx��Ǭ�;Ђ|���a���o��_���_9N�u�s��/�� ;��n���+���Q�<ٝ]�,��!~�ua����ˏ]K2�x����zѿ�x��sIf��E�FC�fB��ۧ��>���mf	p�@���� O-�5�i+��ƎUO2�9�,���@��@=>���hF�.�J�夘.�6F[MEJ��&eNz�7+&m��>W���Iǿ�ڜ�j���11.�/�)xV�s��n��E�jK&�Iz��zd\�8��aVO�'G�������@���8*�騈�|����vHu\�N3�|���f#3F�>^>g���~�������H��p_{��Y��z��mFQ뻁��⒬+0�]k;F���ƈ�?�y]��b�}g���z�nK�e��Bd�S��H�:��o�x�<4��)H�s���z�L7�Jغ#��4�E� D2�����P�V��=D�P#����� Y�9��I�����J�E���_->2"��1�d��3�<<<<<<<<<<<<<<<<<<� 
N͛�m�$#)��F�êx��d��Ẑq��u��_���8��Ua�lm	s�c���q�]� �E�a@f��Ģ[�f �/���8_�˗�IB�L�{f�!��}���>�w�!�i�iꌉ���hA�(K���s�x�T���9���@I�wAy8H(�gJgMU�3`v�ifϑ���X������N�iĲ_e�G��wS�kA#�݆e��!������c��$�ZF�?���Ͼ�sa�����?�?����O~>,���ÒڕMh�����/���������P���rS�J���fm�������n�Aӏew�"��p�h�,�r�u0�ţ����������ˏ~D��kk�}�}��Ű���0���0 �yg4�v�(C[�.���Jy������&�d�u۝���y^^OY�X�Mk� d$��Q#���H�EO1��,��8N���lo`n))Q���H�����ӣXE��=0Y����)=g-|߂G�Y�6�@��_��q�3Y�p=�s��+����O����[3,���}��?�����/�"̿K�.�e���M͇��A]�Gj��Յf	߇W�H�]�-�za~Ѫ�.�3/⺪�Ԃ��k�3~+�>41�W�=��*����6�5q�ٝ[�r�� �z�o|nA��|�'P��h0�m^��D���$͞�}z8S+-#�_�&�i����K:�S�OEh�{�2>��7�V�YgF7�m'�M7���^;�tC3�ƅ#}����U
��"�,��2��D~��'�|֮�\-��yw�N������~��iW?u�/��RL݁=�1�t}�a���F��zq����3Rv0�o4QO9N_���R[���5�W`���k�E�x���e%̫��yW�bG�� ��!�gsE0I1o���e�Jm���u\/5��>���yn^�uq��7^���<sqA滌`�u�^]D��lK�#�8��������d�ߋD�@úѐHF�P����.MI;س�d6��i�/�׌f�ɾ[��*"3��*��K&.#���4>*<����������������������4:�j5��.���jF,ϵ	Ȯ�4��K�{1'�֥s�u��@��0!��C�v�YZLv� �.�]�r��qfo���B�X��,�o�b�w�QV3��L�U$�a�o<̶'�������J}���g�Pg����2��0�NFY�Ml8n5�&����SA�q����h�AD-&�c?�ώ�̬����Ц[���7�ϗ��0�Ȫ4���E�<�h2����V}F�lȬBv�>6�g��X��S_�tX���0n~�/}X��?�W���/~1,��u��w�]���ާ~?,?��N ������S�^5\&̪{a^<1|�w�#�<-ϻ��f|�ߍ�Y��Ea@���@X~Ƿ{X�;�����^X��ٕ���1,L���5q�����:]�狞��BN�j��zx�g;���&Tfn�~F��Y���i���U;b{j��ٚlW�����M�?���Q���0L܂�j$��?���<_���7{Ȇ��e�|�j�"��]fKG;]C�����~M������AX�?/���2��^y�����\=��`ƭݒ盞G�-���8#Qfc[g�ݞ�U=�x���@#����E��{G���+��]z���49���5!f�o�uʼ�~ �V�aUk�^��v=��v��2g�KP�-0/^z'2.ޑH��J��%1��f�t���3��Ÿ��b�l�z��$L�]��x����}�>oiqT��IA�/�|V��y�0s��̤`�c=�qm�gd�9����/�ih"��Sۙ� mD*���{�6'� j -`Ǹ���K�i��\�,�D�6�~/p���*��Ǧ�RD�?�,��7����A=YQ)�<h��n�L��:+W�y����2?Z^�u5���[[_�>�����D���sд���F�@��[�PS��HH6��Da�0/��F��a�t�������
�@��Y��nw��`?�CyjBk���<��V*���\F��6�}��FN��Ⱦ�u�}�nK�W�I���%�yF�������������������Y@!��"%&��b.W�s�K:6�쳒��GECkqNb����[�};,��Ęm2粰���m��?jc�q�(Wa�����J���y0:�(���[F�/oǮdO�� 0;�Pi�s�63�چ�l�E��Zvq�Xr&��?�xD�	�4��FÏ����5�����x�	b}M�|������o���N���vt[ԬJ��f��}(�&bd���V�=X����������fm@㹳�jK�D�m
��'�'������=��갬|���:<p����������aY=/��\٪W�x��l��(�D��r� �^7�O��Sw��h4|��+W.���0�v���>�ԓr>���'�q�9}�y�,��&Od�MM��,�<}���C##�_���8����o�I$q�)j�1!�`�&UK��6ОR�{`�]{챰�Gvݞ��sJ-���r\��"����Z��dh6��j<r8.�p]�$���z���~/�*�O~�Sa����]�������4,�g���я��Y�w7_�~�l���s�̾&���L�������8���3�Qg��k���$��{�-�lE��^���%�/2���a���������}0�
`��z]�w�-�1K���˩�&@?��=wIZnN�܄�eM�����u=�2�bYq��q7�y��'=�>���@S����~��A�����I?��wڮ/�C�;*�/:_���ȉ�Z|����w���u��Ȋ-S�>��cD�Z/��|���^�<���hNRt~�0pԏߏ��\f�N����d��q�eܬ�:�}9fc�p|�Q/�ss�\9��y����|�ޒy05�mLm�h2�`�K�mG.�2[�N9��D�`��J��^{�歰�����L�"#Y��������Y�ݝ�^�g	D��2r6�ڲ>��g�~�y� ���xwV�s�̺"�������g��������������������qPЖ��Aa[.ɨYX�/�nw����X�w��kò�������Lڇ�����`��QŒ�SS�6��Udi-���OfB^�ۅ�yoW(d9��d��j����8�+F=�Ԉ�ź�/]�4�t��b�E�R1ah7��(ݯ}rN��]���>n��6� �^{|�3??��0�..ӄ��W�)���v�_�2��.��h����������`�D��EĐ$� *;T,����[����0��xR�mExtJ�U��z��G�d<�1i�2pM<T��&O/o3����Sg�KH&��S?�3��������!�d�=��h�����C��z��zUQU�CNy�N��!ϩ�y�p��!=����Y���A��v�Zf�K�o���0���`RS����|S����d/�Lg������ի������M�ې�6��������?�3?,?�я�%�}ud�=���h���I_����,5RT�Z�L(�y���ޣ^���Ӎ�`Z��ݽ��ԅyX�{y�s�r}�#�&5t�Q.A��_2���ngp\xv��j^��K�f���]
j
���0�q�j`v1W�j����K�I3��#0	�j���8\��q��&1SkY=���9.���Y'm?J[����<.�z�j��v��"Z��{]s��[����G�/����:��g3���W�)�5l���M;�&]w�I�����seݍ�?�Vl���D6���7O`�u[2���_�H���^?�;�Gu�5��s3`�e�K�l�N���u<F�D�{��ICf����]fvF"f���"�g̦���͐/�Iس�u�@\0Z�l��>�Ռ�r���zR���Ѓ�m���m�A��*@�.�� <*��[�3�<<<<<<<<<<<<<<<<<<� 
NO��<0����%d�=�K��-�6b6�a�bư����e�1�u0��`��Ń,�dB\z衰l���,.�b	�rI~���� �����0�����62@�10ZJFۃ���zЀ#��P���Q��tA��$�*��f�Šn'�]�,��x������@S��!V_����i%��:�93�ҏ�d�R�><�B������U�5@��ivU/�ZZA�4"�!(qح�~�=f�q�c�����O��O=��?�k�N�|�%a������a��O��w}�w��~N4�����a��	��0��I��P/����2����bيx8����˒��[��[��g��|���L�׮_˯�ׅ�ׄ�X�G�m�247�d~i�D|�e�R{�m�䃦�g�N�|��x�=�:���R��m�T&c��؈�+���P�I{��^�����D�_���a��9�����a���τ���
�����7��	�~��?,��{�U��KK�>�����[���S���ζ0��9���b�E0���Yu������ݦ��W��v�5��`�N��I>h�jf_=f5�v-��-C�<�f85�;�b>���ccR�ո̾I�uZ�`�u�<jv]&��<|��3i�\׸�̣⸞S���>���IL�Ӫ�w�0ק����/4�N��k\:��c��W���a�c�KM6	�NS�0�$��8���]/W�te�M�X�E���	�)�*b��0�Rv1�\���J�@;H�}hA�<-v0�h�`��m���X����6��6����R�����>eD�.���>j������)�C� �uȸ�X�[Z���TM�j[We�}=��e�����$�:��;;D��S�Q'APR��PË��g�>�y:<���������������������i�[�c����_	��ۢ����|L����?N � 3`��dݬS#��ih�T��Ӂ%�3D�0. K_�c�؏Y8���"��ښO����"������R@�#/��E�خ���5��0�2�R��]\CT#s,�J�_�l�y��E1tL�b��L�BCOʤL>�L��F߀1�����'�"����AQ6���_ߕ~QAv����5A!/�!��ch��Rې?�frQ�`��;jw�/;d�@��?��7���`W�������|�1a}��/��?���\_f�4����_������o
���o�tX~��χ���",��hȢ929���U���'E;��O��ţ�� �h0��]y����W�?�g�y��s�FV��/��׮>�_�_���� ��V̪J�����kԞРg�����܎߳ti���?��qڠX&�Ǖ�Ɋkg��,��1{�52��ʬY܎�5�p��>�.g{�]��XY^�&��G����w�oK?n����]�^~��G?�_�nɂ����}a�+���aIf��uh����^��������gUy<���8�<�q�� o��C����&�wf��Be����
���_�0�>����t�����h:����0��� �Ŵfϱ�!�V�G�I3e��<Z�7{x��3ĳ����!�Č:*��~]׸�\3�5N�:��Y8ip���|���Os���]G`���2H��m���b��sZ��u=���l1�<�t��븤�O:>��g>��+�o���[	cO�:����B~�d~�.a���9��X��!�uz����<�15����:�m�;�/S{���l6��M���Q�s0G�H/ο+��4���J8�ԃv�v�{��灑\<o��u���9�E.#�r&Rr�:��S4�`0g���qb�����a��W?8�3�ύ�@)xF�������������������@���x `Q���!h��>/���=��/����>uM��
0Hno���R8��� s������UV��>,�w�F�����ޛY��e��Ηｼ3+��/u���ZB �$�i`�	À�ݵ���]�Yf�cV�f��,ư�,�"�"$�@��V�Z�������>^�\,~��Q�{�+��Q����������.#�}'G�2��Z[���8KfHM�|��a��*��99��(3��4�y6�.Ҿ�҅�D ��U��^F���0��.�Ib�L�4A�԰#U��]а#c�g����L�Uj$�-�3ޏ���$2r�4Ë탮<<�H$#�
�^C1�4Z~������_���������SO=H#�q�3֗�����0D}�� ��c�L���|"Hz�� ��_�� ��_�9��O�gA;���w�m���0��eyN���z����z:H�տ��t�1S���9a8�����|[�;,��d�6�.�&�u��0�y�yF&+#0�(M�)��ۍ�R�h��qٞQ���K�ХU�����t2J0.��ZC�X�{�F�$sI��9�=	�qU�u֔�Yc�C�X�iA���*��`�Zv$���`���
C��r�����c�߅��s�	�0Z�73H��� ���� ��?�� =y�mA�������_Gy�{E�>���>-��h���L$�LH�!�~��"��ەa�%�D�ǁ1��]�Ot�]h��V�6.��,g�a׭]�	8��i�e�S3e[���{��Ű��:fV8WQ2�7���^w؝���.W=�e�E�&����;6���q}��_�{�i��s�4�v�U���]3�5\k:ʙTZw<M:]~�3��Q�Ŗ��Ԏl�;y��֠v~�`��q�O1���a�����?5.��WW��w`�	ץϻ
F Η�
F��s��k`�E�������>7.&�q1�i�-]�7\�e�1��}Y�U�c�̿�q$�&�ZK�V�,c��5X�S�t?�����J�2S�XJ�ӡ�W<F�m&�n_d,jt�2���!���2�<�������������������c c��"�����0\R�����{??���&.��U�� �� ��4�1�)-d�Ѝ�l��^�旙!WL2v8Ck4�P�r��=#�/5���	j��qk`������p�O�m-1���ן!�����b.h_U�e7L#�B匄4����ϸF2"��L��0?�v3��s������4���ڕ��
#�	'"(-bAmL�0��3F&ƅqV�A�9�?-U?dp�������9H�\��'���DPF��\� �H�lֲ����o����_�?�Q������U���*\n<$�����S�t�B�?!���[��p�S��sO���=".���D#mnO3S�@so���U[�oȄqU����}��?i��$�"��>Օ���kk�s�B̿�&�D[Z�$��\�Os�My�ܦ�]��]pF~,7ܭ�д;�j%!ѕ�@$���|֠)�kT���К�s�R��=8��M2ٮ�J�-�D�{6��|o��^g}%����*�'�!�qrJ"�g�ID���A0TwAk�]������0��ſ	����_������1���� �ٟ�� }�Qa���w H�_�� �7��/X�S*I}���MJ�Y0���IE�Z߿*Bn~�4ҧ_�f_���x3	��]�{p���ѕ�9<'U����$�'�#ʹ��ܾ[.��w��̋b�������]w�܀��<&_-e�!Qh��j-�`f��|ⶃ�vӌh�ׇ�?.F�븛��j7�،C��Ҍ�]�Ìc�Gy�;�"���G�j�4��8i=AT���]_�x2"�(�_\~Ǖ��9I�.w]g����0�X����^o<�7V�χ�ig���F��BI�������]*���������6@�˨��q}��4��l����M���Fe��
}�+2�ʪJU�c��%�8�����K��V�:��-�М߱���#j$��ޝ����T����O�}; �>���3��̧̘<|0H��$���KA��SO�؈0(��Џ�Yq���G�����5մ�Ư��)!&2e&�e[kp�~�^����x���N&�VN�V��Z��P3��"\u�hIE��i%�@��f���-z?l�ȇkb�5�mvT����1az�MH$be��=r_�_�v���e�1���	��$�Z��ZS�#%��>�!r�MɃS���f`? Z�¸I*� �!�\��fFi���b8ßT�CӲO�CK|N@�)��cG�������uL�?��?�U<7݈�L�
Sj~I�t�ǟ���n��W_}%H����C��q>9��{g�E㋮�+�r��Ľ���p�B���#4���=����y��U0��Rg�*��Ţ�_�6�K��$�Ζ�삛4#V�*�=����1hϑ���y]ܟ����\�\W̫���>y��K�al��f�/�oF�u̿1�h���`~�%�ߏ0_�n�G2�r]�Rۣ�H�q��ݥK�~(l��e0����MLL�<r���3�ȑ#A��o� �O��g��hh�ݻ�)��3�����*H�^\���fߏ�؏���Z��hQ2�Jw�$���R���� \�sѬ�}�10�P�޻I�&����<?oP����mA���.�S��YDd��-�F��̑�����ߩ繅iSCh�\.�����:�a���6%��q��q���
o���7
�}N�j���d���ŀ���-wf?�|/6v�����aY�_��Ӥ�{"b?���j�d%ۦ��˘��	G;vm�E�ff���z��'��o�B�K&�k�Ch��sX��~t�9 -�:W��~�V�)����pe0��ҥ���xt�-b�ɡ�lk�sj�g��(��i_M�/�?����e+n���U+$9n�aeH7Vt.�AH?#ͨ��Ԧ�"�z��>�ۮ9��������z�yf�c%C���>����>w�TR��K��"2�0��*���O�������~�{�4f�Ј0?����GI�M��ڌ>�,�L3fF��>庮��k���(s��ᅙ�50�V�2#=0"���>��Fjł�[��p-����h5�Y�P5Ɓ�F�p'� �[2< v&��s@�v�
��P�Xkߨ3t�r5�ӥ���[i����O"�~hK!ra\T���R�y�����$��]ZA<�4`��"�L>�C�Z[Sk�UF�XO�T�F��7ٯ�Hղ��/���l���w�s���}�w�Qa(���0��^�ҷ���A:}UT9h��NC�<-�qEͲ��r5�*5ٟ����,q]�}�ED�r�;���l�&�����+ܭ�4�Z5u%�
�]ayj�����O�5��X޳5��P��uK;�_��I�Hj�-��!h�������*"��d`��:6�om��$���g?��cc´;{�L���F�D��ox�79��/j�����f��a�.�����^G�����V�H=�W���ܳ��ܜ�;�������o������#�]���o��o�?�� =}Z��h�=�ЃA��c�K���,[��tY���p�@���7�4W������3
f]e��ܵ�F���9�m��ѭ,���s�v�G{^�:m����g����&�:��s0[�w>
�x'�O�˅N��Y�*g��hchݮr.�S܌\�S��Y֩�^��m�m��rq�o���F���Q���0���Ւ��ruz>�q�ٷY�����ƏQ0{<OS�Ǧ<m���w�6�~��3����,�!&�������]��[�c�K�g���BR=�ZM�*)��鑚���-��|���Ru��q)Wv>d�q���X��,��l!C�+s�g֠���U��^W:�c���qry��
�Y���
j$S�P��<4�9����2��,��RL��Wj�J�岌�^yYƇ��?se��l_��q\�B�FG��
�(7�П5n��faכT�#+2��JMn+�i� L���VڍDdjO=�7@��Qpͻ�՚��>�����&��q1�&F@���#2C{�0�^�� }��SA:�(Rǎ���l�`�xen.��FP�HS�emugZ,�=���"*�i��\3�k	�9��a�����6֬�����4�sa�H3՘8c1CSf���MD%��4o:�R��������`NQ��hG�8��N["��?��*��%۴��hP3!��c�z�	�����6��20�g�yT-Kd$��S�nd2%Q��4\O�v{�N����b�q���ljZ��|��LV2�~�{�4�%���n�s�X@�g��L>2ɨ�GM�nDp���S�0�='��A���p`��12���T�)׿��i����F�%�TF~%0�x<5	�.����"ň5������p��&#Xt�5�*H�lcİ���\W�%[˃�����f}��֠���H\
��.���+��01q�(�<ץ���nL���wi7��d��d���0�#�</�tu�k[����s�=�CC��#�|8H�|S������|��E��A:99!��l�ˇ�S��	ѪeĒ�˸��z�2��6I�O�+�v�8�<�0��J{��i<�)0�R�n���C���zR.����`"Ǧ���Z���?�|{�K�=�sXo�gʯ�-w�1��N�V7ZKm�I�[͸�T�o��U]̥d\��#?WyR[����j�uz_\۝��U�w,�6�-ڰ���=n>�o���7�`�:��2tUu���9 ��y���NI0�3��Ԭ�24��䂳�;�n-��L�(W�d2жN�Z�dT5q��?�~BR���mf.���ICD�������`?;��|������a���fs8��jg�?J&YeF����Bj�s���g�c�L��XI2��Nd�q?���5�������?j�s��_\a��)�ZZ����Ç�����>w\��aVVqY���f���GMnΫT��ؖ�S�o���t��M�W���IF WqE�W:e3�\@��yQ$�G�����������������������Ș�t�9��3Ѐ�Z3�������w�[�NO^���A��&�l�<\B�p0�{tm�P=sj"��23���N2���3�����*�xg�� iS������%��s������-�|���p��ƍ4��Ռ���u�8�\c�FJS�pƟ������$6��c���o4-�˓jg�d�BG0��lN"�z{�Mԝ��$���y��T��H�1��v�_w�DF��5�V�����ӫ�4����+��������ŋ�ZJ��"?�ny�f��D'j6�F�<j���.I�A��;�w�����)�+2ƴ��%�}���P���KX�g�!��رcAJf!#O<��R_t�mW�$�-�v������%�;4(̽���Rj�:�ac�0���zSd
�A	& #|��r����UDήB�q���e��>�-�z��]c���(m��!���=<�
�/�rP���O杉�!����3O?�{���G�H�>��cA:9)�}`f~�_���	ҷ�>�w�qW��8qk����KAz��� =��hWy�����󼲴�t�����5~�WLj�d�'���)���^Sn����M�6P�3.��f3ܢ��Zr�T�W+������N�Q��cQL3��B��Sq�7�������1�#4).�0.n:�8.������?�j-A���2��Ԡ�����-m=�iS�!�(��
�������q������%!:lf.&1���.�R��%�8L������`��̯�V ��,��d
���LIw��r�q29���
H��opYiD������g+��4I*c���R��q�$4�W�����/�]X9���3���
{��Sb^���H��﷎�]��*��4��iX�
��/�R�� ���?'�a���L�7���
t
ɂݿM�~d��LXi���]���Vx�r�፰Ůu?��{Ҽ?4��+����dcχ�]��}; f�/*b��s*3��!_����	#���}��,�b�=/�}�2�z�	a6�+L�}�ȟ3嘙�Li���j�S��O��7��?�^��GF#��8�^�uv���̢>
R΁�q��P+��p<���`�1뚠�ɗ�pf��5�F�`���Ү:%��E�3�nO�kf�q_��yD����<�����*�U��ŽI�.��9~ua�ۮN	���Aaʮ,J�h�}c��l�}BFd����#<MDܞy��r�.�$MO�6�>�YD�N�~+H��f��.Ѫ[Cn������F]��X�0��vD�	�'��R/��3�7;3�r�y1c������� ��������,2�.]���Kyn=q�J��կ�sg����|D�c�H���~8H�����3R����������a�1�L-AF������N-2�^ed�M�'���o3#���-z��c}�
t�*X�����J�A^G�EF�M{����X��-�=О�ɟ�� ��_�wA:��������R2���'?��A��o�ٳg���g�FF�����s�c5�-��`���z"C��g�� �O�/	s�����0N螟���as;:����yLh�~C�:���r�\/���f�F3�6����l7บs��S��~�λU��Q�#Wک�f�)��db���"�^�g��)v~�[���R��ߚ-Z�-�8��uR����,4��h�b�E�}I]!��í����h���]�[·�P���y��\�gV�j6+~�Kr^��e�[�G�j��uJ�OMM	�����z���t����p7]�����������F��Kc�G��"���Ϻ.��>�so���0�Σ���o�� ���ih��M���Y�K0��R���oiIV�U*м.�>����P�Q���/��a��q�PS�o�����T�_�,�U,�q�+B��g�yxxxxxxxxxxxxxxxxx� d\ ��'+5[*W�n�v�U"�08$3�_��G�tfJ�:�w��w�~O��
S"�|kX�Ě�l3�XC݄���Ũ����5�C�mFC�[�3Mq��L������{�I����f�ʧ��X�,_Ci�5�K�fEH7��\3��T\{`5S�2s.i���ܧ�ʅ*�0%�w[�C3�x?�M_�h�yS�4I�5u�����kp]���"d�!�s�� =z�`���\Z[�|�JyI����B��}����y0��\]�w��Y�$�v�#A:55�rH>'Oؑ�����=f"#lk�7��E��6 ���HƖv�*#bD�&F��?#d�`���:E�^ehX��Hd�0�q�	ڽG���>��3#`dp�c,�ܩN��G���/�`]{����921�"����AFߕ+�ȜVZ��2��,�"p���Em
2Lɨ3��a�̺�?�o��R,��?�H&5���d49*���Ŷ�q�e�,"wo��w��� ݿO���L��Y�q}T�kw�-�12j���;�3H_}�� ݷo_�V�jfܣ�}�M��� �/��o�9#���ǈ����gj�I�\�\˦�g�Ը�{4&n/�8��_'�:��lE䳂�CøG�m�&�V����f3۶+Sn��fݷ�b�E����^�F��:>.��SD�sT���(����Q7g��SZ{+�%7̨��7˅��jM>��l�N����mΌ�ͥ����;�ظb�h�����
�:�?}H�MM�(�Q��0�{'�{x���8g>����hn���jj�esR�=p���Kǯ����o�֦�n�)�^�Q@?�
���@L�+~8���Ѩ�8��%�q|A�d�Z�u������g����xk��
X���]921���yn�㗥?[���F=���z�ե�L���h�c~*��A��سS��1��F��.��o����>�z�A�͈�'��C�%�Mk�N�|=�������������������c �*`�Yo٦[lCfbW��Z��߳Y�)�a���aY�=�.�����>HR4��e���;���cA�B�!�f9d�zk�M(�
�Ȯ&���*���,7#Z��03۴Mz�H�K���Q.�AӋ�|u宫��s����NAT�Q3A��=%�5�q.wڸPN���3�ޡ�l��vX,�}_����� i�&�^3���I_�s�>���I�Q<F)�$QBd�����#5���0�j���Ѐh�"r���1a��5���oi7�@w�).�_��/�~�h8r�P��yC�Fu��^��얡�@����o����DfS2|֌6����S-R@��P���U��[W��l,g�D2o�M���W^	R2�Ȭ������ňR�s����㾓1V���E���!RFw_2��f���1�HU:�>�s�С ]�����O�ܲ�9r��6�RO����1�*i�E̻H�"#���/G��Zdı�`4�<�<��Ii'_��?��?�� ��#�l��~���C�产����|I4{��ˀ�z���)}`�R3q}3h7=�����_�����G�������r�@�x �Gj����]��Z�M��6Ӫ>�Ω�]܈��`QH����/f��ȕ۷�(����i>���Z�V���S�W��t�N��{�����;=�F���|�"��s���̾p�X��l&ߖCU���8A�gM�5.0��$��(���܏�H�-��r����e���
���Nr�Q�w6�J&���Q#E���{+�:j��S�J&�K[��d�w�D��Qo�=��ܩ�i�^]i9�����P���(������E�we^�-���*�k����e\@->���;��f�d��~$���
V�P��,4DZE;bz�(��Ǌ�h���"��@YX��ร�!뫂�N�f����.��}���<v��U��Y��"丑�s��� +�VV�p~9]W7����_����r+��5�8l��i�gQ��;��1.�k�ڿb�i����H�|�G�/xF�����������������������4gI��w�̐3� �k5ΰ�i:�5͘��dd&��w���{��'���S�Jx��Az��6�=&�*j�[�M6��@�j3q8��t�zp��&]Q�� ��]4Ӆ��2\��]q��=]o�L>3SKƘC#`ہ�U?w������D��TFj�q;��nՌ�p/��6�f&%b�lP�\X�Y[��f�E�Zs9�DBs̴z�h�-/J��5y.`����H�DrJݢ�Н�R�$�!F���\^��F7��ɗ̿�9a"�}�)WI�D�{��p|BE��b�*$A��d=����F�?"���M��D�A��+ݛ4�m��<������U�Kʹ��������Iq]= M���z��*���-�����Qp̹5\o?4�!g���=+��F#�.�ߣ���&!���clnn�:>���0�*�v�.M2�x=�n����f��4Z�Y2Cmm�WFd���m�3#�d�����zᅗ��;�M�;/���a|�΂�����'����_םs����ИݳG����0	?&��;?/��-�7� 3"|��� ���v���/5c
��}Ӛ47Y�mj#�r5Q���^��=|��D1�\L�(��F��:e����YZ�[�\��F���}�)�46�ρ���Z�z�|Z�f����$���PjZ�kg#Q��o��D��Z�J�2���h����m0�_�{�YYc��63���p�A�����5�����nol�d�5��N�������Ei�</d^��Ƭ�C��r.���dk������Zz{�Jn�r5H9�+�d<F����W֤�q�Vb����&��#+���פ�_�~5ƹ����#��� ݽ[�e�Of��~���^���5O����Ʈa<Lw��{$�м~σ)Wh-.����8V���|n������A:3=����W�K>2�����yd��f}H�D����H�8~��e"�H�u�|hW�͆g�yxxxxxxxxxxxxxxxxx� ��>gDK�1ҥ�3��=��LR3�GPc�n�2�z�{d&� 4�N�z3H/`yjR\/>�\��qV��{L1�����#��3m$�^�EuI��5�]%��-�1�/Bs0Ow^�$�L>F j�.�����V��o��U� JZ�s(�\3y��������d��l�|��#<d�"�B�DL�e�<��J�R�HQҸ�[F,�h�ղ����_��dR���U�����&�ʊDHz�d��3�j� B�����7��ҙ�{�{�Rj�1v`�Dd&� �R��-Ê��5)w��#"�V�.�R�%0��<�"r���F��$����~�s�+n741��#��le��j���r���������� }��tzZ�g_��W��2Vh��</�I���F��C&�Kf��t��Z'<�4߮NH�q.V�)G�C��b,hF �خ|W�tnt�u1L�ި=���q�D����wg=�Ř���1q���"�|.]�hOm�R��G��AMJ��%h��G�y�E��V
���uh��;w^�_�ߣ4^l+e9�-�BV�AM���\��cA���1�(\�>㺻Iخ����z����f�mn�lT9��wA\�[�q����}Zo��U�zq�f�s�KM.�gC�~�����^i�'���?$���Yy��W�p��t0�Z4����7�6V.�&;9>��|���W����H�d�7mf!B&�Ok���V���^�/��ײҋ�5�`��N=_���˰���N�Ј�^�mp��%0���6W2��E��2%�O�^��Z���9�]�R�X������}{e%	�~�������}8������װ�&�q%�߼�2V�����8����P;������8N~�kJ����`X��|n�ss2^��^/���
=2n(���x#��K}��1����`����E�0#%��������l}�l�w�3�<<<<<<<<<<<<<<<<<<v 2�R��� ����d�.52�L�G*��<v�����C�t��� ]��g���)ٞ�f���04�/��-]H3d,���j9uu�Lx7\T{��ĵ��pg���Ԑ�����ŰI�$0�t�UL����>l�@�a�%��y�
�4�B�������>�l\�o�OR���ih����5�3����ZE��d��#{p��+�|�oyy�\f�+��:yH"/w�����|�Y����r>h�%ў�4������vUŬ�{��/S����A��C����"8+e9xdv��Fʹ9�PQs��V�%�Zo,� \�WW$E��̬�F9�U��x���W@�dZ�Ck�C�� ��,A�#Ld��ݼ��h����f���j7�Uh^��-�RQ��"\_�E�^�ȭ�I���s��=�q�(�@�D�VL���e���\}=����.�Sp��w�� ������Q�x��KmFj52F,	^�io�~2��~-���4��sp.���w�
�oɈ��􀉌h��sҾ�M���Qy�]w����gF-j,��߾=q��g�4H�y&fj��8�;�[��)��DA3�]��8���,7ӛ��{�w�L3�:e�m������j������Ԍ�����4]�m�j��\��LFV݌+���l�˶js�d�6Xw���e��v@��{П�JkX������[ܕ��\��p�N�韒~�R�.�*�l�W\��61��5k?���������T3�R)�l�@l�
T��Z�Zyȗ�M�a�ֺ��W q��4,�U���W�S�a�e4���rP��N���Ǌ-����c?����Y��4��}��� �qOWV�e��Ǿ��K~'íQĊ��\��
��ؖ����W�|\��Z�\���s�)W>�B���Q�V3ؿQ��/�K;*`'_��,Vb��lG�mN���u�>3I��bnZ�~o+o�iѴ��Zӱ�c��Z��~U=�������������������c�9���i7^=�XI� �<��$I�)G�\2�KWIfV���Ñ[�4|�32�;7%i�\#���/�|P�0Hz�8)��"�.�A�Hr�f*j&5��
}2�8���;%��en2Z�iv�[z�=am7U0��W ө��U�1b�g�^'����0��F���U��\4k�\� ^�:���i?\V�$�۵������2�%V slۼ?|0����̇L.�VS���)Cہ�Y0�4�4;#�D2��d#cpm�va���f(����1{�������O)]���B��ȗD�Fw���n��[*H=��E�|/Ck���t�F� �#A��r&�[2A��75�x2�Z�
�ׅr,�5��H2��#ӯE��D㲜��48$6Ծ�� ۩9�m0�POlG��.��K�E�v����t~l�+���A��O�f�TFl�^_~Y\~�y�� ���;p�e��_{�� %���yy�g��QHd-�`l����4m��S���m�dӸ�L�U7[��F]�F]n���GD1(��dIs�pi��t��_��7L��c��7�o5&_��OX�5{H���V2t	����f�m�x� Iנ%m��!H����70~�����T�nU,'��e��h�{x�\��?�����T3�S��gV��y #.a��9i�����v�}�
�(m>S^�_�u%T*��V_��<p_�<A��]��.�<B"�qYC�o�k�/K���q�n�@Ċ�9jk�}��e�{s�����|W��0ޘ�x���8"������?yUVҼ��x!P�ی'
t�-�|��2��2������<�'&�</��r�r��kl��Y69��_��b�'��"��2�g�.J�+�,�l-t�͗��b�%u�5��b&��������Q�!1��>��L�E�b��i3����3���Hc�;M�h��k�eyZG���Uy��H���	5̔+�YaD��\C�ૣ\t3�7m2��fUTĭ%��P��aA�t7[[Q�=��5�4G��4��"����n��H�Y�fJ-�Wg_	�?���O|�A�E��̰Z�vSZ��[WN"M�pD�ȠZZ�5:�)�Ք��X㚭\5���c��(S2i"���$�`�1����t�5�`�(�yV�@L+�����������@޿_"W����g�	R2�*��{��0�zP�y|�� ]��Y_�Ј�pA\]�VE�Q��_�������0��aY���2?���|d��FDe�ڈ<�����Ԟc��\����c��go"ɸ��<��x�x�,4�=:*"㈄R��R���Q�ÌT��-������~h@�[�)0@��F��5��X���������烔�Ϗ|�#A��/}1Ho���U|p��>�(�)�@�]�c���v��L����ڪ�UQn���\�ʧSt��u=;M�m��ͪ��j��tm��"n��uc��|n���bb~��EKK!d���O�?LP+N}��BSY�Ǖ�*��Uٟ+Z��S[:����M5~��|���������7��I�iw�Lg�M�hg��'Rf	���q�����g]�:�~]
�����R�/���/�`x���.9_6�W�?��d�4��kqI��i\~���_72"��~̏Lc��Ҽ�i=6&�:2����䩯?�d ���~짇����y���_�Z�r��A�Z�M��Ą��^|�� �z^�>�����S�����rY��+������+��v	�s����q^�Z���|V�K'�v�\��u���������!����wq�}; f�/.)j~QG������H���@�L*#��$��C�J�*�k��	j��c��A`����G&���cǸ2"rB��aD$.�O����M��ݬ�wJ8�b����p���I$�ąL�PG�7zF{m?#Mtb� m�4"LS	�o�a�Yt��wXgy���qv�Oƪ�����, 3W�ѕ�~R1uG�0���π	̈�ꪭ���.���h�AK�0����|d�D��`$2⥯��4�����>Hw�Mj�l�}��q���p~��׬r�I7��Ih�Y���'<jԱ��={�%/���`=���kV��N2��#Ƞd�0RM�|���y��v`�d�q?2y|�s��5$���f���f�������I�65E����������`ܱ=h�%5
�c�@DDy����&PA2f _�����{��ҥKV��M-f�=�z"E���c�mwͰ�2x40.�(.�'��:� �bB�lMŭ�V1�֫�~�N��;幋���u����j���L��q�;���5��{V��R�]kM��r�M&ڟ_k�S{����2+��������짇�d�9��:�ACw�?��h�o�>t�1;��N߃�Y�}\���?__�O�{���?�����_�����i����:�i#c��v�Ξna�5֤|s`�uAk�� �8j
����O�vw��S3��|�M�ڛ����Ǻj����A���(�PZ��a?�+�;������I��'&�x�� }���Q~h�sEV��J�I�MMK>K`:f��7,��b��c�\oo����F_ZikR������R�ݠ�����>3V���Y��h��Ux�:����������������������}-�<t�5n��;d3�LSj��~��&�MQQ�`�rp��a�ٚR!�IG`V��2��R(�`�$q}D�l5t�7[�a����yh�Qa1+̙�y����ٺ(?�ӵ�Hb���n@0��J��0�+ZcŴD$n��� =��H�Ρ��g��f���G&�\N�i"#���<�L�l��-y�w�U��s]c��lƭ��_��"rҋ���DE����n��AS�׮@�L9��-�2������3�C���eD��;q�-8N���GF���5�ԃ�z�_����Օ���]tfy���bm3�F�"#|溌��ܟ�[�p�_�A�XCi#2j��^�Rk�h�|�\d�Z��Z�Z[c��"�����S��L>j����>��3q�*�'�� m?FGw�5�uR3ωܗ1���^خx�Y�sp�e;�A�R�}�|��I�s2�湗v�W%~�?�� }�� G$���x���@,�HD4�ɛ���(�o�#J�O�j��c�l���	�Ӵ�Z��֩�"�����7K#n�����s=?�y�j��<���f1n��^�qJ��\N������I5�.����9�R�5��JkO#�x�Y?��3��p�Ef�ߛ�*ҭm?�/�`F|����tqk�	'ד�sE����&�9����
�������+r�������[�{���{�x�]�f!�wO}�� �|�r�b�֍���w�h}/b�z2�d�{s�q>���5�g9l��W��B��ؓWǃ�M0����Tƞ���uʸւ�7)L��I��5](��khL����a��ze\�qD6C-�,�%�&�f�eP�d2��iVz��+h�ϔo�	�Z��c�>�����������������������E[��9�V�02ψ���+� 3#O�����>�F�5�P3��~f)��Zk,6�/���b�5���nV�d{�_o��ܖ�HbġR_��#Z#֛���U�s f_S�%h9$ք�S����0zJ9�T,.������hI����i���-W'������`���h+��X�JF��� "D�S6�E0�Ȑ#���_�����ߞ={��]�l�	ňԑÇ��ɯ=Hs�Rj���AWY��.���{(��u�y�`��'E##t��VF"L�S6�0d���iA&�~���r�<����b�����V)�~te��+��*6�!d��{��e3 �IG�Z�:�n[�>_.�����ѣ�$}�r���Ña�Q#����݆��,�����]B��Z{tcd�夶#���U��{d��'�K�Z/2O�.�'�.ԆɎ��m��K�������]`��1������
��d�������y���=��|Z�P�9h^��zƧ�Q.T��$�̾�����
���Ao��}��׌��=����]�^�b��ֈ�Zz���Fi�i�ӞO�v�F|��wV�s�J�������b�5c�Oo����M����j��0Ÿ@��k�z�������N(���m�mC�����R��F�,���W{��>��-�E�����u�2Q��[Z��3Y)l�韥1~�^��K�&����b�4�'��[NȊ������c?��9a��c���6��f�3lԘ����1f^Fi��{e����Ê�"V���"�/H��8�_\�2�ޛo�
�K���x��� -/K�oH����
��Q����/!?���.hx������.�%\wnĹ<�ߺ����x5:Sm�CWf�>�3��|7��}; �O�u(�ƙ�p����N������".�����Pg/��*�3_M�sR;��s &��u��N�,�7r��{�H9�����SCi��0v{o��s��8MZ�==�A@	2�RH�aH�k�}��0�����H��~��A����o���GPZ�x|\?d�Q��i"-><��pm�A�b(��ý�L��2O��f`����q�.0����7P>٦��>����Fm�0�Ȉ2`�Q�"o�v���xК}<�7�~�:?5�zz$RT.����$�ԔjJ�>m3�����9���(�ע�G2���O<�K�<v�X��~�0�^z�� e; �L�3p�%���O�=�&�z��<'�KܝY�o�m�Zx� dDp�����������Wjj�B�L�����+`���+LչyɗZ���i��:�i�.�oE0�x�=��u���RҜ_�ovV4R�\��a�D`�0��s��\�~���yd�J�ff�������qi7�o��������R?�0��$p�6����f}k<�d<��NGS�����	����"F��<�tf_\l�����Q����b���[o9�{���t��ɜ��N�s� ���3-u~Q�w�z�lƥ���0ĭ_}���!/�ySJ��h7�|����V�+�6�56[�ϙ�/]w�:m����M�>��ɺ����H�[�l�������d�k�,�v7V��U�}>�'��W^�~�K/��7屢��y���1�uQ۝�Tja�j���.ż���q�8��@	Z�kk+(���>hSk|~QV~�>}:Hg��G��*�|#��C�/��� �|���s9�_̻ӕ���)R{K�G�1���q��.9�mn���}; �uπw��w��c��*8C����v���x�f��w�����o�l��c{�`:�oq�Jڻ�?k��9�eh)(f���ף"������!{?Fڸ��i���]���9{U��}�T �5��H�IU��ܔDF�� �;��O������#���ͧŵ����K�����J��.CȸM8��Ct��ơ�|S2M�\/���ٗB$޸p���0�����4��#ptY�Bd�ZfiD���F-8j��w�(���	��m��p���WX��^�K,5�X�+#i�VG�[�D�d�Qh[LM
C.eڭ�����1��RQ�[^�� \��:;�[��V$�.M:��4������kt�G��*�E�$�����p�F#�g�ƈ�2�S�<�f�n2lr��!a��5��=]�� ��lW�2�'�Do�0	gЎ��� }����1�W���;��<����[����K�0<t�P�΃IZAD���C����x�B���`�{p��S��~�'��e��ˏ	��\���m�x���S4�� ���ޤ�T�P�G����`���(^w�o���nf_��N��FtQp.����f�mWf��)�]z��$��Ø�n���ݰ7����/2}���ZQ�r��o-K�T��t��+�\�������|��!�.���\�V܏�s�qd6��q�_���糑$�W3���r�4���OH~C���_/���󢽝��k+G�� ͺ_z�-��J�c�` ��K�2���JJ�A͕G�rܔ@9#��{oo��s�!�����K�+��>sF�|�^{M�)�]Y��g���û������������	�͠���1~��"�|�'u{2�k�0w����������?�>WQ�k�x��>���O�]?PTH�$q#��xF.�� � ��S��\7��;ū�ס=î����:��_�@uU����jr��AS�c��v$��i��7��Z�b��m2�]��u�JgiZ�I�����%������ۏ��i?b��9xL"��qh�����W^	�o<+�r����#i��e���Gܹ��C�Yg$G��R�h�A�,	Z]�d�~+�g�tǕzF@�hO0����S��3�D+@[�L<F�q��D�j���by�`����-����;E�nnV�X=(Lʹ9��?���?#>t���]b�8�wjrʺ^2뺺�z��z;x@��ի¸+�I�qr���!8l�_/4 y�$ʑ�S�f$��j����##�Zr�� �.��h�*���-�1F�~/����QE��&�FK���vI�v��I2P{�Ү����v ���R��{�7H��uON�%��yJ��["�Y�'�2Y�
���O3��""�U��4���q�����OI~e0H�溻P/�{��j�^g�2$� ��O�43��A)_�(�(�]��oq�?-�j!U��{$�B3��21�)�n��[��:_o�Z�dm26�q���빽�L�hm6A�u��ǅ��n�22o�w�R��W�
�]�P�:��0��d�4���ʠ��&�_ҡ�ƕ0��W?���gn�w՞4���L?0�Z�M{�����u��ƩvJf^�%�~�݀��_c�S�Y����
�;�*�a����k�K�Js]�cf �9�wf��gt��f��8j�u��}�_��)W�d22nɃ)73-����v�n�e��z�,5����Ǳ0�X���1���'je�v���? ぉ	�h�"��2Ɨ�.�u<��7%0��`T�e<������R?��d�RO�� L��3hu0��74(���xL1@��2V�q�^�Y��7�09Sd�u(����9���}; 7n��Ql�V�.�Z����^�'��Ei�m���{$�/�̫3���5��|"}-�*�:#�-�ٞa��f���wiF��Z#�v����Y�f�F`[�Oׇ
����P[̹L�0Y���S�{Ѿ#�����Eɇ�
\�V��Y��"4�(Z�{m�.h�MH���Qqݝ�@�>9%̣�9�Ç�p^-C[��iТ`�m����3�~O�����N`v�IE��$�K�*"n�pA]���TY�G��h[�=�%2 ����FF���p�-bje�����ɓR�_|I��{�q��[�V�v�:�j�i��̹˗%2��{���>�X��ݵ��_�f 54SnA�ueD�^��\�7���۴�sd<���w[�\�tٺN>�5������W�����k-���w�%��/%��̌܇y\�q�CD��nj�����
�A2���4�)����o	̿�G�!G���q��RÑngdp��9f#��G�����%�˗��� �����*���[�v�3G0?��z"H��D��kR����e��b7���n�z����g��b������������:������si�|/���_I�/S�W�ݸ���V�ss�1�\3�6��b��e���@�j_��N��2rCw��m���h��|6�%�fi�,��������0��[+;��\�k�f�2_j<��I�8~u����$/�����f�����+�x~��2Ò-nOQ�q�i�27$HL7Ō�p���}&BB�`��KF�jl_�Үfl��4�]t�Ma`Z��ʌ4��I�Ǘ��� ��jE�3�W���K����g��Ӣa�jX�K�mpH}lGd��NI��Z�\�C���-���L��N����|F���7 �L����x+vv�M������%G~�)�K���}(�H9��qO
ҽ���G��bIΗÊ���(w+b��VL&_Ji*�����fc�t��3�9��J���(%�����z.M	�s��w	���1_=�������������������c �~&Y<��Ik�u:� �Q��5c�����V̮�l�3������4c'�ps��~�Cm�(�G�*���T�E_��rԈ2�*�����ɤ��Z�-4����s�%�3� �j�Q��Qټ��m��u��;��.h������hA�a\Zf���	��#A��$��p{���Dr�\������m��*�F�fđ!F�:F�
`��劑�a���P댌,2�9�#S�`�Q�o�(���f�u)7#^԰�n�D��)��.\��dֵ���2�׃=�d�M���vKd�ʸh]��x.\���Z�a���*�uSK����t�"ÑZs���5�L7j���s����ƛ�u3�N&�Ԕ�2?ɤ{��ۨ)/�	�|ɀ+�=�H����0��.�̷�P�T��<\�q�)�y�~a2>��C��S��g�H���~臂��g�E��V~�Ғ��͐BA�khX����������R����)��1R�1��=F&]ך��G_-ή^9�oL��fLǢ0�|�ˋ8?�H�EC(��y0eɠ�Q�[�=%���#����������F[K���F����N����HZ732����o�..6�y�^8��[4^�(:�/�P�g���F�{�eeT���;�~���hʙ��{x6���S���%'3�q=M���f����Z���idl�qQE^K����[�~6ǣ���q@���fL�IMF���V���C��>��V2���ʫjJ��s+2�K���-��i��B{���!�뻱"%��p\�rs�O>/�gj.sE�����_䊧��� A��㛕U���{�oJ�����?w��k+u)G�ӡ���`c�dܳ̾�!o�RN2��R+��05����
��S��*��a4����I�`��6ϫ���r�2��۴�]ҵT���g�yxxxxxxxxxxxxxxxxx� d�<�k��7�F4�A[�&�ftCI�x�D�|��:y�߷I@���#K��fG�<�����m���ܐYj��U�$Y��R}�/��]�zF$2QY��Iyf���n�)k�I	27��j��&�F����_�|�� �����Wz1H����D���+V�%$C��"�c��t�v3f�iL�}�ۃ��99?5��*d�	c����02��J���Ek���W^}5Hg�|#Í� ����������V9Y�0���f��C�����&�/FʨA�
�Z������0��0��1G���"#s���u=����/X�1R�����׫2�;�Fj%�>���
�����8��F�_>�t!���]�d�p���{p��)�s�.�3�JSen�d8��B=H=���i��GP�d>�w�{�(���qu�\�'�xQ��~[�Sfm߰<��V��%mG:�D�i[��ڂ+p5N�~����z*/�n��
]���޳e��|a{z[��b��h�`\�ElO�]����t���nn���nn���C�IG�� �-����ǶF\wcͤ	t6���\�=s"�{��ÓVy�|'�.�+\�`���hM�IF&�#�����������&Q���V�b���/5�)���A��N��-�0���k�Z}!���ʆ���Rlg-�>�H�K?6�-�޼�{���W�~cb+T�R�����\vǆ��6�-�;v�@��ݽϺNjw���N��j�^��~<����\�+b�?欬�y㔌cΞ�qɥq_��K{uM����N�<.�~��w�J��Aٯ -�<ƭ\�D=f1>�x��Wӏ����݉���\?5�RM�l�u7m>����ߥ�ɧ�}�́g�yxxxxxxxxxxxxxxxxx� �L���F#�N7���oz$�����N��}"���@1��u��]�+W��QF�<9g�q<#(d�HX�}�6[:cD�._��R�DV��ݴK�z�vo�D(��H�&m��a�0X����{աYWco�_�d5��fRO��������� ݷO��΁�����{�c¨+/I��7D���l'O���ߒHN�ϨH���"+Ý�Z}d����1�79�4���2�8�۫��;�S��Q3��{W'D�j,W_��gF|��2�~to���{�����3m�v��
Ud��r�� %�oy���C=H>d���	��Vt����o�E�^]r��Ldyo�;+����:}Z"u��.�Ggff��ujw�[o��+L5>�,'�������0G2㨱1�����0���_���sY���V�����5�rB����.���|��S�u�ȏ�H�>���A�H��/����ԧ���菬���k>/�S��=��?��?���~E�'ʹ�<�w��7bZ'�톦b�_�o�-�.;bk�@ԇ�P��3n��x�����w�F#�a��e�������4�[��d$(�����*�4�n��fk�m��o��`���}�����-�5����phWy��aV�$�g��o)�f�q.u��KdȘo��*��d�Ȥ��-E�)��8����d���X>���W�E|����ߴݵk��!s����A��J����I����sX_R\���i�]�\C���
J�����J;(H��؝�?N@����H���?Рf|�WƇ���,�y��9���X�vt��Uhb�R�H��s�2N��F�q���F�.�xy	�ĥwdrRoc�e�Ҿc�8<t���釛nw��K�.��w��5L;�c�����n��&��������7i�Aj�+&�y\ۯ���5c���$�	���������������������ؼ�>��_i�3�[�u1��)#DIFN���؞�����b����b�T����>G~
����4v�-w�*�A�R1�%` �R{��W�B��-f"؁.��5D>��Wk�(��w��1d ��]utT��~F�;��� ��qZ���	���A�;2���e�	�vP͆����0�.\�١�a�G�aZnd��#�ͅ�[��""N`�]�()j�1r70 �tY��n坙��ZY�֮"2֫\x/_�AFY^�	Ӆ��*F��]��wi�t���3��D�r8N���=%���\���U��������_�D��D�ey��$�74$�%�ofF�Ϝh��U�,���D�?���;����d����Kd����q^9�L��^���ya$>�^���맬r��15
_|I4,�a%sp�E����>���]����)zqV4�-�i�������`6�)S�EG�[}�?�F�&i?�-���HD1�Z���-5�!<|}7"��]��4-���f1l���3�\�0�}5�"�+G?3���W�|�0 ��l�qX������Nh����5�N3�3J�M�LJ*M���9���hk:���F��-��J�w(Z���t]?�;�Vi)[��t]���m*S�3�r~�h����@�ohT�[͔0�v�~�̄�KϞ>��'e\49)���Y�NO�J��Z\�j_��4����d��6�.犚�y�QC{����I	��������h<~(H���+�I?�4 ��h�ߘh҅VʙG?�i��Z>�湵L���rŬkr��.�` ���m�e��MB?���U{�^������>� �F�:#=&R�g8�95j�t��SNi5��k���n�p۹F�����nS탍"�v���b�5��3��JSBk�m#@3Z�S�{>��~���%�Bf�	p`����w2���.�y0��F��¸z����xO�f�d<
^xQL��L4� d�U+��WЊa^�qmD���G�e�e��(�@Q���ih��=ԡm��&.�h���kp�Cϸ���d�1���"2����H���K�ãXn�ђH�]k��pl4ڿ_��� T�j�#�I��������]ɨ1�]�Оp�}iў�}9{�l��ox=�R�Ü�mվ��a�h�F� 먇jM����0���c�G�m��hQ�8!ڒdj�e�Ǒ1����/H�WE˒��^0\?��O���O)#�]����	5��p��ڌ%h�U��b��n���#ǈ|6��M��/k��Q[���M��?�yS����f��es�_�73� �����KFd���?8���(&�vc�}�0��.oU�[�o��|��p�T;�L-ìB��j�X�ٙ�c��Y�^L��ߵ�[�+S�kN��.��9�X�����E����i�=1�-n������4wj	�c�
$���k�#�e�F�Ơ�%X��0S�C~C���80(��BA���X�4����¸�8#n�/�pѺ ��ؿ�!j��},.�x��jNM��%2��?�������7�OV��UV���x$����J��oP��w���zh��r�v�[uhzM�-���2�8�ku�]�sh�����n�a�7��j���ҏ��>���'�B�^{�,��Z
��� M��q���A˫R��fk䱆;E7��d��fD.okT�gxɼ�[#9��h(.�6�{�pDE���|QL��H�q9J���:A�#
U��J�.�r�2�e�h��㸋���q��"bU�߇�$�w�h&Ѝ6|���Q�5"=���q�� %���Hι�AڷG�R����Ԥh�ѥI3?v��WVV���y�&�e��4������.X�0�<�d��R�|y��p�n�$�j�1�K�@�ڎ��"4��c��)��/�ܠ��r?�?|�I9�Km�b�v�G��^�
SK��v���$���U�#�32"źq�e��Åy.�����P���ϙ�Z��g.�a{n��V�剫�~idzj>|(H�󞇂�L��ya6^�2��Ky~� H����<H������k�����b�?҃Y�Ӭ+&@Ү/2������"�@1�ˀ1�_��iW@ׇ�0j���f���ס����:#�7Z���]r2�"��I�blD}O\�iW��+W>z;����v:f�8�m��?���QZ��4�(�����i�/��~�z��L�8�L�m7�֤]���`Fk��i:��H��Dykd�����o�.wϰ�i�`Fn���*��ynah:������0ĨgD�_�|�q�n�.��������2���}A?0�Kҿ%ï+@�G���1�����?_����Դ0�VW���%3��w�WX��{:M��\�(4�Gw	s�+e��d;[ 3�.�`�u�\�=�z�>8�c��J�z�=�C&)��+6��Chw]�|�uW3<�׌��)�5L>��KX��(xF�����������������������J�f"Pp0���3�M���⬬�����qa��-ˁ��� �V�PIfv/_:�O>������08�E���#n/�C�VZ��E� �BQf����D�$3���;M���
���t�J�f��a��w\G�⺟���5O�յ�f����U��Ő���m�Z����B��lVɸ0���G�Z��l���`����R��$�E����A�{����t�ޢ<'���s��/Zq3�z�ɧ�����m�/NP��'��ma��������Az��0u�h��[-�_�hE�q^)/5�i#ò5rfG\�6�p�a622�h�ɚ�]�>?]���d�I�Ţ��3@5&olF��Ԅ��#n̟�;2��A2�8mG�݊a���{�.j�M��G�%�cdV^F����9��v����"���]��"c��!���Ȉh���J� ���w�y;�O�s��I���:�tKx�?��+/����������� ���߂thP�����#��V�IO3z3��4ݾ	L=�c����V֖��bL�R���A���z�.u(>��(3��+��<�����%p��d�p�����g���.;ݓc^w��F!�|�L��*o���ݴ�\=��ѕ����L�
t���e`^�;�����\n��������u��ҚZ�/�Q2#���C;2d��χr�Q�l�v����z��1���;�9�a�+f��L���r)�S�T�Z�`���|�,�b|h�H���@��U��TK�f�Ǆ�o�%�����¤K�~�ݒVW�?��,�[]���{+�k�]�+`�q�E?���
�LV�]�.��D���\Y�zɚ�w�Qg�G��Y)�q	�-JK���:�����Rv�∌@s�x�մ@�c����a7���������������������2���wF����c��	IL���	co���ü����{EfZO�7Ho?yg��-��0,.^<�3��1�#k�E�x��iH5�e*vzE,��BK.�Eha�	Sf�ah���Lx:g��6k�vD'��ٔ+w$�Ei�hF�}k�E�S�<�.t��{$�xQ��:U�K�sj�NP����c���_��?8K��""M{��՚�a$�},H��ٿ��a�
�W�0�^|A�w�z�Ѓ��0\NKy���Ma��8q"H��q���̳�ia�--I��:�OM�tQ�vS׵�hk�5�v�'Lmm����"^Y�7���r�.�`p!�E�
��%�nhx�*���c�~�KV>�K�\_�(���}�n���%s�̹ƚ�g� ��q�����Wg>ccRN����}!A�f�u�>�Ua����r���� =�_��9�sfV��90�^zI�zoý�;��CAz�}����/|)H{�q��r����nҟ��O����F�&S��|.�V}���yZ3��ٵEhX,���t��GF�IuAH@��"����f�I��F�L��f����Ԩ��z#�.ͦ�2��~�bc�����3~�P7<n(��<�s�r��H�W�8W����8&�����N��{�c��Ls���ݿ�w��zI�ךi�y��=�H7^0������&'��N[��F1�\㹛�D��|D����y���R3�y2p[M��C��	2�*�'��F���ˣ��KNM[�;�+G��ac9�g�l��(�����X�Ԁ��Z��W+XyT��U�m�r��WK6錽�vNf�i����x��0ϝf2:��53��������`���U���%sv׸~��}��}; ��>��vʹ[�a �5�jf�Zg����_��&E�"E��?�/����_
؄#\�.^��y�ƪ,�Z�[��!q]\]&K�.�{a��
~_���BY�WfDsj�h�> .�Go#�@WC̴�]��9����������"@�<����ȕ�|���m;r]wh�it�a�⪥Mш����,�gl��������UL�Ç��w挸�.-
3�����6��9�33��w����CH�q~az�	588h�7�"9���w�vR��yk�z!ӯU�����nq��>�r�2if���e��(M-���5��m�7��a������v53R�C��Hڍ���~�����;��0B���*�0=%��G�����ҷ�z+H�W-H�%HM?F<��{����}"H�&_o_�U�v�n`����~7�|'����z�)�,\Ժ�bs6�h2{67��X���e�Z*���`y�>�[�CFΛ���ʋ�l���E��!�N.�(�_�Dp�+����$F�fv%:=�jm�(��H��3"�����N�}��#�90�im���s���;cɣ3D1�BW��2Z�������.�	j��g�ΗT�����3Z}l֩���a$�n}����M6
.&Y8n�^��F߃d����rq�r�g5S���h����zi����wwq��Y�L�lVZ�
�!m
��yX�P>��K����=0K����+s�����ƽ�����+=B�ͤ%�u���o�@Jj�%t�>�����4���X6����̋9ʳ�h�oӿ+xF�������������������@�KW�T��d2��`[@��q�E>���dS{��+o��O<#�/����@8|H?ͪ0�&'��w��� �FTyA�vC��-�f_wVf��
��bF{��\��k��c&wX�"�ʐ���,̆�`��y���wI�{�]�%և�7Q_�63ű�n��u�I%:�2�r�s��n4�C&V�K��*O��aGǶ��V����(�9��5"1��*��W_y%H�|�;+Q7�aк@d� ��3��/%H?�����r[��*�g����;#Re0�H�����aҐr)��r�jO�]���U�U�Y�:�Wk�F[���ڿX>j�E���a�P�<�C�r��'!5;������_�L���\�^�jS���z�assҾ&'ŝ��#�(���� ����g?�� =}�t����d�^�8��D���-�����H9��Y_� �2�o7�W��L�t�g���B䱈|~��5H}�� ��?���w�hd��V/K=�O?��R?U��_�7��?��
�cw���/��/道�[���VG�]�t�U���yT+Z`3���l����l�e��C����k͌��N���'��tZi8n7��;E�j� 6�piai�����9�s1�_�n\�Ps�bZ�{O?��}��O����ϋ2'S�BU��?2�?��2��MR��5��������.�j�s��1���ʕ~���W�d�����i�R�f4�~v��
VZ�2���nF�;�gm��\1�����q�$W����o����n�Ff4�Ȁ�b%@f��2��,+���-�]a�'� BZ@�4�Fލ���LOOO�iS�嫮˷�<��q�Fe�[Uݭ����S�"###"����;`�1zmZ����:v=(F� ��N)�]��K����5����'}�&}��!�gmd�W�u;��g+F����t��y ܦ�������%��t�m������10�� dN���>&,K�YVL�NK<'�	�������O~!���
�gr�����㰢5t��c�^��=)L�[oxJbw�Q���g�h��8q,����5:$�6��+�L�(今�h4df~|��gv����m��}I����jy��!VB4M�G'��3~�1��§��c�ej*y�E���痞x�\ �Ci��D��}�v�7�d��ژF{Έ���T��0��f�_<�>��u�֚���8_�6W�CUFx�!h���>��?��H�|�+�߾��Μ� �Ba�%L�|��~`�Vi�O�N�E#S���RJ�_x��aD5}6��c�̒a��X`,-O�)j������Lȶ�
l�|��f��"�/���P�t�V~�>��waa��q�ؤg�S�e�8Kes3>L�]�wK����z���Q���k�1>5%��s���O|"����f��M�q�0����g>��t��=�O,���&���E0U��.6XU1����/#_?��ľ���%�K;|�;ޖؑ����/��������ω��#��xCbO-K���{�07�3?�������[OT��qx�6��j��&���C�a#�a�e���"�W��{^��������`�ʏ��Z���ђ�2����z��&q�h����0�T9���F��O�g�LB�/��yyA3�F���v�#3T1�ɰ/2�<��K����S�1nD}&�/ծU�+<�X�������!�[Ie�#�v����}S�ݶj�@i�fh�1~#�/Z����f?�\J�}���+�^�jG��c�X������5+��b������
b��c�i�e�)�=��]��~*�Tr��&��	FF�2����a�ؚ�g~���N9�^!���ԗl<�w~#�/                 �
@��>��S#2��ψ��_�Fb���{{�0��°��c[%�LN�&��Va^�kv��ģ��,��jU����D�N�.����h#��GJ�L/<�����������	����{����T��f0�r]���(�뎍I�_O�ϣ��@Y۩�f��&�pն��t���3�m'j��#�A���C���>�k%��u�ܔ榉��ԱY����*���/-�s�B�������&YQ���z�;�gb��_��7����h�w}���=yB��k�a�^I��?F���ڎ�;�O��`d�c��-S�y��hb�y����`��s+R>]0�f����9����3jj^د�0�\���`��f��6ñ�F��.��}C��L�9�T�-S��8m#�U0��=z@����fQ�\�+��wob#�3=|���O�I0��b���Ab|@��g<��{뭷&v̺2�U��|)Ol�(}������(������7ߖ�;o{zb����;��qh�M�>���y�sd��|ߺx%ӯ�����f3 �~盨jܡ<�$��	�cj�Ξ����[��������3��i��������ց�r��`����]�c��봆���H���RF���gP��T;�
\,��a�(&v�����h�7����cZ���Y�zy���׾��"!��;��8<?V���	�2�`�hZ�/K���^���T���2�W����Z��e�A�Vi�QW�C�����9ۅo��/9���8R�~�Ǖ8E�����i���X��0�q|��/��<�ʡZG���Z�f��1��;����kƟ,����i/q>�0�J$�~�ڏי�پ5������d�-00a��V.�C�]2��pն�0ܨy����}W ܉>τ%�ZB@9�GN��_�?��>(�5Ѻ۱���^�(���0�f���"������}J�;r\�>�v�N,�Wv��ư0iff%��<��+0��}��1Z�f��9�]���ں?��΋f�7�Gt���46!���Q3��1�טk����Y�{#/3ωf�<����zj��G�:#�L���(B��N3�p���u��,�O��_�b�5������6-<����ȹ�	���䛢)Y�[�7Q��+�(����I�"�L=-�,B�ba��Y5^�����*�˿zOb+`��t�0bo��6��ǎ��&��.,,X�BO�i0�VVd{�f��4��C�l�	�r�z�W�??/Zv�!aOM�	!��|���9K�]ﵶ_^8��U0��?b�B�z�9ëVa�/�S���T{D�cT[��9���(�J�Q���t=�Q}`���Jch8��G(�M����s7-�4z4V"yj���R�|�w$v�?��?J�;����^{�|���O50�K(��}`��m|�(�*�%�״���RE�3�!���>|H4-��w�=�?�J�/���Iy��{��჉��?~ �۠m�<'��5/��A�����T�D|/M�B�&���ѧ7�xcbOO�(�Ԫ����|a�NV�0H�z���g~o{'�v�o���|E���0�S�ڟ�Q��^g1���Y��,F�催��>�a���9�6q�4��ZzYZ��fT�v��P}QVu�������ׯF�eO��E�����K��▩W��g�%�c{4��2W!=U����/�~o�wM�.��h�1�'fLN'ֶ?���3}����ߩ��Q�}ߝ�և��t��U������~��h��h�Ǚ��0m��m��u�f_�!�=��$�`�V�?
�޲:D5�vVJ���%fNu�wt3�+i�k;C���Q����Q+Вo�V�����-���B;�q�~�
�u?]�x��j�N�>0�� dN�i��n�C^�xP��>���&�����-�}{��؛�z{b�O
�`��=�}���{�}�%���h+��r�q��{�q��ڳG�}���gn^
 ���ʙs淨�bd.���!h��0��mD 50~�F�C�K���o�蠣`U�X[�h���x6�L������5�S���pz�Upz	̴b���Qg��u�x��&��d��0�=#d�t���Ct�
=j��у��Лq��q�D|Ֆ��.F�!���PKp���������� !uY����?!�M�_z����
ʧ+��L�*�+�u�wߙ�?���&��g���5?�`��D����Zvd��	�h����;����}�6���r�'?�I��2�+�O��Y����~��a�_ΝC�^���0�V�Y�|N����$wQ�΁��3�Z~-ԧ�%����jw������+Vm�s�J&[�6��m �1�G�ڌZ�HU�_kQ��:7-�c�x`�@k�0F�"�mEiQ��v���K�nϟ�򞝕�m�nN1��Z��;.��3g���o�U�<��ظh�v�Ơ�Ƭ��w������a�e������%�]�z�/ߝ'=Q�c�hV����k�'í��
4_��VѮ�h��%R�H��!y]|�&vI���wI�������r������{����������h������W5���w�h��LnO^���#�1ܶ�ݷ�rsb�z�M�O0Z�􏄹x��Q��v���ځWS��s����=_p4�i���%����7�zl�?/#����1��x�oZ���`z�/r_�4{KJ�V3&���`�,������1\|?·�C�x��2�4 u}�7��o�Ɇ��j��������]:�����W��L-f�s��W\	Ļ&��j���RF�J���(O�����mf��;֛Q�J����F44v�[NG���p�*���3���t;�>��AS��{2ϡ]&#v?�Vt2��d��<4��U�������FbL����p�+v>;X��F�7��X��Id���i�CW��|����w����hº<����wW=?��rU_#·�s�i�����>3�H���0�0_T��F���iG���s�8���$�n"���tS��������9��Dς��0�`�|�~�Jx�Q�ҫ��Yp�U�%���?%�����h�'��W���|K��{̛M������N�!=�]'�x]0#��̌W��(��6�f<��;��ã�(�d��e�XEҽ�:y�#gK��i2V�"})�"f�;�����g����v�G��l�	~}<�$�s�)��fH��Df��$R��fT�ر��8��hj�@���ַ3G&
p�+ͯR�ִjw%�;������)̴*�+Cа�5���!�<��Jj��0�b���#�<ai�I\f{����0�"z�Č4�}T�e�&v�&�gciW��ڤGD챣`�n�v�o~�͉���%�;fVp~��W��$�Ct)�Qg���F����s����Pb�~F����#�_2�������%v�5��fS��:5��JƖ�[{�u�M�ݔ��ccr���yk[c�3j�����?���#{��M죏��v9�?/LFj�1�9D��ja�m�$��Eh...Z�#�rl＞�!���qj$6Q1���/�a���j��������26*��Q��;w��8|D���}�t��G>��*�d0�jb�d���Y�'�o��5�oj����}�{z뭷�sof�r�[�'èg1��x���[�c�C�f�K^,�v��G�y>�E�a��xZ��"4r�7I9ҡi�����t�g��vj������:�����x��^,�Ynd��$��n�!�,��QɮȚ����w.ՀY���=�>�~�Mz�WgteE3͋�����ej��}��0�5�IU�55I p�S1�\�d�ӽڐ��ON�c�7���8�^���͇I��h����ӼUyAmT�d\��Z���կ��'u�TkS��� ��{��f��Q�Tz�w�թ��a6�S�_,�}t�|�=�M5�����bn9�_���_1p
Fˎ�ߛ�����h���	F���v��x��
����P_Xy^��f��b��}�/p%�����X��-S�d������ńe��q5�M��z���_�sv��W3���7���s~�ud�!_��s�����{0+�4�ʌ#0�k��|~���������h��x���#,�uY�9���J;_�љ=����t�~�ի�,i6<����Cq|e������ގS�u?�V���LO�#W��	�0�R� ��x"�����h�������Pv<Jڳ��p�4��:rHY�}�=s�����d�ع��Tسm_b'Ƅ�W�����0�&�q�i3�i.�L���mV�f�$\BM�3���a���!�u�v!���B[�L j�t���*�v5�"x�8S�m\<?��
���)a�Ml���HWky4��{{ �YY�%�g�I�7��{�� gҩŲ �&��"0"�Kr���=���p��n��M��2.�.����i{<�<c&�.�=h�ܨ�C%��uDQO�
��`P�M{$�	Z����5�:6c��m�)��`�׿0K�1\%�5����s�m������/je���,L�_�O���7����
rnZ<V����
J���dpb{	�h9��u�h���4%eʓ��s-0��r|��x�i3��=wO2߫{Lu��G��2�*���u�W�)���Xusb���XZ���/#?�~0�q^f��]�$�0jT��kI=�^iY��(���8=mGOe���a����	61Ϳӧ�{�f�Ȩ\����|OMxr_��.�?��W��d�Dwvel��g{�Y��V�	Wʒ���O%����|�N�a��T4�L"jq�+h14��	k��񺢪��S�2�<�x�m�f\���ֆ�}~��w'�_�\bO=)����_��a�Ѯa0�1�*J�a(���a ���xz=�+ń�1ea;g������I�+�����Ϙo���#\}U�Z�Ԍ2�.U:�G�7��S�ʉ�j�_#��z��d�g+Ʀb����Y!/#Eǣ����Q�����{�_k�m�,x8y�ctR�ux͚���:�G�s�CP�<���y�BFÙ��t�<���(��v����G��g�|���c�eEIM����Hڞ��+Ųu��~J6��|��+�>,��ڸp� �S���F�yd���0�{�g�OֿZ��}`����(����v?��i:�{T}��Z���e����ߋ��@&o���4P��t~���Dd��F]Sqq9��A}2�#U����ߓm2Ì��d�7c����<�w4�xd������wA���������{?cs~׽�Gz�>���(z�- �|_�4�n����Qr=���7������p����yTV��)#
���p�§����S��س�����a�횒h�C%�@�5��f��I�ܷ�ȩU�2�I��g$�bS�S[��R�T�Ң�kjB��K�x;
F�6h{U�n�"�V� ��Y�=f��,�3В�a0��ba��>"�G����Qi׊��x��5�mX�f��4K��qO�=���֜3Z�0"z������gd�����:Η|\��GG	��x��/��$Dm�Գ�(�� �n�_i������M	��KKMX���C�lf^C���������K��v���-��w�r=��"<|���`�}T�LU�`A}�g�]'��=��_��}�Ӟ��믾^Ϋ�m33¨�v�5w!���C�;�.��R[��2��w�����O~����Fbw�(�;�#�Zn�BF���zyz�m�$��n�)�n쏈���{�R��e  ��IDATSnH��h9b�'f%xn�yW]�|I?�z�(]Æ�)`T�jUʻ-I�A��I���7���9��ۼ{Һ�c�oکǎ	c{�0�E��u�J���s-lo�v�u��֪�����Z�o��e:uj����*�i��g������y�J>Q��`���8�~�/��e�#�g߽&�m��#�O�?�7���-��y����j������;��O���c����J�NG�1J? ֶ��9��'����N	�<�o{�0�O9���=F��Ұ�eL�������f���o������ƃ^����,S��%��3F�� �7�x��>����SĚT�����_]5�*)&�ft]�a�1b�o��w��O�/������m�j����vXo�5�г"C3�}=����A�ɩ����o�����C��D��#�ܡ�[�����F�\˕�����υ�ϭ��ƾ��~L/����E��Ԝ�ױ�Ò�h�����oh��aW}���N��W�:%+G8�:�?5xϞ�������Y�����*~Շ����֡��g��=��)�:�}�����K���~oT�¤�;�����ks?��\YR�+��A	�&jnyuN�Mf�w-�+&,o�~����QZ{jR���Ȋ�k��LTe5Nv�OoƬ�m���8�]������(o�����NM|���+�_��;��~n�&jr~�t��
{�.�0p>5t����������������������+ f�ϧ�afn1��F4��O�N�7�{ ��eٿ�a���&�zQoW�$�vD+��`�g�����F����m`�T�����'2�8QJ�7c�l*aF��5��8�	OL�Y��F��ѓ5��D�]>/ϱu\�:%L��Iw���f���g�ωqz�8_�(c��m3s~���s�����0�N-�[�Ѥ�8>m�;���>�aΝ8-L̃G"�d����8���*j=&F��*3��Ƞ�]�����0������y�B4�eh�-Bl�� ##� �����xwbwN���,�_E�����Pgg�@B���ya|mn��m�~�<ψ��ۨ�~��PL�v�}���D��/����~���sz�O�1�9L{SL�7H���$l"�n���� !�1DF��@�f�j�8�Ф[�ӅBh-���)��e�G��GKg�`{ʲ�17��J�������}Q4���`��A��v	ڏ㻅�Z�"?F��fԙ��h��m_��Ǎ$��NL��6	�E���Nfs��Jhm��cj3��,:?+	F	.a��^��wxB���ي�-|�SG-�����}@�\S��XkϤ�)w9,�|Z5�~|�c��=����,�u�J5����9�)8���|)&���en��"�|sZ��aZ�}Eݞ�}�!�w}<���W9ݕ]Ni2j�g/����Y<"��e^{�|d24�S�r��Mn������'�P�u7J��1�*�ɯ�O��b��f��w��wD7���X73�p���J�
~��ۻ7��v����-���ab��d�@+��P+�*5�C�Z��e�<�m���_죸�߭��5#I�0��8Mk��1f4��m{��A�<��(��1�~��]�Ve�v�t��]�h|�5��|>�q:�躾u;��H����K�w,�tLzHG��1ز�������4�2�8�4�y�a��C���{�����v��T�З�NPW�'ӎz���x�=��j��K*��!��qdP�r`l	���/                 �
��ѧ={Fr�ÇK��ێ��v��]�[GT]zҹ$�m�z��l2�5�`�l����h/=��G�|�_��9zL�܊�����k{Z	d�4�2��(}��"��P�Cz0�x~jD�(�A�j�YI���S��Ihd��U��=��C:!�����|��h���3�]�Uю�������I=>̖�)ў�(�VA�"�]{�hsM�
s�����Qg�L��l,�M2����Q���<��2ZY�h�d 1J�mi������=rT�_�=/���
 ����u2�ˌ*��&�}��+�a��t�1f<��������l7ψ��O�-��-� ���@��X�v>���ۘ@�SŤp�s@8��BN��(WUht-��!0��e7:"��eh'���(iW�~�>]�
�Q�֋���ܨ�O� �����4R3��zP��_34aͶU�=�dZ�G�W����N[Ȩ�FS������&vqI�Û�]�hh�0��m��G�i�c����D��g��4�Te�D9N&���ϭ&�~�o������d��HI٢������z���v'y1�y0F���pr��8gG��X���a<��;m���h�GQy��Uk�9+T6��������8�a���L����L���r�����ǤZ7x��+���s�7�;�U>�F`�t��0���n�z5nٞp=�7��4�����;�x�Zّ~��?��~�~�^Ѣ���>�X�P���L6�2�h��+0z�؝��xÍ�5=������Ɗ��Ѿ&-_���>~w�C򻻂�k�aLi4��ﳧ�"?X	��5?Qk����el�q/��%{\��i�"�/��(2,�y��9E�{���Z�U�Z��/ٟ/'_�;�cVr��j�>-��ncEb�BΎM#����e������w�=\���E���>h~X�:ZxIiಾu�,W\���X�Ɲ~G��V��c��ձ2��R��b���~�Q���7X������\���D��������������������oy�u�T���k2����w��֊x�G���$��R�$�*f�u47jl� �b�����;e4�S���O׼s&�ܴ0�M���
:��P�oQS�f±�����N�|-Q��^�͙��e9>>&ѕ�`��!
��E����c��|Qܴv�9�hX�����%�^Ϯ�詩}z0��h�|��j���d=�<'�=4ʃG�!�/�+�f�4��|0��n�P`�F0U�d�tTA�҂���LR�.�#Dۭt�Q�-u-[�Ȓ�jfJ����u0� 5ѳzk2xa����.4�F%�@M�ڨ0&;i�����]���^��ʗ]�'�s��Ҋ0�ȨrWl�j[�mU��k���sa3��-'9�[�&���
�����f�v���JL���a�h�� '߆iN-N��ܧ?.��l��l��	����/�4�`�O��m�&���qXi k�z̋���'u�=�S�w�-�Q��$�n��lj�pЧ+�-e1��Z~�U��P�"�������+����;����~_�o��>����HS�t�{��#�z_}�����ge��ՙzi��g ����w����ǠD��K4�u����n�gy+��Ə��R�&#JlJ�g����ӎ��'(I27C���	��"�`s�o��q~o�N���"���]ڦ���"�!	Ϝ�߷͖�NnB۞+�t�Kd�aEΰ���J�\?6>��Z��("?r�����mk���"ahX������1�=<4����o4��,H5�+��`��G�c�hk�q�QQ1��צ���vx��<}}���W4�>�~����e�;hk�y�~=��o��J%־����J~PB�aĕU�|�v9C�킿�h�E�)ZCl>��X�z�fd�'�;��L�������v+X0��p�d~�I����L׭D��*�����F��x|8�$���fD#fZhe0��&�[� :g�c��W�t�v��h�F33���+��0���3���'3꜉=wN< -x@���X�v@�E�\cO&�a_X@M3�nS�Xj�F�(q&�,�-�QA�,�}���5�&�5���"�<z�YkU�QQq~��v�� ��:��(ReΜۚ��*�@9�v��ڞ�4�#�kߟ0��a��`3pQb�èC>��������vͨ���u24*��ij6�#h��%a���tR���Js��FMjj��MfD�5�0�IS�B3���׮-���u�|�ٰӨQ�ij31�}j��e$��� ��_37s2��)�bDf1P�A�w4��TP*2�SF�9���V���1��-��K��&SD�!D��<��|�ox�T.<L#�6���f;��w����$V3َ}~�h*Ễ�I�n{�;��!/3K{�U��b�d��	�F�	�5k~fv���S<hg�2؉T{V���D��g�w�r�i�ź�z���a����z�j�Z-n���}��։�1�f�y��n[���U�v�����=��6ke��ݞh�kM�9�d3]������PTL#���ͬJ�%`x��4��tz3�F��fx��;��T�(銝��0ǩ}��/)�ø}tX��W�4U���dk���Mf_��3�&J���u�.y.�^��m��W��a�1E�	��v����=l�syY�3���}Z~8>2&��ah�
�o���:~��w�~��{k!��5�}��Uk�q�֢��̻�u]� ]��&Xd3�|�v���׹'4�O5Ģn�N�ko<���a�{J�P'SM?[���^��S3�ώ=0�U?�v83'ѹ����_jI{]lɼ�BS�Oǻ��C"&���������t6դ�V&�@�|F_@@@@@@@@@@@@@@@@@� 7�Z�l��b
��ɓ�]��[k�w��)�Q���zŎ6C]�b�7��+��ŠPmۺU�|,,�(�����1Zj�=�}���`%zf�d��q2ߨ-WS�2gΉv�<d$Vv	Q@遈��w�u��׃m4�<��LO�}[��2��|u���g'Ǩ���ԏ�)'F�[�rZ���9���
��pf=���5����g��O�7�=��aD�^�u��!ќXXj"ra����4}ދ^�؏��?%���niG3��v9(F\�`;�
�������_�tb������"�C�d3mY^fH�����<�;�{��y/�y�����Sm�L��`�3�5c4S�������f\z�?��:�����U/t}%ӫk�����ǋYQ�<��a"�t�at�e`(��unu��*Nos�j��Xv=�;mk?�~�S�z�/�{e�����~���3ڸqCcӔ�&���*�a�]�v���e.i8�x@ͱ(���w �M}�jr�m�����_�s"��q4�
*� N����]h�����L��"�dA?�/�a1g����*\ZD�n�8�>�w~v�v�����i��=Ns�껖�\�b�v�^�I&ͧ���U���q���J��ge�~��W������n�FαcG�Ҕ���3g;fP�e�&�;�ж��\j�Q���bxf��)�~r���?=�'��<@����
��Ԇ��?�?��@T]�~/�YH&�a���a���2%+���Gq����>]��a���ߪq��^�����K�>�rM��Z�%�?%�ی�+�J�8s-���l�z_=���x�@Q���iʸS-X����rV`z�Q�K����{k���-�}��}�T-��������>y�qٞ���X� �15��Z����*�-4�'c+O���L�+h%����P���Vc`3!Ξ�5��O�L<M�H<[���^��F=�)b�s��qf[EO!C���b�w�Į���}����c�b[f6�5�M0�*&
���*0�	��t=� X;�j�!_�	c�3ã`:r&w���4�|�	����f��r�]�g��&
!=K8�x0X����p<���&3��"</]jMhO��|&������MD��;��T�`U=�$є�'�Q�\��̃Ѻ�(�]jF����[���(���[�I��>㹉}1�����%��q��1��
�c���yI�<<|cU�����[;1$��Y���)�}���4�3��ȸ�Ţ?���C�E�i�N�h�Qsȩ��p���m�d�Qp�����O�/�9��O3��L��菱�y���ۈBV�G�Ӷ=S�)⫏z[�?s��^�ӆHT���TB��D���Οʗ��D�ͨ2�bF�"��ax���2U�����$�91���"������v���e�W4�y��ϫat��WZ�:�W���v�R�VoO�����3��������:��D��Ɲ�;��Q�r������������l��0{lk�������y_����2K�������}�>��f��,��;��ɭ����]l�� �!��	�Z��L���;)c����ܕY5���}�M�T��*]���ߥǏ�H��4��Ebrsb���	�mu��6;/L�3g�9��祒���ҭ�-���1+��-X[,��d������"��t���[�]�uU��e�)���wB�Z�N�����-Ṗ��8���1�^��0È�]�ʿ܈�|`w8�&DKm|��
��hV1?Q.�Q`��|~7Ǡ|��V�����H�/�f�'��3��S�y�XY��>�ץ+�򕫎���
G��5j�#�-�Ws� gtӖĞ:#+�=�����������e�uvN~w��d�L`28��<��
���,�
V�1�c�mtcԗ��	�F_@@@@@@@@@@@@@@@@@��4�b2�ڥe�)$#��5�u��&C!uhK
�a��9��a��3��	�0:
��Z]9�����Y�K<�+b˥�u_槁������z�3�i{<�
�A���cT%2�9a@U�}{ba�ϒ��V�}i4�����203���Iw�f6p����,Oj(������<�Y'�6#�x�4#���cە%�'g�[Mh=vl�@ϣ1-�sg����������4������>xB�Y��o�Zb�)��Y��\��_��7%��~[bG�R���+�_{쫉ݲ[�uϝb�ź|���G�:/���u���=v^F��d24#�C8r<��B�y��hr�7�#������8֛y���i4��i�h�N�2�<'��hz��L7�e�t���X��nZ��������D��J��x�x}I�;Z};+J����wE�4��L1RO.ۥ͘�ڊ�]l��a��� ��R�v����jO�������������v���ʩM�h\9��*O?��z9N�4���s~�zz�noށL^�=��Ο�O����ƚ5�.nv�垉|����E.��p�8kE���L�+&���v���z����G��67�}��-��q��7��X���o����ݎ��s%���*R^�:���J���U0�{����������ǻa�-�x+�JeI��G$��2V*��+Jֶ��4�{hin��b� �8��.d�vl�=5��<�'o���=��]�@�� �g������Z�V���(47O���v[�/�YY-cE%�~EEy��_'[y�m�yV��т��G�Z��3f�'ڝB�x9�Q�(c��a���n�.��O"���Ya�.-ȼѹ%i&J���5��{��+��_����2v��/z����@`�\�N���F6#�0հ��}��(�f���=�(9<Z4.v��Y�U�Qƌ�#�e6:.k�z�@b7aF���S3ovVf�g�F{�fY3����|>F!"�2�Z`4rƺ͙��ο��S����N��v��HK��`����(q�8N��e�!���X*Z�QC��"�2�c���RM�21�.B�-@z�ZЎ�>0��v��2Γ�O̊����_M�K�/̾���%��/��W��O&�s�|泿=�W�:���#�}�{ߓ��-�!0:��z�|H�6#�h:���8E���d�זף�F��c�2�0?�U�_.`��e��W��5w&]���	��(%FeD���"_�h��L�#�����n�dh}n����C?E-��L~��!�%Zc>�6�l6Ls��������Y�&�J��g��i�dX;�>�U
�73���|��ut[��V�,Oz�p����;#(��I����{��{�(m^��{m����g���|]6�h���Rי~��ti&��_��"�/=�'2�\����_:nA�Mf�A�FE]@c��}�Z�	O3���N���.�l�N�;V��mE]*R���>GT�Jui�yQ������rF÷`�}?r�V��8�^�q�V,�w���Ğ��r9y\�)�6	���&�?��2U̻��X����:�߰WL��j���v�ͼ�ђ��m���h��s�����Je���<�����yk�$l����|��_��v�R�1�Ś������9a�>��<_��Q���L0�`նg|�vCz�c��}W �'�R
Zb�
�,O f(9�蝜�-a���cÈ�2<��zVf^x4��&$
��G%vb�0���'Qy������Y+˲]T3Ǯ�g�e�l��p��h&xe���[ϝ��4x˫�>؆<|��8�}���v�&�тS�M:�kꙢ���
��L�)�hUK_�&Zx���t�G��hu���.�C�[������������`���ZF��������G���ѭ���ST�����蔃fnh5+�)v�ٗ2j���JT����eyL��9�Q�nyZ6k��Z��Wߟ2��#��Q��}�(���ӌ�_C�7JL:Wk��y��-�HG������#k�غT�Z��{����iҎ61&J��+FIv6$��9����ւTcE1
v��P�6��X������򗍨���w���>��w��qFkv\۞��m6�=/"�������uʉ�������oL�b@f�^3�R-����L�2��љ3��7�{��Da՚_*]�ޠ��C�oZi]� =���?6����p����f�
��ܶßw�
��L>�<�~���A����)+���Ձ�e��{�n������9Y��d�R���,/qe�D�={�<�'SL7jΩ�e����v%��C��!�A��Vg�+&"3b�T�c5�L@0�L;/`��t,��g���b1T1�41���l9�XY�>����-��6�8*ѬK(�ջS��ߕ����N�W荬����@`�\p&�RO��_3��Ĥ+�S�Tlv�Ǝvy2�P�g��؅Y�OML&��&Y�>}vں�7��@bw�؞�V�l�D?ݍ���֣��0O��+��R�]h����2�fXn�H坙eB��p�1>�d@"l�фC6����Ɲ�h�$CT�����S䱞�/h�T���Q��{�G�JO	\���G4��q9�*�z6�h�m����
�G&�&Mt�no�����Թ��O�}�}�b�F��٧��?���jFy=?ނ�=��`Z7��%�f���G��z#��<RQ�"�k��D�󔻏0�^��f28Q�y�e֯�9~d�9�Kj�F��6�����\�^z��I<-`7�3�����\�~�������q���a�C�ghD��9���� �n�
�K����0����b�����~^ݟ�W�ɗ/[�g�v�c
8�Z[������g0��f��~�����栭e�{��S��<��q��;+&�E�S<�5�?�xtj��Ğ>~Ln�G(P㬫We��p3���$l&�3�v[y�`�1�S����{_�������H�U��|+�2	w9�w?_y�e�����Y��>w)�1�C�ᕕ�}���{aY�=]��d��z�ŉU�j�5�j%��(Waz>���uo���T�m#C8�6�%q�G��vi�b�_[j��ڙ*���0�S�#ݼy8�5����/                 �
@�>%E��v��=�K�C��@fƗk���rF�e�[��ƌ�	�B3O�	x���ݗ؇��`b�N�o��m���M������W_���D[YX���è�%����zF��T0Qe8�m���w��r���8�V�HM4��e)�rE�$� 1�1��r�h|�2�=q�^�p\�j[QPjC6���x�������%_�
�Y��x�����gߙ��{�+{�Dq��ݟJ����\}�_����M��;�$�_�jK=���э՘Q�����s`:�J�u�F�a��E���D@|-�#��.��v��Gy��O�J����Ķ��:�]��6�R�"��m��ys����s#R�jƜ��V�:�o�~|��R��+�4*��:'��m����}2��&��Z�'�M������Y���V��i7�;���m��J����ɓ��'��Ӧ	؛����e�C�adx[9���m��i��B��!*�~	���_�q_V:.c(���Ȣ8���羝N��������{�ȳb�9�ǰ�7;Y�6�߻�Ǯ��^��q�f��|k�ijp��c����\�+_)����&����6��gV`Ž��m�TV�����US���y����S7��w��)��8o���N3*̪�٦�_�4��b�O}}>��
ǂOsS�3mo9�KF�ѓ;����}ATo|o���(�Y
����H�\��G`�ƥb��7"u>�����5׵N��p`��>N���Մ�T��3�df-cM�HI<ɕ*fH9�L���Yz�}�+��`|��D*�h,b'6K���g$Ji�.�g[&�&�k�V_�#�"j��ڛ��ߦM��Y��
��R)aƗ�#˘6��p^�!̪���?*v}a���Կry1F��G|�5�����`蔚8.%If$�Oʤ����5ɨ��A�c3�����2� �Gc��maRP���?]x ۋ��
Q*J{X>/Q�������-���*�����K��?{ן&����t��D������������u���>x���n�>���ym�砷FC�=yxN��|�̋靎��0�<$ktP��z�/3���=!L��4O�ȥ�ѧݨ���[ŵjl�ɻ;���OC/�zV��;�T̰�H� �Q���)�۬݌��,Ϟ=�ؙ�gz�^�I�;4:*vl�Jgqvv��y:V~�ʈ����&�,����@q��ݽ_&����;1V�}�g�ē��x(v��귽E�uG9��
�j-fif0Q���Z�ݍ*ǜ�sP-��6Ѻ��К��ɗ�=�q��Z㹗r���̍�r7?�8�|��0�)���z\^X#1��2��j<c���G�O�ޅ����@k��:���4v���w����p��p~'���܆�D�}in������\���ь��kR�����������iw�q��o<��Ӧ�>�Gqeeɾ^G�NW�����ծ2�y8}W rO��-4ed�'�oK��2M�x�.�1#ڵgF��-��F�ل�������V��1j�M7ߜ�/|�Ӊ=O}c�V�)�;4$����������[\\���V~�����c"�d�u�`�U��*S�M?qޙ�8�~sʇAg����=v]����3�����&�.n�Z��P.�*!�
m��3Q�mF��H*�|2�x��j@�!��k�g��g�	!���2�rXA}�����"L��D���w�Qb?�z;�C�w�'#pzY�%�������mw$�u������7�4����x��2�c�ޞF2�g���:�b�z^�-P���wT1WÊ�8�ک�<�~����S��5��|�\2���q��x���&w�H�ʢ�sF��k/C+�Qv]�s���S�d��<�E�w;�Q�G[��
��!~�<~^�#����jY��yMF3�c��>��-f����_���EQ] s��1aVO�ڙءq�����r��g�^a�R����ȟ�]�h��w4ݨ�9���g׭��i��~�G�=���3���p�;"͌ꝟ4J�ec�v�U|���,�����&�6�[�3Ɖ����Qs�s<=P�w�\���{y�{�<�G��|P<��g�]��?��/3��4�w{\��m:_���u}��s���!��r�'�Gf+
��=+��P��%��0���ˈ�y�>S�<�3�8j�-��>������ڛq����>����������������������+ މ>�ƘQn�oߞX2���¤:7#QAwN�q2��`$U���N�df���+5���%D)�}wtBx���[�軻�\���W]-�͞O,Qg�
#j'����,<�d�ի´�!J���"�[��`����L��Ͳ��>"�/��V-�E��9��xf8Sܛ��6�,撊v�^��坯��+S��h$ɉ%D՝_��rW�ud�h;?�Xb�ċ��+�ЅY��n�u%�Y���.�������|�r���_ռ0J��O}��a2XKx�m�P�sw�-�O�!��������?�X2Gw��%6��3
#�QM���|2���׳_�\�_S�W�׍�bƑi����H{����xi�#����n�]_L=�����1S��z��<�Q��T�KkԼ�2PM�j2X��4�IY�v^�$�i�>��#���|ޢ�f�g2������5d۔钑=���]�<����AL'�ӽ+�l��{�?�&88�]��T�K�Y�X/�0�_c��`�w�&�]/���@E��9�0ی�8o�}�=u�������L�^k#���!��/!�]�����]������w��&�/�:��9�|����m������L�0}}��5m-�//�f �w�����>����o}kۮ9�=��o�[�Skf>Gq��덺��\�v�z�{�BN83ܯ��3���3��>o�?�<<�gObO9RX�Z�]����>����oSu<�;�q~��J[/��IW.ȉd�i���;�VMM7��s���z/Z�Д�G[����ٌ�k�lc|�q?�ƚy�������"����t���^F_@@@@@@@@@@@@@@@@@��̉>zNuw'����/�2��hb���'^���.u���j#:*nU�L��VK�n�=<�5�m�O�R1j�;'�½��&��cr�4�*8�Q�����'���� �V�9�F�HS�����SJ���(��vk6S����q'�����?��[�����;c�hb���T�M��kF�����9a�:t �M0���d�1��P��=�g#��F��4$�G��M�ʲ�סFS�5�ڨϨ�������`�F���������(d�f����.�Ѥ!<��$:�̢�����B�r��|���x:a5c�x<l�RZ�Z�ΆI�D�A���1�r�|��ǵg>e��La��h�y4��q�*��E��[3X~>�i��]+���h/�C�^z{�r{�3^�_jCi��|���4C�Љ�j�ݟf֫�V�r�'��,M�Na �vq7�l�dm%�{��^�҉;�Gʌ�N�0ūr����V5�����12�#�?���Աc��dBi�[?��H1L�����C	+��� SIg#���QYL��h��N����F&a{�/���O����#Ί�=(��|�~7�̰�n~?2����d�d�A�8�0����Y���kf;��c3�g�0?�nXj�z�N=�~f<���G{^�ۻ��{WK�`mG���}�o�，��qK��Z��_�eYߵ�ߋ���	�Wg��M�0�x���=�>^��|��dz;oy��_��_*F_@@@@@@@@@@@@@@@@@��r��)K�T����u�NѶ������C�{�0���YT��G*���n�'�W̌v<ZnY��RS�T50�`*�ܱ-��ϞI�SEw�~Ѿ��m�Y0��l��W��'S���Ӊ�_��wdt�];�`T��ߨ��<4Ѻ��^)H��aD���h3��.ߚu���mǡA�xN��ϓf�;L>�p�.�O嶼,�`F́��E]J���Q2چz�_-��0�m���dwJ{���zM>�:�����vQ/��L�l׺�h0�:Z(�R���0����z
����+���>��π�*��s(w�3f<�Z�I{��&߅G.<�Xʩ�gyd�s���M��(��㸴�A��!�'#�є�L&��n�=j���f?Nw��v�$�c�n��. e��N��[������e?ܵ=�ipo�'�F��"�E�:�2\���w�Z����W��v�i݇�R��V������0����z��A y��0���EԋK$�K-?/�`��&�|L/�����ŉJX�b���(�����ԟ_fz����Z���{��v�~\3k��>����\�����'���~��}�{�:��37c�w]�@�{^F����A
���Kq��l���2����jK��t��+��!�C:n�J��V�����گ�k�����̉��s���p 3�.5p�qŨ�S۶���lϝ&ܩia�Mlޒ�&=ڸU�HF��q���ǖQT��c���E�_	Qx�e��0��ydޝ:s6�;�J�WV��5>.�s2�N�8��;vX١������*����x�;`f-vD�<�f;���h����95z�4��������(�A�$��\��vɀ���#ʹ�rݺG�����"��M%����F�O��M���W>���&v��v�l�z.�t�7������Z����f�s{�zÕ[ۋf�g�:ZJ��#HyNL:�O�H5 3<0��>�՗���p���f�I�(T�<�����TT�nG�j����d����O�흐�ѧ���x�ѣx�0X>M��Q�p<;��!�j�5�}*a|q�4~M���Ʊ���k�K�����b�{S�\K�=�=����Mϻ)���x��G}]�u�iw�����v^�8N�?�{�����Ȋ���x�V�2����O.O�e�9�[r�/�yYL�~�|K��d���Ĥ��U�^w�������O�F3��E�ʌ���ͼH�V?�����+#Zx!Ss7⍭�����>�, �0�ڂ*��`�E��/F9�1/�/                 �
�����׌�RY�u�'�5�y<�s3��v����^�D�m��!UfT�=��jGyZ+`�����n�a%Kj��5>1�ؑ��-��|�[�d���o�UќFm��)a$��+Q{�#rߙs�Y r='�a�6��R��q�H�񼚀T��a���˂F<�|�,�"����c��97ы[�܁��h�5����-['V�d�EU�'���*��0M�� 4�E�?�=�i�&��.��&a��Fk�Km�B.h�G��Ȉ����ǈў�����A������k�ۦHF�P�&7c���CѴ��0Oh��Ebs���bQ?43�<ך-}=�eQ��4�b���4Y�1�����/%�L*n���6��Ԫ����)S�w���%���N���K��_�Fb���l���	�DŸk�@�V�A) �d�ď܌���*�%�/�Ǭ/ԆM��6�ǀϧy���Ȋ��g�q�߀��0;=m�K��&�e��j(����)�o`F߀���q�mo>�^fF׽T�}6.Ry8�9np>�ﶵF�^�|�K�
��L�5�7e�y懲V���&��?镥j�g~��w��«�1Z�Fc�Ώ���\�ٵ�.�Ͼ�բ�}bz���C��p���|Nt@����ݾs{b�~�5�=}R��>v��>~�0�vO��]��L*n���c.F%��Ңh�K��b�R��Ȱ0�vl���<%�³�DKgώ���0�ffgp��O���؅ya.A��Qu�p�W��
fڸ0��<�\s�E�R�"�rN�rf�F��Q<������N���yw��{<(d��C˱Z�r�A[��cx���:�'��JS�(gjˡ��&�����n��H_�Z�y�.���3����1��qS�e���:0�G@k䌺�;+�:��/9�Z�ag��IVfxJ���ٞ���EN���Fk�8�����e �h�>�>����4�_>և�6#oK���ً˝`���3�5l���'�����Nl��ª+���o�����C��5�#V�E��1��]�V^��j�n��0RZ��?�Z?ث{�c�;��]7�^���9�X��e�L6�RY�c�v�V����Ske*Ͽ7�Y��>&_2����VS��YN�2W(PO��x�9�¼�Չ-�c����Kt?_t]ﶮǫ7�+>�3��8L1��z������
��x�N�+�����s�]Ε��/�hv���Ӛ��oSN��6�;���Q�������9���tؼysbo��Ğ<.x�~ �< �6c7
���}��Y&�a�hͯȎ�BfV��
�q������eB�3�&��s��JS�y����_7�n='�GG%Z�ɓ�{�UW��2�K�P.���2*������)I��ÒN�QA>�5Hm����X��x�y�F�!�����b�/& <�Hά���eh�Uk`�l�5���.*����s�s+���T0f7e���v�0�$0Q��Y(2;�'LS�}q�Y5�jE��r�k�L�Lϛ���>��ꩤۙ������0�F�?O��yJU�s;��bN�|]�ʳ�h]ٗ]29/%��LY���
k�j��u�D�Q�=q�O����1�n��b��?������Pdbe�۩���MF�%��}	�,���j�����ƨh�v�?`E5�*y��m2~x���o&Ѱoh����x��&B�����To�wl��m���Qx�>V��ì[����s���Q�|��A�S����JZ�
���>�����LK4'�d�m8�BU�G���#6�W6r2e|+|L?���8�yU���]y�Mo�r�̻�a�g�d�����o����Y�T�N�`�]p���i��~�3ʸ���3��k�׬w���������������������+ �D��9�0;�}����ԛnL������c�%v�l�5���"�=�.=͈j
���h�1�.g�%��]�h�	*�g�X��^�yQ������~��O�2�_ZO~�#L�	�ΝK��So��fW�y5j����܌E;elR��Z���h�������xW�����ؤ�d��f�p�;�ʹ�(���	0�n;F^G�OS�4S.C��S@)��N.�0�����S�2�2,�!��QM��]�	sdiq�z����&Ѱ\^��%h�,��LLm�q��Ժ����S#*�	���`�.�7F�-t����LKj%,nS���fsQ�QgE�k.K���N�~�� ���=KU�󒕯"�L��"�i��I�|��R��|`>KU2P�Q��+�m�����=T��Yiؚ���h0�8�����Ppl�}�L)���ym�a������w��P,W2nL��r�6)�[G�c~;m�\�:��I7�������)�f2�z�`�z�f��=�F*���1M��}^�$���~ήg��0�i����oo�����*U��:��M?�rnF�%���f�
6�R���{C}���g�xޡ-��۔�����ɧK�]F�_@��Ż���W�q�aZE�#l�E���1�?2�7+���c'�/�0��*Rf.W�H�-�|�j�������hzź��h�m��A�H�T5��kf���#�8���A7c�,7YQ,���u����<ω���ᗝ���Vo���w�Q�.�_t��a������N?����~����/e��q�Z��ػ����������������������+ f��a��zF�̝ZM�+w<��6����������Hl'��MO�߮��%���f�b���b\er����Ğ��:|K���'�Q����7�Y���f��S�#}0�p����&��ia&8 ��;���,�O�b,L�6�7m����y-���0�<L��	i�H�m��R�3�E2��yHf�b���?�voƀ�̙t����o�PA<3�F��܉7�7�6���6�x�ybG�5,ا�$�ι9�b\X����,�����q�}=�g�����g<;��}��;VhX�(�I�������-������w��;会��&ߛ��&v�ĮĎD#�R`�g�tA��s��~��}�؇��fc�p��Xa���G���W�<�3h�|Y�d`��R^��i7oxݏ%��Ox��esK��w��_'���$�
ߣ��ӌ�7���z}b��~��ph\���{�*�w���ܓR^0�+��}����^��	�}�^�ةm�L�F���Rb���$�I�(Vm�J�0pV�Ӽi۶�E��oޒ؃������� �ی��G�{�-7'�ęc�m��k�.��o��w/|��{��3zX�r�?􏉝Y��+�X�VZ�sg�۟����x�䧊�ʧ?����s�ԫ�m¸*���!Ӕ5� �o����R.K���!08Ӓ��i0`�-N��eǔԧ[n�|NNN%��~�#w}8���	�|�a��~�4���+��E}X8+�����	��Ș���g�}{D�����Ht]�r;Ō�[v�4�K;Z����C�\��XB�=u�hbo������ ���1��zb'��"FE=]<���fs}�n�בz��<~F��y�����Ξ��??+ھ-h햋���ʀVK�ͦmR�R#�c�����;+�۶mGbGF��ΝǊh���<�`�6�|��仆qG���P���'��a�c|���O;קF�5�k�~�t��3L���_��� 1Qj5Ӹ_�}��N�f�g�w�nk4�}+�Ȉ��1 �oà>�ٗ�~?���\/F�>?�F_��?��3�k��2�/Ep��v� ��:�x��̥nXy���ךn����k�vF�f|�M��3���.��S�:�P�p���̭>v�V���u�w�����L�O'fV�5nl�l��Q9��j�x��mA����\bzX�%hoU��{J�E�iF�12����A���߃_��S°���'O$�,5��h8t�����!������&��g~aE����Bӯ.����s!�n�.7^i�yq���dAo>o!^�n�)w�&FިYz�X__T�{z����v��\p�7G�<�5�OGA�D�q%;z@�oZA�6�c�@�����Ն�Y��������NC���	m��jb���g&v���0f�|��$��w	��ޯ���G�!��e��R��l�n��q�wݙ��ozZb�y�� �61K`�<���H�+�-���慑���T��E��^At�_{�����`Z������}7��y���ub�wޒؙyi�4��諁��3?��r�����9�I��{�	c�G_��Ķ�й��}�A&����ľ�e?�سs�Ɓ�9��{�w=7��\smb��G�#ϱY�^�˼�a�G��}�����Wb����{��bb���ޖg�������;��y����aa0Wet	��_�������;|��n��[���������뉝]&�ʜ����e����G�wH}��W�,��i��ׇ�|Wb���"��)Q�e���n�)������e�}�~0��뽉������n����KO��Uԯ_�y����g��wa�f�_w�&���������J��9NFj����6���Yw��°�+ߘ؅�r�џ</�����7;f_�0� ��i3��x��?���L�[��[{����e�v�0-��u^��g~��{�u7%�ّ�5��~�������zb7o���Y����%�۞zkbk���rI�'H����]������%i7�Qi��L���헿�5����oK�>�������F�X1�q��z�<��OƸa�;�~���s�+���'���c'��U�`G��z���Q�qF&c&�}��nk>�v���Q���}]0�KE��RfN��6������W�(�� �xm@&_&�������cpə|�Cxڅ3��+5�g~�>+��>?Sgm�IOț�g?W|���ons�ӻ�].�TL�~5"�l��(��,������Q֎5֋��k��&6��>������ΰw/TlO^fk��� *�q=_P�����'v �����������������������+ e�xs&0���K%zHq���g\i�MN
C��z���������|�Ď��44"v�&�sj�D��P��ӭ�
3�`f�Lb+в!�drR<�s�	���žk�I��>�˶k�N���������=rB��ǭ5��14.���ɔ �O2܁H˳�f\����i&�d8#���1cn� ��O�f�w&ܓ�>=���_Л��1>Jpyֲ&�a��V�M&�z���>�e���:<!�BևGN	s�!0�Ș�G�d{��X{�M��j�VQQ��z�0ж����>��6�V��TJ�$�
կK��a���P[
��ˣ�tN>.����0g�l�K����i�ǥ���*��[�}���������]�`|��ʿx��'�m�r�M`ʀYy�UU�ڭb��>��r�	9�����J�+^�}������n��������΂���$�s�gq���=�y���m�m���D˰:\+�B�V��ɺ���|���^_�Rр��'?��
���{��=xH���~FH{�$����7� ̨���<o�0Q?y��%ݪ��Z����_I���T��o�)�q�]&��g�{�^a2��'�6���?
c��,�o|Sb_t�s[�g���#̾M;'�rh.
�����'�5/x�\񺩆0W���j`dl�y�g��F��_$����z�0 �~m3�?�����׽�U�=Fm�8"��J�0���>��w�'��;~�pb��=�N잽�h}�wJ=�n�l��Ǥ����#��S���ݳ��C�^��oHlT��1y/���Zy�/��9ߝ�;��z��/���{�#ڜO�F���Џ$�5/&����D[2B�ާ\��Ďդ�����G>"ډcc��"���9<����f�`�-Ή�!�r3��So�%��z���&���w���R�Ȩs4`P�>�ɏ'��w
��~��yl��)��}�0p��=(Ƕ���Yo$k<_M�S�3�0���>�y8��5�o84Q�͸�f��<�g=�m��{.�߾�I���V�R����f�3�.29Y�G�.��k����a�8�{�{��^&e��2���;{L�/5h�^,�&z�2�|7쾗���)���_��}��j�VD}n{��짼�U��N��������Ջ[�ת�wABvzx�nK�/������L���fJ�/՚㌨0$���+����ۅit�3E��Q�}_ͬŃ���-7�G�@ �smF�E�l1��
�JQp���3oӄ�`"��-��D���:a����߅�|�vY(O��%���h��r�Z��Xk夙|췵��/>��`�X/�/J��������<�l.8�weaMЮz��/"�]	d���wL�2�k�+T��|L�A|�^�!�bF���y)��â�����h?嚴��y�<AH�B4Rܷ�I�[�`B3Sj	L�f��>z��𴣏N�Fޫ^���Vc�G{EN8M;�c����F�����> �|_�W�hۮ�JZ��3Ҟ;�P��`Z\�������>rR4},�c[E�m��+���\�rݲC�sR�Z,���4�:*��?�sa�5�v]/��֒�����'x���?���
"�C'�a��a�~���$��h������?���X�U������:۴U�����an^M_���ݟ�Ԗ�¸,A�ԣҿ>����ͷ�}wl��vzF��O}�D]�f׾Ğ�����>��k�I��h���G{+4̞w�0�>�I����
���U��J�0���%�PԂM�����Z�O�Y��o���'��!���4%L��G����G$���|�v��y�zP��B������"����&�[��ۉ]B���â-y�����<W��7� �e�>a�O/J{7��Za�<v<�oxÿJ�HQ�g���,vۈ�����
<6$������L�=-�������
��_��ݿM�������}���W-��e�w��ԋ�}J�6?,̌�OK�C�7F��CK�h�����(�JCҟ=%���?!Z��"�P�X]a�*��ݎ�g���}�k�|%�����~�+HO��җH����ÏՅ}���d�J�Oz@�Tz�m��F!�O���,^_b�U�c=���:1����N�]͈����������s@�Ŋ���f��π���(�A��FQo&_�|l0�O�&V��ٷe��_���M����riyg^���e�mxT�~|}�e g4��o��W�����?�IͤS�w�V/��� �pd����'A�/   ��g��9���V�gv6G猍s�q��m�1��G�;�8�qG6��h́��1�9�u���9�N���S�����+iF�;;��Ǿ+������Z����ZYYYYYYYYYYYYYMby�>�<	�	!�䁡,<��,�K?�����ԙ>s��m�jz�Y�<��׹Y��?����{��ϰ�I9z�9V�Q�`�Ӕl�\ze��Sk "��}@����G����
��W)� �P�gX>ODA<�4�G��`>)�A2�@ͬ����}7��O�-O�ˑ{��R������<���!��I���:]`?EH����Y> ϊ�&dx`z��o�Qq�TSu� _V��|=�|�3F���'�@��N���ì���uOIvX��΁d�;NA��n�M�ÏEV�|H�E��$P��n4�z���(ބ�F%��:��>�|NO���Z��G��P���vuls��߃��iS@������r�!�;��\$$[{;H��4�_��Y�I�d�@�Y�����9_D,�Xz��e�� N��V��k��!���Ϫ��3@��0N�{<Ů��*��X�b�䑮(�3�v3��/~oĖ��G�t8��S�7c��D��)��|<w:��o�=	1LbJ�ͦF������ Γ�r߲cI/�����Vq�J�gW~��T���Mσn��T3��jf��˪��ɑԪk����+\�Bu�2�4⎐l�����s߆�e��'b��݀q��5�o:
Y�ϒEڃ�0�n�w��w�/��n���[Ά�e&��$�Üo�0�������������c�m.�'t� nn�v��Ǣ�$�/E�ϕ�p:�v45�}���]{�J���O�<owޏ�.]"6�_��	��b��<�>���3;z�T|��q�����S�~-��V���,^g{��Ax
�0��]^��@�W���p/��4�@��We�	��tg��d_�����{��g569>o���iq�/�O�lG�xUW���O�J��Uzm��T5�<d�@7�W��;����B�͜0��(��<Yի���y�j�d�/�Vs�����%?�:L*ݿJ±(�H��!���x�Mo=]����ǽϼd�>+++++++++++++++++�I ��O?�6�ӴW��~��ȓO�� �C��X!?�cT�M�o�˯��l�"�]����6�4in8�+�-$=b$�
$p��ʑ��"W������^Yz��N�gS>�a������W�ɽ�������ui��6+A&�Wn��<[�����{����/͗"n��~�^�7�nb1����m�lGrQO���w����r#$W$�_�<3��Px�L?H���X{���,BO����F%�'K��݃= W�@�}�3Ȫ9���~�^_|	Dm�)������Q�fxR}�_�%u�j\���Ϸ�N8�	qg/!@�2�~��#P���3�S�F���E�o��V�ק�ws�� ��l�]�����
��/�5�@�M�7�%��O��)D�Y�M�g>�b�d�@/�������]��_+3Tx��#�^�d���kU��א��C�����4{�	I�6���"�hy$Y��}W���g����b�9z�u�t��i�G�ꫛ�[$��c�}�
d7�։�WG�>��*�t}J� ��z�5�x�[�c9	b2��mq������}� �8_������Q�j���1ګ�Ff��az��p_;��#U<�x��$�U�	z�I��҃s����_U\����<��t���9$���x�y�$��1o����k�q9ԋ�W��<!�w�@r$��Z���ӧ���s<xw�Y���O��@�����{*._�H�_�d�g5ü���Խ���	hmms������9yfa�<��$� f��Y�7��/C�AX�L0�2�l�E�~���x�iz���R����w�y�4e����5&Wʒ|���2�I���ƹ?G]|���빼w�h�H�w�\WeC�,����;~`|�!�ʑ�;J;k����������gn��s�/T�~g��ߡV��TI��>]�=�s�ў��v��ҮRO�r�o�����z�e�>+++++++++++++++++�I������-�}BД?y�)+�|����3��
\��9s6#���V�׭��N/I��xv�.ߤb�^i�� �u.&YI�}1Ǭ�Y�̚�b� ������`E8���=qr�|��8��`�
B��W�;�>�����W�L�ʨ�>_�g�����r|@B�x�+A��U��ŕ����ĘX�I�]M���j��� I�H�D	SGg�/ 7�&嵵�Xm ���)r{�e��8!�Tp�����7��7@`�w��4��F����=��@���?QQ�M&# MR!�7�(���d;�Y���f{q�}����y�! ?�����߁��<�D���7W^��o�ld�
I�g�����~]ųOyt���� BB�7N<�8�8�f��� � ����!����ˌw=�H��1?���·An�y�Y*�����v	zI�C̑iM�&k$kr=�>��W�ȃ0>��N]����Y���!�i�x��u���CQ߯|�'D��oYX/y/��n?�U/]]��ҳ����%�����~Ym�b����q���7�1ٗ�'���Q���I�o���xs�fxܽ��]Ŭކ���k0.���>��H���/^�ל�>{%^�4�>,֜�C�z�����:4�,�i�8/������G?�b�~����i��*W�!I�G�A��orü�9��= ��/\�կ�x�������V��Y�c��^A��"'��0��s0�DS8�+�ѣ�dj몧�)�=��ɣ�S���s��s�Z���6�����D�Iذ[����ob�B�߼������u��ΓdS����d_k�a~����`h�ĭ��ήn�k��ė���U5"�Dr����G����'�<�u��}�T�Y���v������1bV)�7Z2���i<��޿��o�c�2�y>9:~ۙ/k��������`u1i��d�>+++++++++++++++++�I���%�W<�59�A����~@i���Nc� �7�s��i�|z�eA��AH��o�Z�� 
��a�Qɂ(�S���T����$�3��
���9Y��K>��a��Y�����Y���k�+F�����#7�W��I>.�r#dR���A*��&Z&a���=?]y��B!d�3G<~�AP{ё��k!�$:�^��2�l�B~���7��O ��>f�<���V�?��Zc��u|!��Iz������/��w��9�moWqK/�ꖯ���]��.��KT�e������:���cO?��O���_~�'���^}�ߑ� ��1G ko�4ds��^Łț�<��:�����$;z{�������������ݵ�Q�y<�u��
�4=���X|�$�^]����- �sØ7�A�3_���x?'�W�����J�.�/��0�,�|�/�yt�V�ѩ����s�h��
q�r�}]��$�Ys��|m<�g���0K���z{\��x��K ���B��1�=��K��?��L���J�s�m�L� Cz��d�@'���~�j�F�n���*�ش�$ɗ`V�b�}\3��GN��ER�
�6��w��.�y �� ��>��*���4�!�{ѻ1Mo�7Ї����Z?}:<w�lׁ�!�u ������zz�oEz6�p}�~�e*��j���{�U*2��o#ѧIt�wz�%S���V���{ ���K�5z�-���я�(��̳��=���IhvX+K��#a,�2��W�}����Î8B�M7��� ������a�21��|m�����h�������^ 1���x�ʼl^w2ow���)MF՚�(C4[��&*�H�FdS�����#�t����N�G���V�;i���=}���Ԛ�/|�S��+ԫ��sX�z�-��硜��NV�X��2K�YYYYYYYYYYYYYYYYYYM��y�7{��<(��9?֞t��T��t����uT�]�M�x��s�B����<o�X��e�]s�d�4�+��| �Wڵ�����76WR�R�a7ɗ�K�]z���=<+^>����O��r+7�y8�~���eUI�G�<�s#+��^>$���c~��o����	�Ƿ��s�q��d�?�8��>f�-�J%��2d�:A�mݸD�$=��$b�ȶ��AW�#$Lb(��$��>}�{A��$1S�
"Y�$*H!V)��P2�~�����G���;Jť�Ab9�-����3O�ؐ�uؖd��A���z�u���dd��M� H��m�!z\^�ݯ����$�- s��ٝA���3�/<ߒe����ۍ���k�M�n*Ȟ-����(ǅ�b��7��](/���|1�Ϸ1+�p�
�aMFj�&�76���g%ٸ4�b�b���0�D6�5���S��[z���Ñ5�����������h���'M�&��YU��:��Q��+��+؏�v�F���Ah:Z�w(����x/�%/��%��&��w]�^�qT����5>��k1��I���x��Y��۪&��|���oy��/�T{i����z�g��$�aQzk���p~I���Go�8=��?� x�0��l�s�;U��f�Q�/QźF�-�� L�r�I*fخo}t�v̋�,�����HN���$+y� ]C1��j�|���a��p���ɧ�5�u6g��f�z�'!+�����CBHy$��U��=�݉8?����*�z�)*n�@�-[��UO�g��U��d2J+!����x}>�Q��|��x�y��BV^�o@r�)P)�0^�(�Y�YV=Ę�A�vIUK��yG9c����=���lw�r�H>����̵ݨe[(T���?�F{��n���瘁2V\�Qֿ��Fyʍ���	N�	�z�t���1���z���i�+���鯝D {*��a��ԫ�w~�TeίΡ!��`�D�������������������$P��I�~��q�:j�O�\��ociӑ,h���'�����(�4�fZ��+�A��sg�5��/���!IPp?��I�<��a#�ƪ��9s���I��܍ �&|B& �y�\�V������A�ɺ�[G��ҍ��"!@����Λe��� <${j{�tĩ��4H�[o�U�� �W�"��Y��1�=��u ɘC~��?���R- W28^*�qP��aCᨠM�����y�������Tij����������y>����dI�,����?\�b���1��^�-d�b�뮃^����ƖF����L�����?��m+H��&�6�ۺY�"��,�� ���o8�(�v��v���z�8�&����{K�`����X�HpR�дu#d*E�0�d�Y���X|���4���P�$����l�/I�s�J�վ.�����d�v��8e.=Ue`��bL�z�uuw��)����Tܸ�T���M��E\���:���C8B��p����f��8��㏀w�k����PK������L�5�q�n>���`Ę%l{S��{��S�>�b�Ld��<��/�������7���A����ݲ	�����g"��Sާ⢕���kD��}�H"���H���W��G�V��x���g�����������Q�32/���f�&Y�a3<{3��z�Gd7Go�h�^~D*K_cx_����!��v�[@@ǒ�?�y#u{�vlC��_yI�s�>G�d<Q��&R6Z��LYR�e��)"�D(��g�@z�B~��{��ĭgGRi�@���һ�9�$�?I3k�JI��BU:��~F;ƍ�+�U�9_�g����5?�K�kV�*��9^�����}�2�`vF{_����ۼ���x��y�߃�e��Fy~I(G�:mqu�D�������������������$P8l<�.h���ɺR�T���'�Ɠd/HX0ޗr}�ۙ@5*y�����;K���2�\䵔#�|)��.G?���ͩRfVy!Ѡ�ixM���A�y8�C�sd��6O�Ͻ�}�ߐxlx�
���.jrT�RR�_��w�q$$hP�w������/�����֮�s��Pq�˯�����gU8"�W<�A�8$�f4��� �V�����Z��|���j�C6ڻ�{��#�!�i����йȂy+=����e
H�K.�D�5] �n��CO�PD���6Yj���vu�}�\�KV��)�X/^o��y_�>�����	6��Q����VD��x���.P�g�QI��"��g�0�����<�iw�Co�n�P�4�H��z�4�u�β�Y	��2,�
7�Y�(s�O��\�3HB���XFe�ʊ����4n�^O:�]�<|؛���g�WqxD��fI	$�Ɗ�0N��`z�	A9@Ͽdo�믱�<M6:� �%��p�drD<�DcCx]�3�tȏ���+��?oi ��`^��f�N��ge�Kg:	*�K�>�:n�(x!C�6�w���z.����x��<4�E<���^�=�������y��C$f���x&���gR��Ĝ�{aΫ�{@��x�i*>�t��O=��晸��;p^�0�h��Ȃ�j�Jԫ	�����x{ｷ��<�l���6؋����ޢ�ab~��x�n���yںn��Gw��}���ShgP�0��&̪��R�k��1����x9�$dN������R1��T�u8Ћ���9��h(��E"�z�8;9�lYRP<�C#׳�L��$�/��mA/�b}��F+!�|��� ���Uf'g��I'�|�����X�o��{���g�r䍾O;#�=Zy��4��Gl՜���r�����sM ��h�F���7\��o��c���s����3��������S|�����<���ه<4��v�����ƴD�������������������$P8,Yq�Ǟ�2,��t����|<LdE$�ɪd�<���&�WN�W�������n�>���} \�Ѻ�"hx��`����D�]����OA��L��DH�������?��xK	�`��] "z�I������10���}$'�˰��KҰ��]�$�,�eH:��d�I3������UlI�Xy���Z:����:�R�rn~��?�E���&~r'�����~Kŏ�ۇU���@{hO��E]9����P�ڕ�ձ�������uz�R�qf�~@tm�eV�0:"3�vz<�^}��=��X�s7x�t�G~����Y��!�w���H�D��L���x��9�?�w��U�Ӱ��l�oa�a��}��ho}�����4�)%	�O9�n��@��"x�=H�A�=1i��6|�ioUq�4���$��Ql'�Z������r��Tܰ~��Qf��ӳN_�$`z0�2my X�������h��眩b��מ{���o�,?��2k�\�z���$�
<�����������r?�����^d�!���Y*�g��~�}�O8MuHƝ�U�/b<����T|�էU��G���b$y3���܁�}�Y�(̑�;��Zw?�?D/�d3����]�^{�c53$�R�|�� �BE����k���f����:����+@ ;$�Fv�SOc�:����NF=9��Zq��4�]�$]O=;����p<��~}#�,Ǚ�7�,���\ܜY�sy��x^�Cx{�u:��N>I���'��>���z��y�7��q�úV�G��r�'99���?�q��?���<~Ω�'N9�t���:7�_�b�t��L�_�%��g��}��$�m ���.�W�>(d0��Y��̂��Gc�;���T���ע}$��8v7�>�ho����U�6�i���j��G:���r]��a~������|Z�Vx #�g�J��������ڮJU%�7^�g�J�+�����EmI>�r�����^w�+86�Բ���ˬ¿��=Ce�1��{X����h�~�ݣ���Iފ�;Z ��L2�cѭ��9#����,�geeeeeeeeeeeeeeeee5	��A���7��Si%�'V��`d��+hz6�,u�,!P��i�l'%rL^2�P�'��N�G/��fgrw�oAc�N{ΉH�d5IH"A�'�azK���0q�	� ���d#6��^T�yH��|^�K��a&Rb�:dC����O¥�$�p+��az8��l�x2f�n/�A�f���x�	��X�dI��bz-E�m5H�@Q����!$�P��) ��|˟T|��q\b��m7�,��ff���= �(�< �芫�Tq���*���4�F���Q�,�.S- b����%�`E.I���k���+��q��ln܈�&ނ�	0?���6������
R���u�2xF���d2 �$릁P���P񨣎Qq���"I�P���<�z��,��K�q]���݈O��v�)J�Mn�����?���qw;���0��s+���u����#��d�̙ ���8���;$Y�32���Bb�yL��쉧A:�Xb�h��T)����p�"d��>�Y��F��>�ӣ,���7�b;p��Z��	�Pno��g�����]
�o
=������w$��O�%D3���r��q��\�b���%�����ŏU�d�_�>%�!��l����%*� �)��q@�(���I�l����_��"�u��뀽�B���o<�����CҖ����(oh�������HF��$>�l����d�&�͸q���_�}��2�[��;�yIH��) �z��xϾrw󖍬�d�%����&!���ϩ8/\'콯����	�a�_��ϩoB}�l���{�B���e�]�ļ�=�!�mƸ��/c|?z��Y�	D1є��A��~�\����4M�����Pl�����AF��x���y�� t�د'� ������'Jt�Vf���P�y&�/�ע���M��l�yr׿�=��J͓�in��0��\穨�~�̨��#!��q�����Y�����>��_v���q=�/�L�'�������®�����1�gz����������&y��Ĕq����~�l��I!K�YYYYYYYYYYYYYYYYYYM��y<�+HY�C�	I�G�2��k�$���d1T���{=�|H���=�~�ߐ�����R9�\�~��Ò()yV	1�u�oz-z���Eϥ��cHV|��K�q��~�k��izmul��vx��ʺ�xY�3LB)K�eX�
��x�7@$i'��d���H�����c �īQ���&x��r Do��C?��R$����l?I!i�\7!��TH�MϬ`��Xĭ]��+7��!�B>d7���'���IoC!��@��xlG��[y����?m�C�g5��%*�I��:c��ݛA6>�"���b�l��$r��̂J"R��B�J�h2��3���b8�P�^<�zz;޸�& �~�M*fy�s�ra�0��:��ų���Q$�qa̓2�ģ*@O�͝��.��6��0=�$_�n�~����� /(����y^�!w�<�,�?����RB ֵ�z�O�h��-�����H��¸��KN�s�2~��'ƃ��B��L1u��w ��v���Ǩn��?��-���[�iy�w���dߕl�y�B/7�+��y%������;��/H+ɐ��]�sɖ\�,�,oӺ5*�S�4	��6�-�B�7���]��C�nz��cOBT�h+�$I��_���A�R��������9}�,nN�Q�I�9�l����/��"�,�ߺ����x���w6���M��}G<9����#xE�.esb��u4��/d��,q�D�v�=x����y^�y!�y�&Ο���!cx�U��34��>M��oX�Gg�vߥ�>���q7U�[H�0bdb�/�_�YI�+�|�NTa�rv�����9�*��%�ɢ[m1����l�㏷�t�Ӈˎ������7Vү1m���T���7��#|Z�<�t,���s=���E����껻�K���,���t�z{���Z�賲�����������������
'x����#1T�D���s�Z�5�!�L�+�ѧA���k���A7�	�R�^�X�G�>_�y�s3�m>odbOV�IPHv?!���I<�2�@1$]����z��]�����$��'ʐT�e�Iy��@��WH;i'=���W���:��2�t����D�U���Hؐ��/��i�K�x"�u*��z�@�h� ��C�$���ZA�䘵Q�#��e�	��]����t�ai��tB#��W�Wǽ"һ�=���&{���
�'W��d��A!��h�+����r����s�fW;����ǚ��Ҟ�,F7}��;���J=�"BH�
�/����B����2+A�q�Z�h?L���6�Y�EWH.�}xV�$�2��"��`��'��S��K#�i��������{Qg�v�?�W���"�a�6��$	�d��>�=n�F��h�,�v��q���.�����/��.���:�+@@=Y��T�,�A����$�O:!f�Im������l���8�7X���n������BX��O�8��Ӹ����:E"7�iX$��[�+>�Y����gi��d��cϑ~5�S9ф�4�ɉ���=��~�� ��8e�q�j��1}����?v�Sγ�RY���o�o�	��&fr^G��k���B¨�l���1Ͽ���+��	�1޳�8t��V�o{�ue�����C��*������U���`__`rhbL̵����K����*�w�x�k�T,���[�{���C�߼^wc�W���X��O����_+<?(�tXk��}VVVVVVVVVVVVVVVVVV�@��M�N�-/�ek�e�s ��%1�oY�.�է�G
� D��38�G�rx?���[O�ט��~�Y�5Wʬ,��-���Ef�A���(��ps��F]��GV��/i1L���0�x�e�D����F�p<#�M�A�ỈH:��sB�O����
�>��U�b�P��T�
�D=�̾��Ǡ �BTtw ��|������PO��r$>B��b��m���@E��Uw�^��u�'YkD&٣=��O[�e� �*^�0�-� {�GT�l��d}%١d��4�H�����t�n�]�AR9�q kr��g�Y&�h�`�M�9F�����A�V��伈�V��pk�,QF;4�&�G��]a�]'�d�=���P����p��ǅ/9��7�e9�m)^t��Cn�����'/�qM�jT���k�G���&G����a�Z���^��P�H��M���9�O8�$������|��3�,I9��ҍ�M�
�-�9$�t d��6�Y媾j�3A�ɼ%��H�K��X�|��9�WJYO�z������s�y���ٷ_Xo�P�ǣ�e,,^wx_�KVd���S���g K2�嗼��ͨ���qx�>=~"��~^�@�_r|���/�u�G��Az�	5&�v�J�����}��!Y�L������U�|���W,���DV���C���ߓ����#�������@����o��Z�U����9������~�+,���N&���_+�q��n��0��q���S�J=���Y�rd�o���<�,�geeeeeeeeeeeeeeeee5	@�DHT,Y�l�{ת�	`���BK^8���ʶ�����WP�B���`ްp�^z$�~&�"�O�ؑI���$�l�swԿm�5�����G�N�=Mbi�@zmq�>�٫��R�'��:N�9!��:A�� "A����%r�B๗ܼY��=�֦R�=D�Q�; |V4�-T�}l<�E����vn�7_��K�$�`/ț�+���0���*���ב\'Y��`�ɶ���}������^Ə��X0I��U��n2P�	@v���u.��r���B�@�#��y:��ٵ���~}�vțUq�}�Uq�� ��-[���U���fvnC9y�O�f��ǻ�0�Gܶ�T�2�J��I4��Ϙ�4���[��J�f�g���ס�sՑ�,���
��Ae=��C=I���C̊*ޑ~�MW<�"ɨ�}z�r&��D������s�ڍ<>��$�mi^r��� ��ڀ�0D��ǛA����z�) �g\�u��mB����!΋C= ���YW'^��ߡa��f��l�ҽ��3�qp���� ��w��g�o��鮷���~�r�Q��V��7�,�ݝ�^B!���Wk��O��AJ/�,��ǘ��s-�\o]�q�I)z��^�i�F�{���8�Y�?r�U��+�Q1����}4Z���|ߔ������]�����&�:�����
G��ud�V�kxߙ�KJ��{��=fvK	�{���Qr������V剏��[�v�8��*%���*[p`L*yUz�	�NM���Xϗ_�f�j5���g��@歑Q��+_/-�ڛo�c�����.{���1Y+պ8gW�P�����1�����}ڍ���=����)�˱����)K�YYYYYYYYYYYYYYYYYYM����2X�J�H��� R$G���mG7�	:�<5V�̾Z̹W��Y_�=!�$���d�Q��L��k�g�kO���"�]�Yz��y����~_&�hxĔ�����^�����d�-��)$�۬L�|JO��'��#b�*C��ȊQT��~2�ʂF?4�s��D�{�}:"�!�'��x�	�'�V�;K��BNV,�}"�jhh�����S{J�W�[E�&��Ӹ��e�ȕ��u(�mx�i�@!Fy9fI�����7?��O�^fq��G�C��I�E�&�~�*&c Ğ~����T|���`�=T�%�P+X��n�Y�����c�������*n�bP�C�Ds>+^�B2�2��������;X��O8Eş���ؘe���뢋?��� e<t������(O9��V�����Tܸd�]w� ��j�O_�Bl���Tz�}�� ���x]��^x�eǉ�!��(�|_��Ϫ8e
H�����f�aS- ��x�Yhy�1�������b�d�~��GUll�u/���͘_�[A~^vѿ�8w��$�^]�H�;�CŎN�o�z�+C��S��n�}���Uq�O��>���o�����j+Y���]�M���!ǝ��$
��=�7������ẓ�T�Tx} k�㯱�b��_��
�8�,�s!��%<��_�8��;ULA\>��<���s�:�r�����w*6Lmb�t:fv��ʬA�K�_��E�}G�e���e���뱺1�[��J;�c�3H=�n���kE�s�v"���	Oj�$�׵!*�q�����G���M|�iW#7|��1z����^'&�c�}��ɦ�O<�b�$��ٱdu�����3���5Rp����g�7�7����c��[���e�Se�W�Oz�M��[+Y�������������������j��O��
I"IWf�Ӟ7��+��E��`X�����x�=h7�����cA��}�E�*Ƴ}����3V��#/(y���!����+�#��8����A�tw��l��8���N�;��4	B�lIGÛMga�&}"�\tg]"IT���Jȳ��}�?B-FS���o���7����S�	�{�tڵ]��c�܋��L�Ɋ��d�M�;+���E9Ł׻�`�L�5�i�7���'B�d=.�����p��zг�^���Z�����Kb1�8�D�����G��N�����;O�)��b�j	��5�aVۣ>L��9FŮ���}�	�ao?��>�E��ڗUL5�Km��M�AX]��+T�L�j��U*ƛp~�$�*eTwRa�EX�g��˧�?����Cf��l�� �woB�Qn����W�-���p6#��:���)(�5*֑ /��.�_������韠���hs��� ���H���(H��ݦ�0{���T�^��7Lz��/]Ŗze˷`<$����/*���*��w 9S�8ߚ�$)��A���y�����KTL�>���%؍$�0=��������W�v�9�������N����P�7��{�1�;}8�	�a�vb޿�6��sg�S���p��I����?�����&ސ���^�ԏ^���OR�g��b]���[�E���z����M;��k������x�7���^���Y��7��X R�������7*6M���b�js�F|�Y���y�>�{�?�F�&&3�۠��MΓ�v�zӍ�&y�&�|H�q��[N՞o��Y��)�\�E�ҷբd���]�j5���e�X�����?���[�������KUzlV���,vF�.}��|�������!����{J���v���%�������������������&�<�JON�[�D���]��e���\0o�e$(B$a��$�H�����rE��Y33����&���t3I6��Z��f}�l����&�K���J���xdϜ�0�H�� ��y�k*�I�HV�X�1kn(�&��쑥l��o���ګ��^K{ �����}��6������Q0�G�8�$�v���x����8�xo�8�Yf��%q݄����]&�A��c�0��|����dv߭����K�A���ױq��~�)F��=E��Kg�5�1M��� �k�x"$���YS@=���*��W�T�}.��>�M7^�gO:�d��A�[�뿿�U/�"H�w���g7��F�y}^�T�b6�+�t����ګ�^�*ysAz^�op�ɣ���<����'��v�����E�!��cNT1�'1�����I]�d'��B9���?_��k*�>}7���o��l<Ԓ$ߊUz�z,w�mY������O��^�!�.N/��ѻ�ۗ?3�l�W_����/c^����}*���7��Ҍ��p�M<�${q�D�y���L�?�Q��,%�-�e_��@���_�^��s~m������?�я����^��Il��~��Fу=��/����C@�s7ȻbL�j��X���H>�"x��� fc9zЅ@�-�3��>k*��i�*�w�T�~���ȼ��[U����T�{��*��b���-8D���f-�!_x�9= ��裏f<Nſ��O*ֵ5�F#�"������<b&)7I�����*�Y�K���X�4j���[m�)��5ڳ�7�F+�r�q[�����M��^�V]�3>ƍ,�������*�w�$��c°���D�%�������������������&����L��2�@$C�7����e��}n7!���l*��u�hZ�*���違H�k,FO�\�M��_	b'�!M'�Y&��& ��'�����$��"���I�yAzq����U 2$�4!H�1X���5ܗcD�uR\�[<S�1MH]�Q^�
A��3+(���WUǢ�����G,�\�(h3�]DƓ�`���f�Rܺۇ����� ̶n`�K�}B\��c0�&+�`����B�}>� ��H�%R ������5���dq��	~�]�� ���<�V���d\�^��/W�c#�s��G�8�r��W@�
�Eo��ۭ�y'ڌ�Y��(ב���w�x��oRQ<1�1\O���o��2�=��s\�M6�yt{e�b$=�3���4��
x�OS��0�i6�v�ch���x<Y��z{�?-SQ�|?�o�]����*Λ>O���|��/�q����AW;<�͔�*ʐpR���Wq���l;�$dv�rv��@��1��ǽw���KȲܾ;5!��	�<DX�Vs��$ķ���:�$ߔ:��C����_/�7��{s�ܯn�VŁ(�Y׆,���u������T��B�u$IO=$j�^�
����8�����A�]�����NC<��¾����G��v�Q�?�|������^�z��p��k��K�~�oeV�%Ͽ��a~���͝�b�'�O7�Eř�A�����?����}����£���� ��j�VxT����n'�[Av�1�r��Ł��<+��W�7��;�d߮��;fbޒ}�J������ņ��h�筜w�(ĸ0����$�d��D������T��gȯ{F{[/�x���<�Γl?Q�Sw��dG�}VVVVVVVVVVVVVVVVVV�@�}Bj�œ� �xT���,�����f'O�����X�$Y.�áWSn�@k
^d��fs���w�F�M�n�3CR&3�(��xߙ+�E�7���z�7>��@ �C���� #���r�~��c!S�NUQ�����%�ӶNdo��GS$AB��8�CO�"H�x*��f6`g�/�����~�?j�Ol��ފ;������1���!H�A���p���n^(B&��/�+���<	М\/\)�I9!���#WL����g��U�ymf[�����د 2kl�4D���T��?��g���qg�E�W^_���5  }�a9��u�'�߯b{
^h瞆��y�����lk'��� �:����Q����ZŐ\�$=��7�u*�ca��}�؇�%��y��c.�H�X�|[Ƞ������ �o��/~�,�/-~A����͒8f����*�h~�r0��u�E�kBf�Z�J�V�ݍr�kd��^�2l��Y)�v�6d��3lݬ,�/ q��� >��Y�����/T�7�AŃ�BM'!���,������Y��h���s���7�����YwS!�O�7���.��}+���V��,|V�#�e��V���oG��x�Ȣ|�g��h����^�B�q<�����D���
y�6ޔ�=����o�u`�{���Rq�l�{�7oF�8Άr ��:�1�x��sо�5:���=�<�ݣC���Q��]r��<����7��͏���D�瘱P�8N�^#��}��Gn��$������������o� �WL��1W~�;�6��d��󗇀�г��E�]���u|�����@�0r�c&�ʐu~+�YΣN^*��r<�R��XU�<�w����Xe�>+++++++++++++++++�I σ>�I���3+�x���P�t���<Pw�>�ѱ+�QQf�MD@0qġ*� dB	������1m��Ͽ
2e�
x�^��V.�q�;Y�bŌ'Ђ`��l�a�'���{o�&x��H�
 '�l��G�P8�0dML��z���<��R�م�fz��U�πʓ0����L�hO�%k��ǲ+�?�D�@���D�$�|k�&�j� ��g%�x-Y��$���L3.V�w�;Kqn$�ì��(H�	�°d����k 95fuX0=�DYp�u�.��,�ܽ�o?���>��0���i���`�m�(ȣ{w���h��L?�����*��@L�?^�"�����w䁘7��;��b�Q0���S����R���y����,����T��?杞N\���gU�m���a�2n�a�>�c��"�)!��0.��]M�O�^g�W�R񤣎W���vq��S����6`�7�0����D�{����O���,ۯӛO�� �?�Yj����8��Ѕ����O�Fw���7��[��9;��J�e��c� ䷻�t���ȃ*�v���B����)����}��L��}���}@ųN����u��w�s����yZ��9	����������ev�ԓ���E?&��M�8���������9����z��&�~EI��q���O�x�;��W<�֭^��G.F��8����wؿ��6�s[ȼL ��}�}���0>�<�z�q<~��v�$�^y�`Q��8���8�C���;�篵	�x�Jܶ�]�dzk���z��<*D_�&=��C�WJ�UzX��v-0d��~���S�~N������	��%ۢ������o͏c�]#Rf���j�Q����\�u^�tP�n���JͿ�;G���v>���3�w������G�9���w�V;O�賲��������������������Ŗz>��JdX�x_����xZ��)$y���,��Y�~8�@��Ka��g�$	I��H��h��b�[����.92�A$�U�����1�|��˓t��Z=�ҽ�Ҋ��ʒ�;��oS�������0�d
	�F/�>��r�3�%�\��/w�@�5�X�y�`7�K6ձ��Q����8Rx�v&��'�~�3ߊ�h�Dc�W3��m1��2�>�`d�d�T���^Bt�kY��`�f����U|�51�_{E�3�@V�"ѤǟE6ѭ��J�dVYo�|�&U�V-8��1~gΚ��/����_�9%+�y�		�D��晘��Z���A��ۄ���d��w*H�Sނ~{��GTL�Eq>r$�r��������,-����!f�N�q�$�3�n�0[p��;��Q��]�庩��7^�/z��;�Ԝ�u|�A���H�����6�V��*Oc�Ƙ���W#��y���1��X��Adk��"K�d�MM�~��Ev� B!02ѧI6�߉S���P��:I��r|F%[�4G��Оn���!�!��<�4WB��{�F\/)���a{!��я���'U�N��n�࿩����L�tc�O��w�R�����Hn��o� �1X@�߸�k��&8�h�D�X޶B1��3�����d��7��1~�����y]�d^�t�O�� 3i����y=<��Z�$��U�f�h�4�5�$`������]���֕(��dk����9��xtl������x�S��c���I��&^Hܛ_��E�ʎ糹gE\����j�'c�r�V�T��p2����}e�;�:ȇ���Qyl�O<>w�K��,��q]�~t*{[H��#�v�v6h;^`f����w�x�uV�����h�Qiy�����K�U{�߻��C��m�s��e�>+++++++++++++++++�I�p��1���n�B�+��RO�M
��W��{�v�]'Y�$��9�T�ԃ8(����c,H�"I� � �I��zAH�E�Z�^\
B*CrG���a�!ɢJ;�'�B,���#�4��=�x-RG�@�\�l��azy�Xh �ұ��<��6 �(=�~;�e�W�R񅥋Q���,�H�M� �,�Z�o�K����W�Ү����u�sm�XSy��W.B���K��}R���y���a��s�]�1�t?���M��w=�6nD�׽��˵��{���+?���v�����R���2��r��ø=���ULIJ�h��)fe��9e��0Ȳ~f���]��W(�zl쀷��7ޠ�e������{�qf��b��]��0+o8���!��H޿�>d5��|c7��ߺ_ˌ{��$[n��G�����nz��A(�q�)*N�Rj8����{A�v0� OD�DY��o���*>��-����T�=o�@�o��[*N�9]�%+AD�_V1�l����܊yzpp��r;�����^x��}���x�Y�G��L�S����kP�c���C�D��k��ܬ�T���d���!=�o�y�Eo�a��r_h�����=w��rH�sĘE;E}�{�~�l\��0���>	�MH�!�S�BP�u�i2M��U֪��~�O>��������0��2+}�@�IP�W�Fx@�M�g^6#�����(���Z�O^���u$^S1����կ#+��ǝ�b�d�^����w�Ws��FH�n�����?L� �������7W�����������t�W
VJ���U�����h��$�ܛ�L@`�����,��%��,�]Y�N���|�w��_M5����>��8��cɩ�UŞ�Օ�Tz�VI�v���U�z��j畀��D�������������������$PɣO/T�#Q���=xW�}yYY�~|?�!�b�R�Q�� �E/�}f����C��H6ZAa$Kc���d�"Q7�
�r�q��+�K׭PQ�Պ�Z��eR��@f�c%%�v9�}�DHI��N=]���L^�[��#y7D/%y0.ف�BXlɰ�Y�$�q�Ŷ0{b(v�/� 	I¦�'�E�����ZH�P���~���]��[�t�]2.�Xq\f�@��� ԊFֹI���J}S$�����f��qݤS2��9�G��Y8u�͕z}!0�_BWt�z{z�����'A4��<�:YN�P��̎�\��� ���Ux����T|�ŗT\���\��k���zlhd�bA贷&b��].0�����$���(3bg?�3Ib,�Y:���H~�!�6��)3�t����[����Eh�)'���� [�Y_׮�<������m�����T�e�WW�p��� ��;o��v��2�pS��;Y�O��{@|��8`�r�r�BA<���P���)���޴�����L�w^2��t�_oD�Ą���yg������1��Ӂ�x�O_�#<��(�6���~L�:z�]��*.ZL���9�Dx���x��7�R1ĉ��?�v#�I_u��*ַ��zI�q�I0+o�Yf���%$d#�{���U<�$�gf5�<�9>�|�i��!;���糉ބ�-8{����򡇮�-SQަ��kV�D?� ds.��_�"�+T@���xO�y^_Y�q.�S���A\Ӧ�=�6�����ۢgs|�)�T-�����X�^����B�Ǐ8�M�.בQ�K	��
�?/G�ֻ����(� �e=zt��s�גG����<^���?o��{'��T([!i�1��Ʀ�=��8N���>�"{v��'�!���j��Z��U���ר�����&j?Ԭ|��G& ����"b��k���/���])�8Ye�>+++++++++++++++++�I ��W 	T�ޓ�YF���:;���(f��:x��5g����A�Շ@j����s L��Sh�6dQ̒�J�ܡ,�t>�=�4D��E��+@�#�4�J�~�ʽ�P�o)6<C���E{b E��!b���Ж- c��@ ��(OV��� \�@":���U z���KT�I��B�8�x&�D�=і�*!5e?�ǟx��D�b?ڥ�J�(*]i3
7Y��*3:y|�|)<�V�^��vF�!z#F�����T�8��� #��*�X�\sfÃ�{�Rq�Y?�"�HI�]�.I^ʸ&HUd6L�J��h>+o'��#��K��|�������c@��?�eSg����@��Db'��us�>�;���T���(-�BY�im zn�r;�R�����ً�!7!,Y�����^d�$�����\���pmMa���t�<�����⾇�b���0��x=�I�e�Y�G)$p��Ax��I�ƛ�~��U|�ч�����G��+@>o�CVh&9}�bxB��y_���I%r�<�?r|��p^?lx��~4�C�Z̟�_��̙�T\��n*���}:�~N%b�7���fW޸�XO�a����/<��HL1[��՘��ʼ��iʉ�Q�A��۳a*��y�!7w��;��������n�R�����ߦ����b#��U�p�<��y����̏�@*Nm�癍2?Jb�kW����7�C��o~W�.zi�X�G/�g��R<c
��NoA�s1=f�rx_<�Px������]7�x�]�m� m�g|ѨR�W���ZΏ�+�_(t��>�q�?>����x��޳�L� ��Ƥ�(�Y� �2�aо暰����v�����ն�8�v���;���v9��1�Cl�H�`�EO�XU-�]6�m����k���*�W�8�:[��� ���#K�YYYYYYYYYYYYYYYYYYM�}��\�YW剨��qE������G��4�W\�t����tȂ��z �s� к��Tq���Y{��~:���dDK3�C�m�t =�0�2�'Ƞ5$-2���ޚ�ӞS��Jڗ�l�|?�E=��cv�DM ��{�͔ ��n=ȭ��=� ,X��lf݌�a�%@T$I����k6���IdK�>�N�k:W���[|?��S�<�/��PyMrO�}|M�.HT����578�q$�r�p��=�DͶx�EI ��(���\�ol��V������T\��\0���Y!�"-vo�O���S�/�$��~��X8��]}��T�׋�U��D���A���w�U1OOȩ�� ����	��b[�#��/�F97��oc7��H�d�b$�1��sk�q��g���c�A�P�v2VgA4:�h�3�1��f����$��1>�|ކ�� )���[��_���h#���+A��@��3f�`o(R-������_��5�{��[v/���YZ%{w6CR8�>�r��ۛu��!;��$� ��[�u<ʎ
�yCx�)�u���͞�b�L�b� ��W�,R�g�����zf�7"��2E��|]׎q���k��Y�������09��W�������U<�(�h����i0���ܪ���C�T;Ƚ��F��.���G��~��x�m.�!`~ش	㦷$�������7�_��p ��<ɼ��=�q���WT<hO�j�_�+�ܾ�h�{�����:�3恠|�T�sd�}w�����y����a����7*.Z��׷�+���=���3͉uC'�͆)��C�� �eez��W�5(Co��1N�t�<�Y���/ۻIVH��[�j��_'����ņY�x>��:Xq���J�x��9?�?�7�.������+�5I��D��s��R��@�����O���|^��+�|Ox�q��x�wy���v
r�6���~�7y�;Զ�v�,�geeeeeeeeeeeeeeeee5	T���K�U��&z�vae>��6e��J�a��3Q/�fW��Y��J5	�4(���^˓�i��}"Ϥ,�<Q]����Y�$H�pd�1o>B�� ��"fA�h��`���d��1��H�0��%5E/>���~
�81f%��8ӧ�ؘ�
�� P�|-ڰ��!��ű�a]`�2�I�H����ƒ�;����#{��Z�OTf���P ����H��.���<A���q��Yf���Kr�:d��5y�Yg��#B7Do�x����S��qܥx��l��=�t��3_P��{A�<��#؀䓌Sw{�j�"�N3��Wq�ܜ;
�4G�MH���R0�[����i ��x�*���$Z$�$�(���yדw���G���:+7Ɍ0b�>�z-�
ư}�����r��}�:�ɮ��#�b�.hxT��h���B��[�ل}�U��H�~����O��J�^���+�-�`��}�v��OB�	�������|յ#�!���
h2խ�J�~��+�lG(��,Yr��o\��.��	�����y��_�^q�MS�Y�k�Y��A�E�EY_b�8��b��?�_I�?�M)w9,6�������o�_ �-GBm�R\w�љ����WϽ"��- t�z3���{���u�u3H�p��1{���uu�C�Jc�x=��,��V�zOȇ�{Lŧ_A�a��-s@�7���_��]}��U��i/�/.E�^���H�����<s�v��l���@�� ��}��Q>�b?���hO� Y����
exEL��,� �˒pQ���3	`�{ɼЄ,4Ⱦb���*�>O�]Tc^q���5����sÃ5��}k_�Ǒc�o��[�y\���.Br��&.�Q)	U��U8�*T���������!�G�Ыu�ݲ?=�1��-~�~ڃ|�H�J�UK�UJf����9��g����>V��N��|9�Rb�8n�$���w�%�������������������&��>y�*Q��0	<y�;}��Xi�)�����1�c����@�����g��I�Ɋ~z�͜7�U�^ ���%���p� �D��s���R�,��i���Td>�@L�]�O�M�QG#��̙��B�T���'�)���`I&]���+'��?I�导�b���I���DK��h�=��}0�[Q�����$"ۦ������A�6����<W�sNA��-$����o�عc�2���@��L�wb��V(�q�[ae3R���s�(�w�ϝ���o9�U�Dȭ��B�`㭿���gA��Ih�t$��^|��7vO)۴\Ǽ��<+5&Ab��托�\,8�?I0�� �	c	!I�������Co|�I�b�M��8�!?/H�40�mI�'J��$�8Ϻ?���|oI��c�&ɧ�!�@��2�<�~W���8��ĳL��E��&�������MPJ���դL�M��I*�AP0�li���^�<�'�oL��:#	w��?I^r[X�~���x��G�>\�9�o����.��ߧ?�*~�_Q1D�� ��Ν�n�S]]���֬���$�z�vu�3�i&;! IF��y�٫׮[��P^����@�q�~q�s*�p�CA!fIj�{����,���Fd����X,��} �#qfO������!YRm�l=d\��������]H�IO��������=����7g��}w�0;�w3����~��h�D��k�s�*�5�b�ёO��n����#Y=�0Ğ�<��������t���6�r��������Q�#�Z_��4����^e(��y#o?�d�>+++++++++++++++++�I�7}#���Ҵ�@�g� ���ʲ<)�3w���V�{��/�L��sT񠊐�
kB�d�ۢxsq�;Hҧ��`=��XOԻ��Á�ᑴ���Xn.P�"�Ɠ'��8B��>a�����y�$z�vcg'�d2�:nHH�h�<}Qzf2��m��~��ܴ�ŁG���(?O�X�ȤQ�\���e�;�
����?�,9�0�+H"���6��)H����c�$ʍ�Q��0a�C�a��~zW��ْ3�7�rI�|��q^֭\�b}�eK�M�O���T��_�Wq	�+��\�}�D�����`vU�`�-v#�3oڼ���&N˓�r��7�c�wo�خ��J�������ۻ��BS�����qa���x)�,Bn��� r<�����Ia� �kfe�_V_y��$M�(�(h�l�g�nǃ�έIJ����.������kَ��齧���4I�J���>�� Q%��@X}QsXD�0Ͽ�^��k3Av_p��U��5W�8u���r���<�᪥KU/�p��#��B��Yf�N��<�pޒ�}c#��V���|Dp&�R�2��lg�B6h^W�l�t��*�s���w�*�gv�����$��O�^c<�1Ƚ�w�i��u������Fr�뿲]��O�U,��c�o%?h|o{����d'�i¶�ٵ�K������`R�lvN�q�D���rkܲd��r���;�Ro��<L�$o`L���Wt/�=g��͗;z��_l?�-��/Ռ_XI�D�������������������$P�}az+�_��gz,�3�u���̑xc�ڧ�Iw�aG���W_	�PU�fA�e��E�af�eE�z��[;�9T$��k�T|�U]�*��I(�����_��hHI(,#>���[�D܌f}>B0�&����@gy��Bf��۶��z�;���)�A �]��	��A��ᐐ���M�yR?2�W���y�v�Q���o�7	&Y�c$���U��UxF�|��Hŋ#%�V��$����NfM�����n��O}RŇ�@�͛6��"�R�Է����@�tw���ԑ�1:�����g��^�p%4L��v��s�fW9ޅcjϩ�I>]�����\���X0I>�z�^w�f%�8��cÂ� /q�J����'^�:;�	����g�2/[�8��k�#�G��\�N��O�(�l���7���c��g%��|����"j�_����d���c>��c~��kW�������Řw�H��Y��|��1Ϭ_��$��"�O��n�<��e����Yw�i��$�#��x��I�;a?<�x���F~�����Bd��.d�o����󸸿����מ߁��f=M��g���̕d��F��{E�$�������u�F�x��;ae���x����x�C`��+�/MT���	��7��d��h���)�]�H>�{�*Ra���)��Y����ĸ^˪���x{���_��^\��|��g���}Qu��2��|<�j�{�d�׋�2�Z5�;�E؇0�|O3���d�>+++++++++++++++++�I����+�/�q:�+��ĻI�'yb�ޫ+��x�ǫc��@�H������r0Մ��!y�p,_�w
�����Z��] ��@��ͺ�!���JIy�A�ߐ,�y�7F/�'�A�C��G/�X�3DR+�,�u$�z�m8��cJV`�K�65c�g�C6յk�`�(������~���[#7����iF��}Y�TG�؍��y����~��gw��2�
�?i��R�j�?�[@HF�Z��^z��7�<.�1W�u+��[7b|i 6$��jB�}�7�q���>�橸G;�N�0�I��$gL�gU<
�%�vg3�g.�(㡡ޔ�ݝ�PW,���P��k�����^	�o��*���]�&Hd�EH���+0�z,x�4��:�y�dfu�5�.�l�q͇�pdޔfyV����M�>_N9��#��As���LF=�I���h�܏�Iva��xW���IB���|ڝ���N���'��������9�~�.FB:���ݏ�(ٻ���u� �f�9_�	��e	����=ԏ����=H3�N,^�� �r$�d��M���y�Z��K*
�'Y���T�i�fzd��`���m�����p䍉�~?�f}�=^{�$�	ɝg4<)!��'۩{��S�컣��kOl�/�d��z�x��;���vB�G���xy���dgT`���D!9�Ʀ��|���WK&&��U�OU}��;�_�{�ƪ5�W�����I�ƪq��S�3�G�m�������ݟ{��0U��6ȷ�Y~}�Wwܪ�r�:8qg�Z�}VVVVVVVVVVVVVVVVVV�@�}|b"Q,��9�x�\�K��?���<����C*�
���n@��H �R�$U� ���G���e�Od��GV�?܌,��mRq ҡm�Ts�L`{����O��v]= ��a�} �{�;﬷�8�l�Sg�o�����2K��gHJj�De�Yo{6��~E��_w��X�1N�'�G)�DJ���kAVrF�5!�9#?/���&|�C	y����f�<>��1h��q���xѻ߫�V]���#;n�&�c�:����;�O9��͟�bg'H��S@��ګ*.Y/��)��������*����uɒlɽ�166�1�1=				!��{)�o޼�p/��%�0c0�F�7Y�,ٲ$�������g��g��3{��]�ѱ�~���Y�f͚5����ߓ�u�W��(QV����*���i�/������ӂ8>��3 6�#��$I���zY?�]���zrYg�,dWX/D�
��Sl�ݨ?zܣ�c�8�0v�v��h2����թk�5W��szٺ�!�!'�3�`ؿ�|(�WZ�����I|��>:?�ߌ?G�k�9�x�L�Ll��ъ�r��b���)��
�Ԁ�{�P���xJҎ�Y�������~�r3�c�# ��D��q�����.Z��}�ݘ $_qd%��S��9��&�أ�H^�9"��ǭ~Y����T^:oz�6�h�Wy1N"��q3BX�k�P�xKJ�YH���}r�@6���p�)�wTSKI�,�q� �W�=м����\�����{�n%&jZ.8Y����*���ƝP�=Z%��q�����3�X��Q;�^w�g�n���8Ϳ�m`[��y�n�;N��`��	���k�;G�999999999999999999�D�g�4�y�}��dn-g|3�T�z������]ۑw����<��(���T�2Q"�&�jD �z�Y*��G?��;@D5�D4�A���H(�AH0����ͳͳ�۩�!W,���e�����? ��_v9�H�"��ÔݰZ5�Y�2T^����[���=[�~�k����A�!��eb�A��a�. ��z՛m���Ye���L��zG�+�So�b(Ȫ��I���C��OY�O;�T���T|�GU\�l��앵v�����F7o�l�Ǻ5 <��^Ļ��z��\���;��U��;ߡ��X��z��q�ܿ�!���q^�Z�7��f����G���rZ�?2C6����87	B2���5�$��0<�5�L�p�0�kD<e�T��j�H���׃qi��[?GY��ATq6���UZSc�*�t&Y��pLk;M�q�m�g��zF={P�Z��3�<N>H^����q:_&fi;9�;E.?h�L�y[K ˚�O���Fϧ�#t}}򜣆a�/�������,�3	ȣ*��eo��)���"��	"�ׯ7�*���#�1��yr����e����+Gσ��u��]A�;]׽;����T�=�|�N�	>��6!a+oD�yd?���B5r���/1E��Zܞ�N�8����RR�	ɾ�*[?�~1����ܒ����&�;��-��kDóM�{�z�:�R9���_hA�"�$�H���Qk�gt����*7�%Yk�y�[�g����)G�999999999999999999:�E��Y����@���h}�����7& dy�fn��m*n�ﺗ_�b��C���)���� ΂�x�{OŹȄe�kPE� `�,��E��g��0Z	�b� Ț2���@�}�_S��;�T���N�|
�)9A$�cf�ʖzǭ?Sq�~y'�8�Q��I�!>y����N�X)P���L�5$��=|�X$O?��f�m~�s��B���Ũ� i�#H1}�\�E�`��2˫n|���=O�Vq�ȽCc���U�Rq�c�U<a�:�(}b;�_�H�u��	��;w��G�J"^�����Xg�K�^S�O���oc�� D9K6πd(�3�<L�D�7�ҕ�,�������r7&L��G�c��\�
��u��*>��U��8������T��Y[���͢����:O;���~�WcȞ���@Ż@���!Y�4���n��+_��*���Tdo��Sn��M*�w?Hўa"�$���D��Ƹ��w���_�"�g�>e6���a�F���R���_U��q��D�m�r�����=V����I�g@��i�z��/W����x� �cz�������*�g�>�Y\�=w戌~r?��b������_��KT\C����0U'���s(�B'�z㉨?�������W�yh/G&�ȓ��nW�x.�)+�	�NR��@�OA���Q���b#��תt!S�)��5��,��
�l�@|�컖��ŉ������3�ӺL���z����E&9ts�>�n��y�DȾ�$_rr�\��ob� �f��y6��_Tx����/?B�,P�i��Yb��K��'�g�
ɟ�9=��]�����.�K⵽_�|�F9�4���v�Ǎ�>'''''''''''''''''��@�}�&����a�<�x�Z�}D8���J9"�); {0U�vN�P������R���=6[�&2����{Ǳ_aTe�� &�W�[��g}�h�B�gr��nCx.q��t���jxuM��D#�}gA��ߣ޽}���x(�Z�����ɳ�@dba ��s����s�m�=�<�ު�P~&R�	LΞ�׏g�5ᦳHRx�ɂ�[�����e���5�S��f���L`\�{d���o�ӧ,��F��^Dβ*������C �^����'�p�
�z�Y6
��A��I"�z�z����u �n��*2����~�r׮Qq�����{���upY�= ���I��[�����jJ:�lS��q�d� ?L�M`<y��/V�_�[*Τ@��~׏U,���g�r�����_T�C��P�G#9�W��s*N�P΃£�M'c����������3�3�G���5*^}	��]��ٖ�,�+����~���8"�� ²t���X�֏S���_���GOS�� ��������ګF��p/�������^�����'�c��W�8�����q�嘇�:5�8�p��w���Nw�|��Y�i�Y�0���mv�� eS/�	��AܿU���>}�v�O����7��7=��ף��Ӈ�����W�}�^���eT�aY���p^{�z�P�}��/�z�8NO?yђ�#�'l�� ���Hή˞����Y��WI���; <;d�}����I���x�l�KU�ē jb���	;���aE�~1�V�$_��W���g�D=ƒ����YUC���q�r�%&S��u�X2��wl��N�yq+��oһ?��~����u�>^�!9�F~1b�#���������������������}:y!g�����S���f ����<��6	�R(�� Ȏ�C��,��E73
��'��t�*�<H��2�'��W�l�U�7~�I'�'�A�6�IE�"��M��>Y���S�C�@hLyS�i�����_4ʙc��QV�7�ذA3A5�V�L��<��O�2Σ^Cl4�y���
D(�g�D�(g�#3S)��H>ތ���#�h� �E/�)��
��v��ȤB�E�Yy��&oH�fd�4n���aHb���!K�k/y�uH��� "��.P��Ƚ�_x���
�����w��n9�gx�ӝ[~�b�HV��c�4K�gm�j�}5��!��Q��c�e	o�c=�4�'-7ȣ�W^�9�����R��-W""���/��b7�	w�O~��o�ᯩ8;����}TTd�
c�{/ȯ_��*>� H��ƻ�\r��sg���ZE�Ⱥk^�J���Z/�Ǿ��N�N��=�s��oy#H��^
��4�z����N��8Y����e��ؗ��w�nU�_���g�s��o����l��s�9�o�n'r��r���zs��G�[�\C��D�i�QΚ���"}?����bO��y�"�������o]ű��Uܴr����w�}w�����C��/���yD����������k��]3E�gp^��w��4��k&��D~sV�|�����L"����;���F0��Q\y"�k��v��(K\���ɒP��d�-7�����x'ɾ��ǣ*0��y��eWʉ%Ļl%ۼ��:�HN��������$_�D���-�{~����%	=���$��%�{r|h�<[X���]/�K�t�^]/���\��;3Z	��N�\���Ad?���:.��R�#���������������������}�+��>" 2D��$=��aY�<�^���# �jD"U�@L�7��0��*y�͔A4T��y1i�Ǌ�����s�!*�ߐ��jz�x�-�m	gz5�)�Ρ3�T�F��a7˗�se"��8N��F�K���\�Z��)�g�Cd��Y8���`{�-�/�x#�3SLը�Q|�/�����B�w�;CY��}3�MH�Z^�"��kȆ�����|�5�{��y�q3�3�8S�;�@��[��,���yF�����;��կ|E��Qx�R͵���u�i��x��&s?f�t�nW��ˏ�g2�:G^\���ϴ���7��>�d�FO�,ym��F��Z�O�~6�o7����[�5R����x������}����O-�	�y�&O9	����-3�H��O��u޶ٙO��^z�KT���H�D��lE=�a��2߿}��W�_��e����d@$��~��W���|�d��V�U���] &�6��zOA�����b��e�?�l�7c���U8���ˇ��'"{�0���]��<�"�$k�Q%O���<5�K�O�@����#��ك�A<?���*����_�2x$�i\��W�Uw���X!O���߫�я���g�v��7~�[TOT0_D=������)�7gQ����m���ЃX�`={�.'���l?����834��W`,�g#��*PD��U�	�n�1���묱���{�|}��s\�ԳZ��&��E�	
�$D�D���:'�<�N8�ȈN�]�E�-�}��!⼘r#dR*n���#����c6�W���6ˏ�R�V��JP.�qc��m�.��Ok{F���YV�~��,�z���{�$�#��������������������E_���L���2�E���{�ьq��}"�BO0�L�N���z�߲b/m�����,U��� ez�h�YYi���C�笹>�pc��c����Q+iGM;08B�� �|ΪX#���ȴZ�F��GH�j���'a�'o����*�  ��#�Z-U���R�F=�M�$�[�&�ֶ'&�4Q@$��E�嵣 ��* �L��*����} S�D*�z(;o��\#�ʤ
�t�!�0"���xW]y���_r��L�Gb�D^�D��&�o�������p~uΦ[&.��~�y��޿����e	��9����*P�i�I�p*���6�flqF6a��n�pYw�U;ׇ~����KڀIR�S����S{U%9����T���v�T��{�V��/�i�Vދ��m�x���T<�t��}�?T��?"��3@ ��u?��O=�X!������<y���xe�}�5�ʛ.�|�鿾��+^���a���#O#2�kZ���8�����3cT��<n�~,�^�݉������O@}
)�ߨ��3N���K.~��c��ۇ�7�u
U�Ώ�� @��yXzޑG�[��U�4�n�s�X^�Z�=���Gf�~�^�E"�<"(o��f��نs9J;O�� ��O����;ߏY���Yvy=�[�+A�MO�>Om}���lƨϪ7P�������dmW��]����� f�T�goˮ+%	?�%1�=p���޸|���ll�ŉ�4�>� ��������qdB4۩� �}�����<��[*?��
!�ĉ����k�x]���k�>��"i�-���.J
�?LlǷ�#Ǒ�!��-0�߶��i�=��K�b�b�����,�A�����	,����H�>!��gG�999999999999999999
_�1	A���2q���R�W���D2͂,����~�H�\�&�jD��L�G�T:�{fv��ȴbts� �z٣�<��D��NGdFa���̀��o����Ҽ,fB�#�H���B:i�f_x5IR*���A�m�6{�Q��2���W�Ző^�<b�Ї�W�u��m�����~�	������Y8rdzj\�lDHeD\o/H�36���N�T��p�Y��B��$����d�,�i�D#�K����vÿ��iک�6�L}�#z�\!C˴9q"CÊ��^[su�$C��dN91I����}��kPG�g�L[�D�(QZ�=SȂ��S=
T�l�0��Ny��# sjD�.����5��t��q�Wc�2��β$��\kS��㈳,�S�D�ڼ'l�&���p�D(f�̪�t��?IY��;D�E�X�o�".��o<q�q��a�OY�ԟ ����zv�v/��7[�};�^��G��6҃�^y��戠�ϯ}	�݁= ��d��+�~����K�"O���<��L�S��&}�(����x�Yk��A�"��ѕ+T�?	B�yȝ�����z��'��6d�ݺ��W��*��[���,x\f�t�}W]Č�1�+&��,�3{w��l���|��w�[���?�x4����m8�矦��`H�C�ƌ�nڌ��mwܪb��GF�E��!/�l�y�B�z��\����~\����T1ߋ�.����G�D��Y�?��f]ϒ(t�x�������a�NIgޙ���hp�u^L�7��1="Y�����M�����T'�f�h���\{Ps������&������
,��L��N<��^J�6l��g�өګW�����!Q�p��;�B�~���d#mz���ߍ)�|�$~��.�ٟ�F<˻�����ً���:} ��1�0�}-�2��>�Z�4~F���J��!n���Ԟ���£Q��Ƕ�;>������w��О�)''''''''''''''''''�g��/���#�A{;�K&Ԉ��6P���wU�#��y�1�t�]�R��c��x��]���r_��WU��:� �ox�[Uܵ�He)�첗�X�,�Y�,����u�P��Ƿ�y��X� �̵�Ï��6���� y�$�{�as�֛���>"?�=З���}��|�֭W�u'��9�B����@��u�]��ȼ,k��?�@�'v�T��Ԯ=�A��J���ݸ.�]z����kU��;������i��Y�vI�w<s!�bF��̙�^�̚��y�"O;�����d/3��DQ�V���o�� ����8����e"Q��|o�%�TF��,�+�Kp���xf�H����!�\�)��֨x����G�N:�d�+@؅�s�y�|�΋Ē!�\@�1�(g�ji���_��1QL��qt��<�a#Th�@dd.���	�8_p�*��@�=���W��,�D��E��}��>4����y���|6����i�F;������?��T�{ �n��O�8�@?���xx�k�Sq��u8��5{����z] �]x��U��my�I�>"Y�d�Z���ׅ=�GA�Ua:2���o��o��7��n��{��/��RW���Ӏ�~5�X(��<2Gޤy��L&��Dw����g��V\u��7��y��#�q��Y����,�Deh�,p=�){8��M߿��ob;� �3��DnօW�Ž� !�z$�ԑ�tB��@�+���7ӳP�2�ې�mq��ޮ9A+�?&u��T�q$,��'����-�s���3?��X'�\��|�)�Q>��Jm�K�b&ڣ��s�lѤE�|?�����Ħ\����8�� r���DŲ���_4���(O��t}��?��/|�Y�O�䋜��������k~&&Ql�nw@�y
h%
�m�T�D�uτ۵W�V�x.4�b-?�I�����(�K랟�P�_�M�:/�G]��ؽy���%���9�͚�P��ކ�}�S��'�'��g��q��@0��q�Ļ�UI�Ʈ��؃|���]c�69��������������������8PF�{�MFψ��70c� /��4H����ߥ�����6p��g�x�k6���O��8�d�\�d���A�=B�_�eúU��,�m+ sDL��@��Ѵo?b>���{)�w<��r��p��b��8�,{#Ѣ|OoV��jy
$�o����q5��{�˧?�)g�kj��ֻ~ۿ�-oQ�_��*>ND��>�Qo"����7����T���U�l?em�윏�ʁ�yީ����O�x�c�X,��z�8:qȰe�R�#@�-߈,��*�7�1�>9s�DW�l09�J��_�j����`��+H>��8m�hV�<���������c{�u�7�v�L���4�j���H�f��y���D8+teٜ�#��A��-w��lp���?��O����7�d�9�ӨG�)��!I�D_�~ҏg,�%B�X�[���K���g��ΞrX��9��)'�~�u"�}z����ߪ���Ҏ���s�woR�W�s��S��cw�z�3��i���F}�>O=�q*CY�����>������35|�����U<0O�ek��5M�W_�rst�� _�2{�\��A���~��gm>Oſ��ߩ�w|o��+�6S�y�L��e�z�q�����b�doʓȻ�=9��_�C��f�*��7����k(�/�^~�t/Փ��(��=�D�����[���$�,�s�/���r��Mه�<H��4��57�s:�-��wp�T��U��ˣܲ�J��g���eigr+W�~��)k2�g���T���q<NHbOng!�"�lq<�I���8".�V�[��
6-?$�%�oWr�	��,4�z�JĐ��q_��b�yyb��y%A@/hޮ��y ��C���h�=� �+onz
�h;-��_�{@�C'e�+nn'��)�y�%���"t�����(���d.�6y�j6�F�8�n5:,�������`������|l;l�J-mu�lMܰ����Q��,�r��J��I ��K:%���絵��^zR.���Z���vo���i;E��uH��
�=�����i�#���������������������}�͠���e3���\s������*�OYe˔p3o�G��|��y"3 AR�_Ͼ=O)B�+��T&��7�"�������7��w����� ���@����d�ܷ�8�Л�f�rf�I�jD�p<�zr 8n��*���T�D�3���s� w��aԃI.��b8 �h�*"�(�d	���a�F�U$��KЮG��n��'T /0�R��Z�<㨜�P����ՠ���A�^�v�
���r��2�@y�:�T����<�b�<��SO[�W��]��K0M�1��7��\+K�)�= U����MS�Fy:�^d�'0b�H��q\�>"(=NrIYB+���JD��ZI}�-s�>�G��v�y;�������IJD�"idzB��	˕ـm�}r�Dzl��gB#h$�RѦ�>��ϳ+^2�MWc;�_�O|���Jܗ�
�#gɾ�!xp2�w�i��_�>y�1�6��u�Y�S5p���[�~�j;q������A5� M��?�#g���S6r�?gfA���?���Y�6K�X�C:y#��#�Ο����	�z�y�!��G�Ԉ0��f%H¼O��k���_p.<����g��A�|�[*��0�#���t�h��O���rO"��;�C۷R{��N@a��kׁ���w�OA��뎟;3���x�^�������'�D�7EΆ;G7x+f�����W�}�橃c�?s�x�ɩ�S"Y*Dz�|d�f���s���0��$�:�oB�$)9�ޅr �젳���"`� �$��=�<�S�^ZR������L?�$�fB\=1�Y  /a3�;��l\���ހA��)�x�a�²�
ګ�L{CJ�M�'�S:4w��K��!�l^���E>,�2򼍐}fy��!�{�وP��P��	�*��d�Z����sNd?��ej����H��~���B������������Dm�����0�%�VL(f�N�����u�٦x/�n��q�gۯ�l�!9��}mK{ۮb~IaݠS?[����~�GpD�������������������q ��'���>�fu�	`�f�2xQ�? O������ї���)÷�𨌃`X�
d�@��������{��7��=|^#����Vj 5ԙ%�l���CV`�>�����2"@N� ��-�^�3���l�m-eD�b��)�z�=�4�z۞�W���:͐�M��;x;����A:?�8c� ���	"fҔ�3K�{��L��)��� �^��W���O�����vx�=��|�Q�<��t߇���F�F�6K���$�l5��^+T^@ٔ�D�	8���W�^�i"C��}���|hƟ��T	��ė�]�Gw<�8��F(��*�pu&��gq]�E�I����Lx�5;B��ȡ4m������ݗ�'�5UA57b���uJe�
�~��d�Mqq��|^�3�N�w���e9�q"����} �����% ��x�����T\6��a�P�yX	;C�q;� �{�&}W_��<��׿�jOY��R�/�����cOế���A�f߾�;*֩CrV[�LMMQV��o* ��^s|��D?�j��;��#O�e�1��λޣ��!�o��-�3r����koy����Կ�����嗁�d����}:����s�ۘ4	�i�}���l��@p˝����s���Q��k_��_�%HƓ�߈�]��]|�T����buǿ�y���"���!��][��86�q�-o�E:ȯ~��*N=���s���>��sU|�ixl:"�o9��{������;x��3>Bdi���I��d3�r"Q�GһƳ��/Y�y��4�X�|��ۼ�b��h������QC�P�ݵ9�c��YE��d��l���42����=���!�h��ͯS`��ynD�p��5��F�E�V�_��}����::�H��RKL{��3j���z�����bG��X�9���/}���>Ѧw\��$�V� c���&>^��BB�.\�|}b2��ܔo�H������]���,ǝf�<�_��I�M������{��.氎�srrrrrrrrrrrrrrrrr:z�Qd2���1%�&�� ����Ld]��,a�֭S�I��H�W\�c�� 0�:�4xm^r�B�#��:|^�]�H������ټ	Y$׬�l�{�r��f|�Mk&��~� �~�ߡ�.~��kOڀ���$΃<���^R�=r���̬���=툜K��V��+�����2x�}�}��8�$��g�(y�9 ���H�l���
;9	������G�z-_nԏɾF��:
�)��3	}���q=��2�96�̲���3�H�[�y3k��p}$�4���W�9��g��-Կu"3�p]�+�2ykMM��Z�r-���g�ST�ח��1H͸��'�^{�Q9��s��� ��0o&%}]�eƦE�y�D��Z ��e+���nÉ*^�}sD��D���u d_�Y[�@v����Ȗ�����7~��*n؄r_q���^�kȇ��|?~��~"��{<N�w��t�ʫ�Az�� ϲ��Q�}�n���Uܱ���'�x|�83;C�SV���t	3�W�
Y{R���(�y/a�͛nTq�)�B=}�����8؏�ϋ>=r�a�&]�}���jP&�����x'�F%���ΐw�K��B�U� ���������/}��*�z���q8q�q�	����.<'��}x��z��q�+_��p�9x~�i�\�����?�3���!�����r���hz�4�\�S}�����,���f��tm�2c�@՞CXf�y�uW{���3�U�h|�|�Ω��g���b��H�I�����O]���>һ�8|����+�aiaM�
3�X�>K����U�'VǑ>O�-��I���{C�$N2/�Xu�A��G��lA�:S��sן���؞=��Rl��#��s�v�Ž���o�$c";r����cӟ�q�x����g�q�C���F����B�%��K�k��b����嗘7��D�5����wD�������������������q��E�~�o���Y��)�P��(�a��q����nȯ�=r��C�O� ��������M�믆G�C�aŞlU&�����V�,�D��@Tԉ0;<R#M�U?fFC~�0cy�MP��?��?��ó�����u�����=��3A�|�&>[�!ґO�	���*�"9�_&�e����h��*H���}*�𑏩x-�D�����`��:|�<�ry&�p<��cϚ�	d��4�ǿ�go:��Y�w�|�S��X���~N���c�O�8קA���u �~�]�D=�|�
E�_�h�"�#2Qz�i�Qg
,�nCh�{ j/���N��9"Y��r�	�%�|��˱S���-W�)�d�\/�D�D�g����l	d�w�Y�!ʚ<<��,���8���di&���$e���P�5�O������/�D�֯Wq�v�����*��km�ܯO�W^�H�4{�eq��8�o��M�r.G^�L�j��=�r���z+�ނC��E�=��)���,��=D�W��>���}ݵ��ܼn�f���(�ѝ�P�����S3yE�\�`�b��{;�����%���r�=w�8>O�[~�,ױ�7���/��e*�{*H��a<Ǟ8����Vx~����� Bz����s�|��S�5�2_�l�O��u���t�k�d�Ll�w�&ϴG+�?����x!'赥��L:�k=�p���-�m��8�yg���D����o���,Wg��x������Oqҫ����= �P�a�uy�_�y7�s{%% �ǣ������N\��̺�@��Ӟ�����y_ő|:k|B/�xB���×��N��h�ȊV�G���.�=��Z�`f�R��V��V#�>��w���e~��[$4wWM�����E��>���Z}^�q3��Z��Wwy<XpүU�/�v�������Y���h��"y]&7O��wD�������������������q��^��A��x����b��9]��X�����M�՗_�b_�$�V�WgO:�{t������T��J�g/<�OLtLM�P��Y�����k�5K����⬫3e({�<m�w䍭F*�?�D�7�L��W�<?��O�840��>�b�����~����Ud"�Gw����[��O�f<����C����ǐ%�DY\���!��Dŷ��T�}<��ɘ�,�� �*u�)�*H��'��g�z/e��i�I7��jܜD;<��9\���:0o��5�LS�[&-�e�Wuq�	kP������p|$�3���9��$�t���u=�G3S�,�~���<�Ѷ��5"Ryy�x�=MYX9Ig��H>�N�EH�E���	'T"DM���9,e��r�P��ҸF�&S�Z�����촽��o��9�C�����3��$,{f��#���A��}�: �g"E�� ő�C j~�Eq�/�:��0�>���/��7R�����~Bǁҽ���3�����A��;�b��a�,��g�|s���C�$M����$Ʒ�n�:ί���{��{T��!x%�b��2lWo�z~���T�+_����'�!zn0�7C�df���AJ����o��}�?���"�;ׇ�P�Q�q�@�?�Ğ&�H[��A��WI6YH�7��o�8�<��jbK�����$��q��Č3��t��y����"�%1���I�KB����������>��q�]ٟ���$C49L�^/˵�z��Q���~�%I�/&��hNN,Uu�s+���Բn.�b�3K������q����T~�D���(��O¯��Y,�s�o�w�߫��Z�Wvî��߅�2��SId�m�����~�x���M�[��V%�EA�?<�*� G�999999999999999999ʄ/�n1�3оI�1)��~yH]x2��.[Rob$Շ>�u+@Z��Wގ�0"EG���Ir�mߧ�X�/���\�����تPy3 ��Uȃ�8���T|d<��5�D� B�Y������ːuqv��]��I������Q?���7���[�*n�O�۶��)O�e��	hJ�2�.�s�X #>enq��bhh�pk6!{��]��z� ��g?	���� �p>%��*!S qz
�+��B�S��>4�&��Y�t6=��Aǚ���Պx`]~�e*~�?>����|u$_�G����*����'�|c2��].O^��~։���p��� p*�C#8��?Cga|�F��E����l����aOI&*xy�)�[���,��ggQ�� e�6�[	���gěI�1��-�L�s/+�Š=�s�]��زN�ڊ�e�G�%g
i|ʒ�h��=��MfRM"����a���J�q~8'��z� � ����������<�V����j���j�w{��ĝ�*&�>g������Z��xS��f������^��]Lx��}ï�k�VET�r���'�N4�,��^�S3���W'W�Fy<0'g}���{���57�<W�h��x\��yR�L�k�Yޟ|���bg^e���%���3���8bsAb�d[U4�=�Ā�O˶�� E>�o"ǳZ�q!�w���ͻO,3Q֮{�Y@�H���3�U(?�y&�_13�����x"����&�w��mn���@�Ci 	�%�9�)�Y��6���л���;.G��l�K��["jۃ/���hY\+�g{^�Hs�3����,=�����;{nD����_0Y�{���6[`b/~�Ԃ�V�N�o�}���s������m"}�뎖�z�rD�������������������q�ѧ���4�~�I9 ���V�8�ܕW�l[=O5���s���aq�#Ȗx�K_���H�F��-����nT�3OW�SNE}
x79MG�+q��6�����F);�k�C�ǡax'��#xnՙ ��W�љ]�,��r�^���W!���g����>�)��Ŗ���K_��,y�}���`"u&'@*�^ ��s֮Y��@Ȣ
6<���vIS:�b?�_��W���q"?r�߫�ۿ�[XOfX�"��O=#O����^D�0��/�Q����^`a���Wӟ�4�W��;ߍv:�")�>�b���n�:�=�Կ������~�O�V���DFN��c�2Ecd�{��*n�����u�0��τ���+M�Y�w����a/.>o�URY�?���߷c[�y\t1ei=i��+@}�Ư���m0�%Ɓ����I�@D�hZȌHA앗�@2ۣ'A5�����_`zF���:Gނ�j����`�υ�o��ѭ*��w�Ǳ��l��^��O���{2�*P?#�UW�$��3On�y`����g������lqS�"˹����Se|;AΠ�&���v��K�\���6I�k^�&h��=%.<ۂFӭm�-��J

���������ϡ�U�к"��V/>�=j]k  ��IDATW��k5LL��T�_�7�\�%��cB7B,5� �>��}ލ��I�^��?���s^��c�1q�^�ҫ��A�z�יts�(���%�`��C-{W�q$R`����j�b���KJ.����(��޹`����#n���/�m�^��%�"��mJ����<Ox�@�o�<,�胾K�uI�q9�.+�G^���V�������8��?⚭M"�����y[�#���������������������}z�ߜ��/N9�&���+����W_z��?��˨<��ȸ�7|�T|x+����>YE�.��K��:��������S���*�< ���"H�'�ޡ�?w��7nTq�J�_%��_>�I�g�����Lϥ�hQO�c�@v����_z���y=����۷�O>��h��?|HE��Z�d�/��}�F@�1A��^���T���]7=�,Wi򺚫�X��C����^ &�/�y󏾣�)瀔��2\�C�Ȃ[%b�/�v.Wp��+P�C���X�Cc��yv���v-�b�L6wt��!R��a�������u*^}%<O_w6��k~ٚ��3���	�|H˩)x�=��Ct8 6�����C*��b\�A����m{���=��Gk5� #�/`�3ʦ�7B�U<נ��=�-�%­w�߼�ע|�
ۓC�V�.���`Ĥ.�� X�'z�̌̀�x�D��R�+lXH��~�>��qx\�~m��nLB�U�2��J� �Ӽ|�F��7Kޟ��=�D9*�^��/4�f1�Z�	~	nE$��`j^&�zj^�~��L� ��:��H�wڍ��������	��\f��ld��$�5�&+�	Z�|�O�noM�3qHd����u���	�����cY�hz�e�:�\oN~0��H��ԓ�P�ė��\q��~�ɾ�Ǘ�^d9-���8[���z�Z%�Z&#���jwթwߢ�e�l�ǋ�6�5{�z��%����r��j���nI1�D^����f��<�����U��pR8�m��_,����~����A{��8�6���㐒�� �w�IJt�/θ�����f�f���b�>'''''''''''''''''��@G�蓤���I7z�GY�y�nw=��̓A��J��ٽw�8KiG��S���:��W�z�ɦV�ݷR�~��GT̥Ad�L�\��F���v��)��	�� ��f@n��w_�:g����K5{���s/��������/~��T, ��z�^?��O�ػY3�V.�<�?��G^t�C��;2���\��k��i��O��X�-w�NSV��G� O~�ӿ��'�r� ��� <�RCtޘ�l��#�e�0ڵF��P�[�?ϼi��g�|ݱT�_�����_}���V�ߡ��ι �w���'Q����^Ұ�53�i�0�F&2y3kq���f��t��ߣ K�g��Vl�:��B���=�(z>Ŕ R��
y9���G��R{�5G�)[p.��5�P�YU��5:c!H=�g�7sj" ��VI|�a�t J\�O4t�aH7�
ܜ|�q2h(E֙��J I�Z�r�:c���wS��3�����a�uԤL��_�g�b�9�EI�c7����ymq�z��cI�e��ZY�ᄷ��[P�.ȫ(�ek_�v<��rS��=���1܍H>�<��͓��V��t-��p��p��|���$��H~�v������r~I=�� k�|� �"|"۲���٢-}�専Fy��^�EK��q��*x��oұ�z�2��Pd�b�4]�/h�`�o�����iz<����_�Q��&��k���z�$c~ٓ�\-�ԩZ���/�,�[��ЋN�=�b}��c������01ɛ�/��_Z$;\��b�#�L����������������������t(c}�g͙W�R��#l9H�ɹ�H�Z�ȼa�כ��Y�Ⱦ[���tZ��y&G$Y�R%��>��Tt�)�}):�=�ë�gd{��yV�i�^+z"W��L�IfǬժ�w�J��.S�{nG�$Z��
5�=�>xu2ec�N�o�$[����([g���$�rm�����G���l��/�)�ai�ak���7���*���<���v���ׂx��u�dQ��� ���yTQn&�r˳hoz�|&���s�9��`�ȵ�<z�6�=���+��NG����[�D�����LX��׊e�ߧ�9ԟ���Q��6���4���*D2�́�,��<3�"E�7U�e%n4�~U����k���������Cd`�<�2Y�3���z�Sx����ao� �$�!�J�?��]L�Ȭ�rf<���'�್\�&Z�҉�j�|^��:[.m�����v�9�ǳ y��Қ��y���5p$�h���}g�ѡw�u��w-�l2������!�՘w;=����3��񢇕�ؼ��is�kR�Ԣ�F�IB�?Y��q�-{,��㾾���wf���	�e%�[�S�$�$�g1�\����-�G/���Jd��e�(Ց�g݀���K�	����-�v�~�D#D�Ԃ*9��DI>R�������@�c��ӻ�=s���v<�u�����~�6��jyI4_L\���p��S��ݸ�È#��������������������E=��7gU�q66����\?�O�}�n�i�,g�o�9�l������/��:</�*y���ɲ�iEf�"?�6��x�?g����}O_�y��e��'�C$V��-�����aW"rrl�y�MM�S.H3�I�VϬ�W_��ٓ�Wóo��\-q���c����=*��Zi�G����wx?��ddՈ�����d2��_qxd$_��H�z�ϑ7��0<������3�V��H���Qd5�r8�B�5M�"Bs)��'\�+/�L�I��c2���/���^���#����� �q���� GFA<f�d҃��s���({��眥�Q��Gef
�=�^Llz���̠��ڰ�/&Y�L�6'���+��^v��fu��KIrO���mn����T�����.��K3G]�����	"_���9jC�WX�,��YH�����c������b�Ǥ/�����ibf�!��&�.$n��2w��596��y����#<Gm����0{��MM^��ձ{���z��6��0����yE�,��K{�6?~$[��3�u��՞|��$ȵV�%[G�I���^�x�dE���{�,6�>KN}�KVt��'�'�fm�6~w�-2��q�/Jh�mo#��H���:T�^1�?���x֢�Dv�9gv�Ȯ�_&t��� ��Yy��	�_>W�[~���M����.�^q$�����e��Ab���!����?8�b���#���������������������}RE�)�3�43۠�t���
���g�+���3�TN�L��8ȥ�� ָX&����f�u�#R���j/A��4O�M��+�@���ą����������e&������8+�&I>n�*y�U��|�U@Fj�>zѝ�%���r	�v{q�tdca�#f��e�K{h���i*�d�/M�{��ʕ��R������8| d_H�8e"��^Y�����*��V���\�D�#�#�wt�B�e�+_����SOUq�4���yթ�3)X� ���4ʧ�Q�4�8�����8�)�`����W��zT�<ܴd^�������z=���>���ի�z�=��X�@,�k�%�K��3��Iz�b2�����c'l�[�#Ē�1\����(˗^S��-�5Xx܉l���'�D��8�\�:�c�q�%���R!���:����J�����Z���Og�E�R/���	��œ�m#�.����x��rL{H3b�&?p�3��j��ds���A�y�L({������E�;t}-�;.ˮ��8��6J�x�v23��gއ����%�"�)�G�i�Ȅ$B����g��TW��l��&���8��v���2����^؍��r\�l�E��Lb�����E��Z�l�T�HV�N	���T��}��^�Z�ry�V=�b��Ā{��N�^�I�o��_���+����e��U217K9��������������������8PԣO�dZ&ػ�=?�{ۈ���g��6�Df(��.������䑣����_��X��YF�GK��K��xӫ�-Q�iOs�	�4e��3̽��Z��n�P�i�/�	"��݉|�oΌq��<�f(;���$U�ȿ���ؘ���������(����o�Z���#]@�?��ϩ8��y�!��=88�����ݗ���q��l7WC�;����ЪQ����܇�)�e�_��A�>L��׏��ܜ#�ăc8~.��[F�z+W�P;��~�^����OÁ�>3D���Ѓ�O�$L��L�f<��X��^�F�I�e~�%���`�P/7�B��0X���+���kN.�"�6�K�;��~��H������^&/f}s6�F�Uc���f�<fJ8S�u4r	�S?7�LJZD<Ә���ܡ�C&�$�!��yi"x~�G�U\��^�LF���[�����I=��}�&�ɶ+�K�1�ޥ�Iîw����u���7�v/F�4�w��SB��S�S/����p>��o�y*��N����͋ϚM�o��I?a{#-��W�X{^����G��@�io�e���L%$�,�Wd�v�׺�)-R5"�/�j}��n�7]//�t�m���X/<�5#�l3;pǲ�@&n;�����rX��mh����P�1,)F�㿿�:�%7�~�f9G�999999999999999999�/�dV~3���z��g�.-k�g�){�x#���!�¤���Tg���GwL�5L�}~�"���<G�"���_��e�_+��{����C�D���4�>����zzA�1a��(�'\XQ&Q��`/g=.�`c2���:y�I��@Yo���$l����_q��9���nl׏����[�ޅؾ؃��U��\!O���+����l�ފ����"H��}DΠ��a3�0g��%��Y��	�֣�
y)R=�����D ֈT��w������ρ`ܰa��_|��y�?�0�"y��p}��`&���e��'�/��f7���$\�jN���S \ܙ�0[�m擷k4_�x��ĲI����V)�����:�֥�^�^�����'&h3y�X<��x�/��d�lgo�3�Z�X�̼�)�5q%��EV�F�fn&fn����3���N�����/�R�}��)�K�@�L�--+21����<�?4�iЮw_�{��\n� �TC�'�.�z�����㭏�<L��k�<�wG�r��K���^���r�W/.)�Ԉ�ny���[�J��{�{�,o�i��R���'&�x{����o�ݭ�M,�����������Jڍ�k�K������i�γ�v���-�����N��$_��	��c�Oڽ�߽�}����2�w��7C�tI��]�K	�:����y<�����P��x嵶\��srrrrrrrrrrrrrrrrr:fݍv憚�&c3���W��d�*�N�^V�@�����3X��PGV�W�&e�e]��$J���x2�g"YE-30�N�P��>�T�A75/�"�8nHhJ/%A��/��9\�kר89�l��#�D�}CD�e(�k/��L���m���f�Po�x��Y$��e���y"�<ꗯ"+.g���0e"��S��ÉU�(�%b.2Q�d�A:�"�G�����ɫ��Wj �g$u�_�,�Zްa���7mR�L�u��ًQ���\G�^k���$%l�$�H���ۈ�ؙ4�n]&�4��3(��M��:�g�L����"��zA�%W��r�yu,�'߾��b�����ՠ������$鼔�/�^���-�D�$o���k!P#�a��g���p댯 �c��4�o���6@$H2VF���8��e�I�C�=d�W��ˋv�/������r?I�2n\�����L��q�ͳ��^��y�*ɧ���g�қ�}ì�-����_Դ�`��Lu����b�0���4�m��m�V;������dOt�v�H����J>�;������K`a��`�ʓ�{�7��&�L�O�yɶ���+���|G�y"�o�G�_R����/v2��#]��.3��Y�����AP5����̴ڷ�����#��������������������e�$�9c�x��xG��M%����,��A�9� ���������mCX��f��L�Vos�5������������  �+Χ�������B�P	���oԚ��쩔����H��x��z&�8K/�||�\o�W���݁={�����fA�e)�p&��z����}��K�V�퐧7�2��>�?g�M��Ӕ�k3L�'ɸl������ccU\�Yv�o\�r�C�^G���<�'_{��E���)1]���X,��ڣ��w$�cni���S6RJxT�2�G�w�6���,�n��)�n^�kʒ5:u5?�!Ǐ���l!a3CfAb4Q#��.�����X�
R5,��[�ٵ�
�&����!yXk�2��<K�����zŐ7]�QO*�}R�;�����L���|z�ٳ�&m'��7�ߩ�h<)�R?�V������3b��CO��#�Ky��ק�����g�]��i�F���d�;�x �Y{�%H:�	I�8�o��2.�x֩��'�%\%$���9�}u�=�����O���>��]m=N�_�{��Q)��ڡdN��R��t���ټ��VxG��������~��T�������,}�go����/��O�������{T�}5>��6�RP�b0fqD�������������������q�H�ݤ�x	��d�����f��ov%����ˏ5�D�ֿ���y����8"��	ۛq�E��09&�^�͂4��t�M���t�E���jU�y���Ӈ�ղ�}�=��Ï=���yͭX�V�#��-�L�s�ۑ�3��!�0��R��>��"y��M�R}�C��op��x�̏���Y��f��8K���}���~�7_���mUq�nd.�J�������<HYy{{�<t��*����=�����De��'%4_�C���b46�+=�$I&	@�X��$Rj^���M�z��] ��<1�R"��mX�Y��zAd���~��-��e
<��d�;�����H�YD��j��Ö�!�l���(��$���\Pc9�*���<K�e�N���?K���~	�k�Ta%���h�z����OĢ�~h�ڋ�eC���OE{4,Ϲh�7���	<o��#�Ȧ�%it8~�.W~��/��d��-B�-t,��O�Ⱦ�&B�0��A��ĥ2L{�ַ��j7m�{��&�~T��7�)?�y���=��}{�|��1���k�Y����Z�d_����-��V�_%�;�lQ�����ҿ��IG�d������_�QN��<"{��T�u�����%�u0Y���9:^�sKpv]�Z���8��������������������8P&�"0f���^U�l��&���:��̖'�(�K9�_�W��������	�;�M�E-����a�Y��~L�P{�W^@75qDEΆ[�����!�y{&�x�AyL�M�c��?���7����GYu�D��f�T�ԛ�l�����QN�`f�e���ب�P����yN����������k�����?������=�D��}Ά��O�]GF�	X%b�T�P{�vذH��O�30<����)S杫=��U��i��s����&2�	�L�+O��,5y��q�`��L��4��gzSƲ��^j~�uu6���)>&bgve6rau�e/����W�X��R�C���(�t���~xG��zm8�Dx�n�<xx�$�g!�4PfY��Y۷�Y"3�]7�%;UؕDı�,�J��eo��ɑ�$�l��N#i��i���p{
1$VēVd��"ϗ5�[�����&��y�-�q�[$^��i���e-���\U�˃���@�m^��~�D���o��n�G�8��5bN<�߻]#�lǷ���H�w��to���'&?�Ԟп��-���&�ϫbE�>Ȃ�[^�/W���k������������M��@�����r=���uE�y�ר]��}���Ҍ��srrrrrrrrrrrrrrrrr:�賐x�S/|����&.����E��d�䌮|���rB%ƻ r �̴4_��g+�KY#%(��t禦��%:�0>�fb/�j�Py�e��͹�]�0[/T�ߢ3��Yw� *͚���rx���LS�����1���1�e�_������y��+DΕJ�T/":�ك��x�Q��� �.z�T|t�c*����+�W�V���_���)���e&�*K�A�_OeI�������krjΨo4k_�k.��yf�HI&��zڷ�4��b�I8�t�'r�#�=:��}���iZ>{��ꘉ	�&����xʒ�C&"r�*���C���;i?�̘�`��I����Z_��W��o?e�>��,G�|i/�'�T;=G�����	�y
zv��~�>�:S��BT[��0��q�T?�}7�\��Ϻk;�6�4��K��~�䖍 l�[k+Q���y;D&���!	/�C-(���6r��|���l��I���8I��.�׋F�-2X�H���-�s�mR��@>qmύ���)ah�]�h�����G�u�<�;�m�oS~���&߼��,�E�򗙭>��U��e~�Uq}���ߚ�X5���}��@��;g�
�&X1��7�&O?�]p��+��w�ޏ5�$Pv����>'''''''''''''''''��@]{��А�,�lBE3�������(N�墓�&$L�t,��j�h7�g����ä�g% �{�2sO�L�S����
�b>��
��z��Èt㬾�Isd�e����r|�]�7�SG&TdϾ*�{���$!f6g����D��P??�?[�qfg�&}�H�w��-t &�^s���r���y�r����^�bb��`�_ ��2ޫAhe>��s9�ZׅA/��՗߼?�	Gj/��|��l�֨�vN���F�ޘ�`�Sg��������4�j:�3��4���<��$������<�7��4]W�����:Lދ3ST.��I�w;�A��v���93E�;]��>�����v��~��>Iž�34 ����T�G��K�Y��ֶ���$o4��������ⅲ�3�!<�,48خb���^H���n{�%��kS�!�Z���Ǌ�n��aqzΒɶ�%uz>��-��f��R�y�L�ŕ�@��yt��������w--����y��Y�3�>��~��&�[��QwK��y��yN
�`�z�1B��[3�o�<�R���V��f����~=�3U���o�3*>v�C*�?�K����싁����}NNNNNNNNNNNNNNNNNNǁ�/�d6�ng�
K.�71�(frBIԇ�x6l�:�{���&V��I��Rh�k��$�3և3Q�DL�̊K�C�;q���C�5�	)&�Ӌ�wo�KD2��#�:&�)�oO?�����xJg���/ϖTd�,�ˁ\�TK�=e�%��g�A&�F�/W������+T\3��3�>L�����������r
�Y��M����O�d_�gR����������S�T�D�4��i=��[�)J�n�l��2�{�ۙ�Gj�>"�z�y��NdF����)\�J	��و��1Q�L�1$�!�Ҭ�=ޞ�1ӌ��.��c�L�t�a}͙>�hd�Q$$������U�D��]~��׿�z�)�Go
��)x�-��ׂr��|*���}R�p6h"h�{5�|��x��8~E��?)��$ԡwϒS�p}����	l~��:q�����w�C�U�/��Ku�:���>��C2-�ˎڲ�ڷo��ӄ�� !)�r�ɼ���eo���}���L��7zX�Ea�Ⱦ�(������Y\ɾ�6�e<i����/�����Iɼ�ݱ��M��X��V�g�}ek>���}M��!�9��H_<�s��WZ�R.C��}��� ��,�{���!��!n���z<�������srrrrrrrrrrrrrrrrr:K��[��
I;�A�%3�M<�3�L���'�M&R�ǔ��<���/�Öm2�?�.�Ʉ/��7��lU��mĢ.�$�r�p���~��ɻ����6�x㜦7�u�<D�u�coj|\�lo��|b򋕣��*���>����Rq��{v�g�5���F��T�8X���߾�i|�o�ٲ����l��%A��	�D�y�>1sǄ_N��T� ����e�>��J��2�Vx���Y��BA��bW�<�bĨ��3{��,����d�M�31e��+�I���ك1���s�S�[_t+�ې�_��'-W�t�Dh���zW�?��y�O`JܿA�QH�L�����s *'�sAe2����e�<!��Ëo��M���׭_�������*A
��Y�5�cɚ�b�����K�h���9��.Y���K^\w	��W��%����K�i���|Ӥ�߁qY��p�
[�綊y��F���|���~ol/�n��m��%=^��2ՙZ,��|]�L��.�}��좑}�wx��ƫ���_0b��p�V��N�ض�ng����-*�{+՞<��FV[>�f��D�tM	/��ǋpGy��v��}3<o�t��~�_F~)I�[���
�^�8�_Lf�'X��hy��WG�999999999999999999�b�]s�E�y�i�U��eϭ��}��>o���$v��	����V�8�z�W�"[d�B����Lz5�I���j��U<����q�7�K�ii{��+�[��!��|pd�vo>3��]6��o�n3��*���}%�v� &H��=���Y�:���2�GD{��{zTd�+��y2����d@3#H3M"�$)�i��\4���O�!�2*�g�|s^��O�{�M����e��Y8���󅟥���,��t�)�5���F��y��'�_�����0iD#5���u����9�t�
8I��V���?nbHg�f ڹD�WĔI,����9�
ˏ?����w�X/�y�p^�ː���Z��*���<r�]��ϻ��*��}�Ak�Yr�"d�yC��a�7�[�I(''C]F!g�e-R��}��zf.���^B���d}��?L�l��}3m~O�xD����e�}�Q��T~/�+�߾ɊT=�=�����8k��/��
"���{����h�DW�=-$S��G���n��j��|V�s~���"�����om�F��_��[%Qmp���/L�Uje*��x��78���K�y�?�u��e�e����{%<������#���������������������z��1o�;�V�̬2��^}�8����'�0ɋ�W�t�/Gm@���l��l�CM��6����7���]˿���7�]"fpld�e9,�$��"��G{��e��Yo����7��V�7ݳ�yO_/���4�����?�H$����ǭӛ�0�l�z�����G=��?r�LΠxfd�����z3� 2��T�gjdE�u����1�#�o�'����S?\Ωؾ�f0���f��zx���~L�Uκ�D"ߟ�m��^�\0e|8^�q��3gu�^���!3��Hp.$J]�L��?g��ۏ��l�-M�X=tٖ{��:;@�K��E�>��y�A�/R6(����t�0f��`^�zM�o�Q�E)'�琺�E����~Z%��~��A�v4n��)�1�'�_z>U�T7��5��{�X���ת��j��%�	�T]��9�����!���?�{��1�w����n�پ_��/R�+�qo��l3�D
����V�}?�t��o�e��~$�4ɔ$_�a��	,��Oד�C��l�;_�W��Yz�1q��z��{T,P{��ߡ�U��u�~��R��}NNNNNNNNNNNNNNNNNNǁ����7���ଖ�C��ؓŋ7��COx��YCmS<���Yq��W��f
l�J�Mx�D��$E������V��X�y�3� ����G�mo��q��k���"M�qV=ΊG3�L�zA�5�����U5����~�^"�t�S�_$�43K5�z&��eΦJk�:��m8[l�w�$l�Kq���iĉ���N�-�"�x�	ńS\/�5��>�l��2��^X�	V�0!�ǟ9��瞡������E<��L�oĒ�㏟kN�Io�4͐p�a��=�~�l�9��z�$@����Q,�#$�h�S� ��G��i��/��ޙ矫�G���멧T��b��wީ����FܹCō炼���qZzC�+�b�Σa� �=����v����-٧y<�v�Th�	�ce]ұ�Y��4�.��۞�n�꒗e��R�����#2��-�׃BC�<�秮��Y*e 7?|��M����Ȳ]�Y{��g`X��X�i�ǃ^�g� �ĊUb<�w��"�����K,j�jux����t�k���2�;����U��|���]������i��ێ�;V�p=N���B���_�b��4/@�=¿X��5��W4��{���/H��qד�;��O��|9��f�=���P�_�u؏�������������������th�^�E����L:��_�+֐<br�$�4)c�|�R�W�r�(n��k���o�[�_+&��&��X�rI�Yf�4���^i�Q��H�H���I��z�t�P-��O�1�Wdg[�sY:��y��8�*��]{:��=6����u��3Ha�3�<��Yz������8�E#e^�3|Tϔ���>"/#"���D=�����|�9*��٫�ړ7�8sdJ�b/H�+W��׏eΎ[.��p��l�t3�3F�{����s��,.�T*�K�V�KL�r��E1�v���j��E3�����\�*���
�ɛށZ��dp?<�u����u�}���n:Yŉ�	lOY��p�]٫U�5p�m[���������\��'�v��j&Q37��|�1Di�gɛ�����{R���)��8J*5�����	������=^�� I$��y�-�ux�/̉/ڌwR=k�T����?��U�����Zt�����m[�LF�tJ�3﹢V��A��������̚]��zP�h�h���:VZ����B����b5#���Ϳ�ۗ��o���g�f�-U��?�ǋ��������r��tOܝ͋�EN	�` I�3%J��`EےmEK�U�e���:=���g��HI�,��DQ�$&1�$��9oޝ�	��뜯�]=��M��Ώ�vf��������;u>��9����}G�*;�m����q\�wuB���������~�l<���P�\?Y|vj��)H�>�賰������������������B_EON�g��h*s"��L�5��k�lJ�Y��m����uh�C/���;�q������I`��ϞA�
ԟh�y���!2�$�mx`\��Ԓ��G�W�H?GF�|6�}¤&�/QS�9ђ����dXI����� 2�mַ��\a<����J�Ȑ��$'E�M��iV��J���:JP�-�(�֟G͵T<�Y`�5���%L���`��my��[���2^�Q�ɨ3�"#"�46��Q�C<V��+��0 C6�l'o�s���[�S�7���ה=��Ca�F��%˕}�-�){��+���R��g���x^�=#:�0��5��W���>����ܻO�'����-��B\V3EF���<x'�j�Ѻ���&'&��B>㏀����	�q��|��2��9�렲� Nԝx�a2�=c�T��2���h���%]���'>�c�0`�e\�0�����ǏjU�6�n0�q�/侇�sܞF��;�B����J�:�j�v1��!#d���V�xח-Vz��
��Gi�+󂑽g��B�-،3Y�,`��صC���#�v?��6({`/v�ESXr�i��iڜ��.9����݃�曐������>,�������������������b
 t��q�3`��X�v��0��1〈�w�X���!��������r[��$l���ޥ�#���AGe�n��Jtq1�?]��K�>�6���+-��<�~0���	=^��<]g�u#
o#^�V����1f9$z��#���0�D�M�S�%��3n������`�qT�h���4=F;2=���n&~f`�BiZ���Y4�VK*^��.C[�12����8�<���Ð*B�m��Y�Κ��m��0�2ګh����h������,?!Q�c	��\��|��ݔ�mԷ�8R��f��mO����s,�C�&�h�,/˟E;D�膖�-7��WF�<���vg�����O2.�x��]����������D�k�\����^�u
H�1z�R�$L;?���V�|v�>;x��Ayjȴ)x���pB��� #D�MU�J©����l�UbDYX�l0.5r��C?���הMR�w�`B��bm�P��ی�gb�-a; ,,��J�Eh���F�T�v<66p�c�%
jݏMza����Oa�M8�^�0��X���DIK���	�.L1M��/�p#8���+P6��u���.F�*b����z�y�1.)ȎE�D�� �]�?q]��qMDvRVҚ�m!;,�������������������b
���7\��H���H4F�Ea�qT�`e4�=�QRSR)h�55#�I�eu��N9��a5� ����Qz���� 4�zz�,�^�C�	s�(V^�U��
�0�����"Ȯ��W�h��>i�чWX�7=�<K�~�n�/2����h��F�� �\�̾^F�5aBe�ч�5H7*�Oy_��>����E2�JK�������hm	�fV��|��&�h����/\��2Fى���˟C۬ �7�)*�2��PA�����e��N��E����ӑ�λ@�Y���3_^����/+�u����s%�P^�{~O��!ES�|�F�0 �s!L�.���d,��IS�{z�yц�����z��C�$���x����h��=���9�F�)�Ԅ�xt
90�v�ީ��h@H�"Q��ܱ�vw�ئ�Y��*;������+ghG���ԡ?}��g�ݿ�>�k�ܫ.G�=�#�ғ�����3���D�~�syBm����}6/���n�c�8���
�I�S�5Vb��U�_�0�א:gx̳PMӊ'��,���I7�=c��I�s7&;P"��F�n}ZLNL-B��̧S�:+t���/�+����pmS-�/d�X�xf'��2L0��!̾���p�����h��N�� �	�E|�����/��@�[~^�\9��KW��"�#�MrZ�̽w�es����C	&�q�0�4������c}S z�O&B4�+Ş�u-�0��^�u�K���/ ?�����
O�� ��҅��mo��l2�gfi?��8��:�RJ�Q�
q�+����9�yX����hں�Me��b+�"���J���}u������k2�􂴱2���Qu�(�F2���̫bѯ�&�6�z!+�b��l��{�u"}��Њ'�Os5u`�%
/W�s����-o�W�T�֗�����u�{2Fޱ=`~v4�){�5�+�f��3�,���s_�Y��L+a�Q�.�0�m8.J����t{�W?fZ���s��>�)eW-�/O���;�*�}��؈�r����z1��n����w��e���h�eQ�)֏�SiGZs�x`5�ڍ=�����/�����棜�_������$"��,�C�7`�T��s��{�#j�����۫0EK�P���,�h�G�x~b5����ج��%��^�Jٟ=�K䓞�"���> M�O|��ʞw�|{��=��}n=�.8O{�|�~K�)|�d���uk��&f����z�~E�3��z�L�� ꩣ��3/U�x'�[g�������mcP��l-=8r�kX�D��Ү��(J{�gD�y��0i���J^dr�ch|_!ͪ=��s��V)���3u���KM���>Ѷ���6�'�e�U[M&Jkΰ������y�,��S?�F�� �Ek�Tb��\LZ-����J�{��W'��*�IÈۿ���a:��~�;���Q���9�
~�8�j6*;2é�;�0�`���6�b�Ӓ��˹3�(;��C��m�������^������ܹ�ݍyC� �)[��Pv��3�ҋp<!;�Jfr��y�^'�<։�NE��a��
ȇ���]vn��Ѯ��`�{?�OW�Ĉ`���QQa\+���������������������ŤGx��0��0�{��@5��\�@㊯�g4�|,K�.S��߫���v�3*�+A]s�$C�g~�n%=c�P&��1Wَh�>w��YF�|q�KʾD;0��傇�:��llM׼��'�qe%���0̕_C�G���/�?��W�*��5ԢX�N1��0����\��[�| �Q��Q��2�6H�;�.��EFWN�z��%���F
���)�=}���0Ơ�O��P짶]��e^��m�#zj*"S?��ϼ򜲿x L�9��&_�IF����9�Yd����I��C�]y�ʞ��|2�~p��}�8���ꠑt��({��W+{�³��x&�Y��:e��&��蹍-��4DP����\ėa��ϧ��217m�v`d.�_l�������!Q�L@�rd47�S�)�p���� �'
Z�����K����K�+jz&��ܺ�=w�Y��jG?�����)۟C;jmmUv�-g*{��k�:����� �Q�^����ct��5���H�s����`Μ�r]y�{�Y�)��]y��H��[��T��?�[��<�K��u��2��R�9��8O6���g+{��=p@�j	0�435�[m�N&*S(t\���c�������0��ɨ��R����}����{�>p�0���5��2��=n��,�&;���ø<��<��?1��*>iڕ���������Uv���8�y85�j��5�a~w��Ӕ�?���z��4�d���eQ�_���)�z=�;9�z�D�>$�q�^�����:�Ifߦ-����0/�b���|_����wh1?2������2~��?�و�;¨ρ�i-�������������������b
��B���
��?��h��S 	nzE8Ӊ���\�=�0����*e�j���*;���#���l��>���Wn����42�~��[��Ǖ��=V��J��\= AT^CH�1������)�~&XP{@~/��'�a'��s�+;sS;�|ӗ�xM��0#3,U�z�0�o� �v��x� �y�Ԗ���9���PGo�'�����M�70�E�t���7��[o�Y��h���0{��h��ޥ��=��}``��er��,W$/���!Q�L�L�˝��s�#���Vv�Q0|�����=���h#�fqj���=x��MM``�Y�tV��v���d������ ���^xT���ߋ�Ҍ�$05�<�'I�Y��#>����>�8�������{�����<t�w���x��Kf#�p=E������OG����&Q�����&�x)��h��~�Fe������~�C��3�E��O��O�8t-�cZ`=���|}(_:]��w�P")qQ��m?���Z�h|�QS3����U٫/�B�&2:��h=2Ɵx��Rxn/��������W�Me��Ac2Z��7,a���/�'���o�P�Sn�{e�م'���a0O�nȃ���'~�5S�d$�b����S�/�G�YO��n11b&�da:YLL�W��ҏ�p^v�E�v���޻-u�a�p�|eW���I3�1��#�/��Qq�; y!W������o��|6��/��m��ڱ�9`nbl��1/=�u����;�IXֳ�����
�i�>�9�l�XF���l`�G�����������������������B���g��E�
Ya�p���z�����ܦ�ZDэQ�,JfST�)
�/$[N0#>�>W�����@ź�승`��+�3g ����=����}6��,ES4��m<���64����1����+��W����%&���E����0o�~�	e�%*�0����^3s��x���"��QN��d��9���d�ԼK���,�wߚ�H!��L�:Ӧ��wpV��a4�w�z��y�=`��4�ֿ�V�aIk���j�C>��f2P��O�Q&�K�I��\�}c��KG�a�gԡ����%ы���Z
�%��ۋz;t�P�m�8^�#��D4e{b�Y��8��D�%Y����D��������2*k��H?� B;I�>ct����ͨ�{��x�lxz2���f��&i�LA}�����Q]+�W�z�Q����e�<�be�u�;�Z�d��]���Ͽ
�5��i��6)�E��>���?��@K��U`�y�p�Ͽ����+����K����a5ݗ��O��'�������}yF�vZ^�r�`0���u��)���K�z��˰]٧��7V0�� a��IS��p��rᚄrǌ��/�����Q|w��|�:�I��7�z�0���~�N,s��0V��6�qE����\�)d0O�u�j�-^���Eg����&����1���nT�P�\�}��k��s.w~�z�l�lOa��2��3�3��Z��:��ٗ0?�w���2�~��iĞ0�z=Ōfl�B;���D�υe�YXXXXXXXXXXXXXXXXXL�����8�{�C	t��r%��P7A�.C�ś��Q�j�9yY�u|6b,��� �0�F��3��I'+��[2Y��	0Sn^�jj��{}���>���F1���p��0y&�1��VrS�Ơ�s�y�=�+�L�P@d�d�17.Qf�L@/�U����D�Lf_vp�w~���'ɜjj�q`D��t#ya�Ʊ.�)�o۩l>��;� i�&h�]A���g"��{�y����\��s�Y��z09�C����* ^�d15%����,�]0D[M�g�b�-�A�b<`	�"��B-?����-S���>��Ne�Y2YڽDϕf�� �#?�ܵ�˒9�5ɴ&c�Q ��7���}`^{�
��c7(�Q���Ff�Dkb�vv���� ��G�1�o�Z�ZG_-=i�|n�v�s$�z�̫X��}4.ڧ����ʨŬ�i�D�A�o�ݾ�Kڜ#���f�C������ݹ����7�@��2��m�(�f'�xr����{��9���3�^O��Pٗ�!=ǔ��o*�Y~a,ɓQ)J�Aӯ��n�粿���y��;$�01�qF ��P������n���dcLV&�S�φ�L��ƞ���[�����G�0���dkWc�䲘��&�֎�=,����$�����}�qɯ{��*���|	�W\|��m2��N�$��9_�r����d�n,a���/PE��8�Wϝ��m�15�����ܬ쳯<��S�O�dQ��:?:wD%��,�,MkZ�賰�����������������(-�1�gx��k.`&"ث� ���wܢ��K/P6.+�M�X��Ĳ�����0�\8�����Jd&X���YY�5�\�ia�I���uԀ9u�ŗ+;���_>������N4�����)���� )��<aQ{�G�^p\�Zw�PaxL����I��q��LJ�$}��eq�E#N3�jk�@�d��K$�.k�r?HFZ>�:���Ct�B��*��lxm��_^�lSj����K.U��5�){�Dc>�AT��w"��cO=�����p�F0�
�_�<Ht#ʏ�*Q�ѣ�f����u������~�>���x��zQ�W�FÊ��Ay�Sk�7���;�t-uy��k��D�Q~y_�#Z��C�<�c�~�礃���/~Y��Z�u�V��Q��+�T����՗�9\~<U{��|}��ִ��z�\0DI5c��hc���xq�!j@�$���� J�o���}�g�I0��A�nuZv;�������l��ޗ�P�YB%��LR�KQ�a���PL���P��$���h��Q�r׮��&�x��y<�F�.��(�S���X�!<�W�95����u>�\_4�����"!�83�ɂJZ&a����qG%�	�0FeiD��1����'~�B���f$����v-�EY�=���1�����Dv��ъ�̈5*'�s9f�a��?��t��|^ql�c�t�1��vG�-@���3��f����֧0/v��W��}�̸��������Λ�߫,O�����S��v?��HvN4g��Fٶvh�?���8l�W������l��u�Q��Ȱ`}S ���
�{aK����+vc���A�ka�@{dNyE���g�L>at�`��Ĉ����3�x/�/������H�R*��}_SXkVtc\�u��M'+�mS���W�r0
)~5�-��/�ͩ:2x~��_(���n^�̮ a+d�7��+�R��b��噀�f�I��LO����W��(���ˊ���q�F����~��a��/��R���7����v�Dݍ��2�(��z9���u�ܧ-�v*�����_?��ٳ�=��s�]EFkmW?����O�1�(�o� �h��T�������w.��38���6���U��Ҁz������/(��@&�`(n��O�|[�H�o��N�U�C1Gʜxx���")��I�ϣ>��h6;>������_���u���|�ܳ�'��{������meo��&e{#h7_���W=5��'��R���^ILGGfV�3*p��o��о8�f������gD�ʲ=2WgM�v��~����\��w)���Ǒ��vTڑ2�X?���	���}���.��~�5����Z�O��<܏3-Sv�Lh������|�	���2��bO��C����Y�=!��2��Ub��c��r��J7@vj�t���&` Z��p���-���!Qʏ�}|(A&ĉoW�ݻ	�2=�[_���7jdJ��F$���m�u`Gԍk�Wvz�����R�:Ԣ�|�m�L�}��7����̳�;�D�?�s�x]�b�ߖ�Yrcg�Y������<̷.�	fc�uX?x�ɇ�=ڋyZ,-��k���U6��Ҏ�
��>�) ��gJ�<}F����%Z�+n�8�������paY�b�T��v���B����m�~z�/�7!����Gy�?<p���g��Em�BhH�6���`fէA�j"�%�'���
3N��F}�����0Mٛ��>e������=����J�l*w���oK(�\b�U�p��0�
��YR���]a�:�hh�E�ȫ�#3L�W��(0��'+�5���#s���	�4���-&�?���gA����[0��&R��,���l�K`�	.�|��P�i>/᪍M���=K�Q���V"��]2�����3��a������^�\��b��j?��8q�5��ud&��P��[w);؋z�z�q�|_���Z(���1�&�����͝�#r�0��*�Fa�v�Ah`�����g.c��q�G��(� ��(���E)�4��S�R�Hj`W�~&�}��O*{���7�]J�����C������N�/~�s�^z>�{���=��E�-a�#S���h0�t�c(��C�x=��sʮ:�|e?���SV��/���`�-Yz�����Q^����٨���[��i��ǉ{a<?Z{��-��{0o4��H�a�H�#p���D[���_��<��Z���Np���8��{!�W�u'��y[�o�6Ĭ��bcb�5���N����p�{뭘�̶������7��d�Ɲi�N���Uʞ��,e[R��9C�N�<Mk�3�w�nی��u��f�������fs�g1o�r�W*�y��={|��3g���3gb]�����Ʉ�8�%;H%��_v�
��;��>/iӱ�j�{�h��?
mt�9U�Dw��!�B��gaaaaaaaaaaaaaaaaa1P�B�0��s�$�naHT\	%q�s�}e��X�cY	�+�Z�ίy%|�3V��ң������;�]�+Z���2ʪh�5�3ʣ�z��+��¤�}e��>��X��M'���Rh��Z�J�K�I2��"�k�	�P��Q�q�4۪)��_T6[ �,R#Z�?4���.1���8lm#�ğ�(���� ^u�hEF}-%S�V��d\������`�ɔ��@\
�u�������y�Q0슃����S��	Qx>����8�p�1\7�z�c;���u�KM����ʾ�:��&p�L��"qa��QՌ%�1c2m�y�(�h��>h�R��7?�Ae�π�@\<��rU���=�Ke����>�l,��R��
�-�G~���+��>�����i��>�F����%e����Z���|��]�+[׊~ ��u��@t�k�A4�K��������p��R#P�ҰE;��kJ��&ϡ���і�(�.�a�#S�>F)O��x<���C�/U��{{��;ލzl�١쬹�@m޾���� �
04��~��M-,z�j����w�}�݂�{��W�8Fa������#�|��5ʊ��O����w��G��^�@�\d�ș�/�O�}aF.1�����@�žchgQ�G:�vK��d�ty�0�%}̈́�2���q!
�&�sP�w��k^���qaݏ~��*����(s'#%<�����3�q�����x���@k���1�a�X��|⊩�i81��ިHu�[XLBh�p�bBc��?�*��X1�d8V�'L���3��j)v����S��?�Z�^Av��g2=�^QvfEq\c$d��۸�5e7l��<�}	2�	���a�׋8�|�Z�����{|�G��W�<�f@�<K��#1r0cԌ�4$R�	���{Q=�WW�Gه�\�7�`���	Hy���nXO���@���gaaaaaaaaaaaaaaaaa1X���	��qe�H-���`���o~F�YI0����<���g��34��QX�+�ϬG�ϟ?t����>cq��N�� J�	�PK���3��v��qO� I&�����=H��!���a�����X�(W��?�|&EV���(�[��%�#�zm�������AN#wlVv��]��g�̊%Yɸ��(jODy�RNӣ��ē�|�
�+�٧Z#t����J���+�¬��	�p(�MS+�+�L�,I��5�d�tC��ч~�7GY��{������#Zr������~6�@��ެ앗���uh��c�#�<ڛhꕖ�C�K�F?�Ь˦P�_�v۱}Ѐ�a{��D+p �X8o���M`,e
�d ���Q��g�.X��מ{Qَy`�IT�D��s:�,&��LF�Yf4��c`����+;����^x^ٶi���3�Ѥn��`WX���ke�����]7�s��$�z��_H2�/�v�ٍ���ijH�e�Y��]f-��0�?{4+,Z��0�lF�IF�C���f,�0ނL:�t`��EW�Fyr��s�<�rԢ��$]�L���{��T����2���q��Þ�0�M����Ja�I��6<��[P��bz�)՞M��k �̖9`���۱�M^��'�u^SH�15Go�i��5OrB�@ScP���F�kф���r�>�|ǻq�ߢS*�~��))�)�[�	���@�������߹ݶR�B�|��L���8�#��aa1�P�s>��$�?N6�9�U�j�`��<6`6K	w�"��0�\���u�':\��q�f����%>�ǋL6r� 4���x��-`��9?nlnT��;�d��S/?${� ١&�-nԿsMnW���g8��:��3��=����4����K���ձ	p_ړ��]��e�ڇ��0�+�8���b]F���qT�,-�������������������b
 |��ZbW�J�}�c�V��D��$?��1����� ������ VD��.ew�ڮl��G����I��${��E6���3=f���v��(�>�����U$e!�Ez���Ǟ�X�޾����&�c��?�G�_=���]ʮ\f^��$݈��'T�8�M��f���ރX1��X�&�K0��,Qr�R�W�%Z����M�O]/�s��b
�p�~�B(��f:LKX�M�>�6`_A���X߇��Iwd�>߅�Q���?���_����l�O�Ϟ�6�}O<�l!Fm2Fy&d����I���?�}畠l����so�v�c4`�X�0�|�~������{v�|tŤ�>��&��W^��Y+�R������c�ܔ����(��k�a��G�L���60)�	(ŉF���b�r����㯽�Je�s��FDg-��|�ޱCٿ����+0��w~�]e�y�|+f��x��)e;�`dI?d�G��2㱐�dD
c��'��o��6e?p�o(;���ʮ}��_$�}8��˕��"�x7�+��
�ϬO���AX*�t�=�E2����#�|XٖH�	d�%��-RVh�ѯ=�;�����쐇��t;�%2BO{�p����s��q�E���"��E��fD	��Ab�7D�e-5Z���]�B��ĸ,�$6��(�*��(_˷����Ǟ~B�׃��:$�=��<z4�yܗ�~����O%��>_1Lk2���茖9e1!`6���L��ϵɔ�t|�N�Qb������U�`�{e ڽ��>�����}x�����7��54M�-��pG��e�e�*�t.vE�c� �<Ѭ3��d>O��@�(�}~�8�3[7�����g���$��2Љyqc)47a^��yK��l��I�;0��i�c�C�V���d��ߏX�P�c�te/��ۚx-ˏ����:�~���.L�~?���/�F�G^��8[��iQ�G�7d`D#�1�������2�,,,,,,,,,,,,,,,,,,� J}z�Q!���h,�j��{I�Bes����I.)�4��YP9�'^��_ݏ��~+@)j�y�X��at�s�+{֥+�=m����FX��|���E泖��FFם?�^����9V�f�=_��7Q����6����*�b)�y�)2��2mj�	��e���v��`T��կ� �P�-%s/���J�w5�#����
]k��gԜ0���^��>J��0=���͚��:j��u���7I��xē�܄�c�Ez0��VX��8/[���k���[�x�sҔ�v@2��<�j�εF�yL&�ɜ1�d�?�Tbvcd�2ʫ0c?���+{���w�����?�(�i�3��R�祥�M�t->GYo�Ԣ;De�Z������2����$�("ȷD[������K���O�K����<�+�G�Y|΅�ԫ�1=��kF��|�J���(�����L�x�6lD��݀����g!_��_�t��"?�vfm�?�����TGm��՞������'���ZFY�G����`��������#*t�޴���S)�ׇv�l$70Db�L�F�7��Ύ#��	F��B3���nP�������k�.hv^p���^���x6�Y�����6�(��O��/}��ʶ%�y�m7�W�id��{}=�ch�G�����矉v��1aF뒔�^X�0D��ّ�#�bT��]�~
t��~MG�Z�-���ńc�V�g���㎉V�!0�����3��֘3Q�����>�0^��z����=oc]�S��ֳG�����7��5�������`^WҌ�3���ΐq0�|u��?{;�D�z>5�c2o��Y�1;��ym����a����K�<Jr�������cǏ){� {���;ޅy���ۃy�k�v�ݼ	���;_�3�N��`�(żV֏D�/*�"�J��3�V��*ex��Ũh
�ƪYTh���gaaaaaaaaaaaaaaaaa1��B=��K�E��KC}X��Zh������G��&�v�������B�n�&hQ�R`�4�Bc-��R�`'Vp[����Bkh�,DA��5̵h'QР.�=LN�#+�)FMrIV4�Ρ]�l?��/����V�����s��^��k�i�,����YO�+�3i�Z0{�B_ʕ�'���{��
D�4$'���E%����Ε���&|��_��}���A�u2��/A������9��u[��CPK�:���fX�g�lDq������rxR����x-�'�%��7�P+�8O�����䨭�	&���9�a͵(��
s�njp�670��&ӯ���~zX��*5;#�����-��(5����?��<{���A�%C��w1Fa*��o���Ou��!���p�Z���v� [��-�t�Gd0HQk+����ѵX?�?���/�E8c�nMM���Iڲ}�����>%�s��f��K�s*�.ߞ���w��ϑ@�k�Ƨb���>�fE�Q���ܩ�n����/Z�l� <r_��W���(���f��ɂ٧}Z��"ů<�	�~�K �A���������^3����teq����pJ�_E}}Ҭ�=������0MF��Gy�s7A��}��({�Jh]�Y	��o�}��[-����	�=H���#��0/hh��2��H>Mr��c2�\Ú��M�5|���bb@k�jM��;�Z��@f�T����*5+��@	hȞdLT�B^�/,���2�N�6����}��GMx���T��N��d��1�N1c�1vr�Oc���b�=�	;�r�f��33L��3�w>�se7q|��u�-��c_v4���`����X��yC��D9q��Q.U���zT��ބ��X���qk7`ܽe���(���	�c�1�_Z�q��];��z��f5Mg}�qϯY��j�P�2�Z�f��3��q�K8K����F�拑��2�,,,,,,,,,,,,,,,,,,� ����%FFa�H�+��:�*;���K�S"��&�p%���ߧ��MШ�跭�`^���f���h����o��qow�+��l9aJ�w���c�sZ>�o���>�GY�=w)^3:������?��O����&e?t�����
M$aXH4^a�E&F}L��ao�O"���^\�3��3K LKњ�GAc�|a�;~&�y�f@���B{^B'��F�8a���!���
qޣ���`Ւx��`�u���y��_������D�����	�%c�?��M��`y�d2jt4*��͵|�`���<���m S�S��fWk
�>o���ieq���f�&�2[��ɧ�Tv�^xD��T����ayR�d�J�x2�8�����w2�zz�$L� �9+�Vv�L�SMIh���B�a�X!������y0�6o#+�Ĩ��M�v+�%-T���=at����[ew��#N�rAkd8����E��yU��Y�����g�}���^Z�y�*}B�c2�B4�B7��co�[��y��/){F�~m��ⷾ�me�(1X�&�D��:
��T�Ն��p����h_�=(Lij�<�_��(`y<?C�)2V�CxAƙp_�V]�O�̟�O;~-���Μ�~�(mo��Ѐ���a��[�K�w���s�]��'o������^����n^�*��tE�s�L�`������1�&�uz�D@3��E)�LF����?	D�'*#��ߘ����ߙ$�uS����8�{�M:�M��&ӸjȰ�Z�-i�.[&���++;4]���e VO�;�~;�^ـu�&·�4����bv �>1d�����R�H@�u�s��nZ+��<�y�/c�����A�ى����P�kޡl���G]2e�C��q�wZ%���h�5������8)���3�;-�������������������b
��B������L�k.���k0�tt�H�g��AbDd3�L�߄�~���ntԁ���,F���ˀ����|Tٖ�f�L����Q)b�'<L�'����]��k8�t=w4#��>�{�~�v0�^ۊ(/�z�ו��羠�h�e�D�O<�L���
�����x��g�=>x�%B
`2���!�!�t��j���q���q:��`B�u*/B�m$a1�%Ff�·�0�[�ma\~���)�Λޣl���a�I0Mz����jh30
�=?A4��и�i�ģk%J�P�M�)`l��%>�S���A32��s����\v��,>>�ɑ˗�.����~f��(ڢu�Ƅ�$%��]�|��)^������`����Ce�w�@z�u�Rv(*�]�<�u�����H�K�P6]�����a�A�{:�/��j>�5qF���Ӗ*������0���ݲQ�B�`{�=�|1��~��#]�L�����P�L��H���(;ԋ��rѿ���]W�&�h�����W���в(&�`��~]2�q����_0(�7F0�}^�X�}d�t��-�e�-V��M`V�q�پ�_{�5e��D�,ƈ�U��,LLX�кx��t�#��{�S�'�=��ի�?�tD�?��y��`��:�=���oͿ��5�S��g$:!����01FD�0f��AW��"2�P9�r�yd��F(��(�oaº�|ׯa�N2�M����7'�{�3��+Z�S�Ac1��S�܀��,p���;U����NF�1�&J��f���l��e�^����
�d�!L�u;����Rv�9j��.&S��ׂ	';��1|K0�}c=����Y�6\�y^���>��4��چu�][�T��j��<1�Q�����:��ۀ�����.���q�'�l}S U3����}3[:�m%F�x���{���S/��&���$���t��ӕ�������_Q������J�{R��Y2Վ�0��0N�F�ф�~�hp��w���V7n�
�ڛH��R�S����H�²���ċO0����j~���xC~%� ɇh�� D+*��6LO��o��y$��ї5(D�����UH�����h��`.����?EfVz�=����y�qekȴ��XF^4yE�R{��Q��b��,I� ��xn��~�d}̞i-h�-�`�֤�yw�(b�d.%�8>لrl?��k�~ݔP��?��U�C�Z��k-��$�S2�u���x�����P�7�|]�`0��L�i�)��F��u�̬Ԝ�� ����D��d,i�<(Qޘ���.�4�w�ڽ�8�(Z���0C�~KQ۴P@�I�!�n@9�z�g�	iW���A�
�_��,���c`x���7e�7�_/��vh/��\x���V���9��6}<bR�7w���̳x��D���J�Ak2���yf�.v�h�o�vD^���M�Q����9�e�"�_k�#X��вg�V}�Dc��(58��W�����v_��Sv�E�v0��oܛa����K���%���w�b?����qD//������X���&t�!7��}#��'�Ȕ���?�=H��)Z?a̾j�(��p&�oj�'�f�3阗üO����s��y��~#������h�-���.[�&Ij����+
E^��ly�3�Lh75��{��b��D-�4����딭�r�섷�a�Ǉ	�����s���h߾}��|��"�-���ɝ�g���-���c���';Z��/��>�r)���؁Z�0���y�XW�e�YXXXXXXXXXXXXXXXXXLT���註Xٝ� �(N��w�`�i�+�*�1��Vh�>�G��8V�[`�h�?���%��4��7⿎�Z3�k��T�	�3קc\�]4w����6e��.e׮{E�s������4"����.��/����^~�G�̩R�C<���A�1~f4^S���ѯ�'.���#ZoJ7���6Od��`jm��'�9W4�x^A�?>7�c���.0�by���t0+�I&�����{v@k��a0���ۥ��;�uP� �*�3)Z�(�Z�J(�7�,��[�3Wr9h=�=<��x5�Z����Q[̘�l�a0�<2JRn�&V7��Z���"Sl�Q�G��s�A'�7*�p��[�<�7Z&�����"�S�lh+ ��60�(w����ɑ99�(����OF����M�z�s�)�� Wˠ0�p��(�0U���֒!Z)7�y����>k���MQ���!$��?�L?��.K��x��Բ_��(0��;�9s����W*�Br�<�\�ںK��>�v��!�pJ��#��H�p�(��ߏ�U-��g.9S�U����>��&]}h�u�.?ސ���h��<x̽�(�5���f�Kqj���0L��BS���o�%�1���\�U�~��}?�/�V��+��{*��+��`�5�af�,*i��߫MP�W��b����i�Ue�����'���1�������D���̝��w�A�U��[�pW�|�t��s����/����&�;�j����i��1�8Ou�����0m%�/�D���q�+;9���'���˛56;�]��o�E1^���mHb���{�z����<��>��T�f�WV֗�����k����5���'��n���]�NeE;��zs|���^}㖶F�=2���H��:96�O�賰������������������Z���
p�L�����s�#D�feO��%Te�}��u`b��:0R��k���=�v������i�7��1��
#]X���?�$��ZM��t)���+{�84�Z�K�1�y~ώ�������pii�y�s`\����C�Jf��	��T�0f�0�J��ݸ���3��݁J7F������~f�D=.�CRd���$��͍m�~������	0d
d���M�Ys񼜾	�Y�����z���̞����ɨ?_��%�M~�����
</CYxbf.^�l���g�����S���H-5��	3�
�e�l���HS����?�<�_���̟�L������
0l��!�F�9���'YK�ψ�}&Qu:���L�+��B����ܺ Zp��a�h�R��"'�w���{��_�ϩ��%�cL��V������@��=Џ���8�!篂g�o���dn4�D+$Amֆ�Ʒ&�������C�0n?�lw�s�ţfd{��c�ch�9,��/U�%���c3��s�y#4W�<�l��a��q����h���K6J���~�����9c�t��8��=��C�8���hd/���GA���W�������/��V���:��^���~�쨴{?�Y3�F�.�ah2��)0VZi���d3<B���~}a0����~m��n�u���p\,l��OG�����y]���*�o�Z��������8��݄�-��f��"�^�/NR*���&��c�Ƅ�������&���z\0��`��9�� �&���������1�UHk���?l�����b������5�0}�W��RٳOGT�Rk���tB>�>�#BLk���x�eo|ǻ�����Pv��ה�t5v�lٲ�w���`J�|(�.��7��B�;e�8;}���� R��[f��2�,,,,,,,,,,,,,,,,,,� */��ɐ�`��9	CGd�'Z:����[��ڮ졃���
�����v�R��u�r������� 
x^&�t���>�\z���5�>�,�����+{�M�UvzZ*���:���4�fO�����]ra�5����D�5�z[kZ���o������Bv���*�|f�o��5�&3 ��������/}Y��Cc�G���2z��:a���3����<�:^��կq��(���5f0ߴvIT�XeZf��#��t#��H@Ө�󜢶������_Etk7��%�4�� }12?|��]��\�Gf�Di��&*�74��W	���E���H�MP�I<-ô(L�o�ZP�Ϝ�l���X��J4)RIԇ���L!�ի5��y1������`ǩ�V���h�E5q�xn-?�j.�;ͨ)Ȉb[����R�Q�#6�	2�?��/(;�Qt��V��e2��/���&�;0 ��|��f�ؾ�)����5knP����"I��א9:0�|ęOyp|?z�̕�������6��Z�r�DC޻7��.e�Z��x珑��v�s����)������(Z�W^�~�߾����?���^~â?{��kj���"�Gݘ�� �it��0��0���{�f�[!��D�p�}a����R��1?v��d�v�G<�Y7Np&�k�c�}��Imբ&[{=i�;��G���N���Ǫ��4�/p�*;O�ì�㽘�z�	�^�/�D'�qSw󒧞��D=Ǎ�(�Gӛ1n\��le]y���<�=0]��/c~�H��5�\���=��ޡ�m��[�p��������9�I�|��A��+�܁0��t�`��3�w�X�d,�������������������b
��B�vx��sO�֊#C!p"�8��i߱{;�g!"Ÿ��k}��b�sՅ2�����D,⯷˯�6��Ce;/��V2���,4�Q���w�M�^S�L�����O3|�uL��\'��B��j愡�&!o�h�}��W6����O?�l�̞d���}������}E�����R��W^��k��	p�����Cdz�#����̅h�L���5����u�8>�i��(Rl�P]���0{�n�����Ԝ��1�	A�L>� 1�<�v�O-�/|���O2�ă%��(�j�j����ؐD��h��4����̎#�=���_��l>>��Hw�������T6O��G>��"����8����Tv뎭�n|u#�_��W@��|��ϩ�W�75h��_w���,~�[M�Y�a��@	۸�'�lt�dZ2�o#��.>m���d�Nkӻ�X�?�c�D����=�|?�^�|�i��w?��q�ا������/G�~=�-���Dk�,v�`���O��]G���ۆh����y�	e���>~Q��]���ׂ�7-f�Kݺ�ѷC]�Uz�5�H3�˿7�B�Y#$�we��ʉO��t���;��l�
�������Q������9����s��E�	�LZ���+EK7���?�Q�Z��)�x3�&�m����ס�)��S��y�(8�$e*���f����v��L����(=^�q�7gc-d��'��s��>E���'�}J�l�wz�<��e˔�KR݌*Z�íߑ�ȝ
��Gz1� ��:D�}�Q���*�Sf��xw�^�Se��xL%����q�56yc�����y�����{�#��u��f c}S UG�MD��5�cO���8�ƙf�p!��̢Cǰr�r���`{��
�P��������m>��$e�hI���?_�{z�����(�� Z�gԯY�x�<0��k����/{�H1\��S�>�?�VX�v��Y��!?:��0)��D#�퍄�zjh�kB����E�j�y/U��(��1%k R>fS��5�\#j_��hV��?.W���/"W�!?3p�n�w�20#����f0�b�$�G�sy���sg�2DY�$Dd�у8>�NF�ɧ=��ׂ��S��;w~[�FjRx�f��ޓ)x^�q�+&Q_sH�.Q�=�h�y2��J�c�x1�*��/�X�_�f��?��'>�Qe�2�Sw�~�̪�qz��E���s:p?���Jeo��w��׉�B��0�0����L�k~�?���s��HF��o�ݩ�}ѭ"�?Ř�����"���OV���'�
A�95$=F�ϱ�.�y(�9X�q������vɺ���G?��3�+{&}��2lhj;FmZӓ�ɞ���?�����#�����y�ʋ����+������@/���50����^�q�����2���L�5y0(%�y���f�^>��$l/�	���3�{�+�FaL�0��j1Y}������]j�zd���=U���U�]|��&�;���&��t�H5���g�m2vTLx��e�O%���©��1Y�\������\��Wu��}NE1�X�~	�!/W,����ˎ�l��ʦk1�MS󯽮U���/��bx����0��HQ~˞�T�;g��+�^���?A=�ܹS�\���*v�\p�55��֢��G~�h�be���~�[F�賰������������������:�nk�Q�������0(<=��+�}`25Q�*���}`�$�b|х��M���%LrO�!�T뀑�|)9�}d|��e���{�rn��5��4�Q��d���c2�4���]�)z!h��&�hv��\fJ`Ϲ?�`pM
/�C �W�J2(�<\�����Lf�ԍ;���|�9�x��صո�0a{� Z����ܧ=����fV����TM�pɛ�;&C����
�I������4o.<y���]��YG��D�(��]2�w��C,���`�F�H3{t��0&_*.��&a�Qj��T����`�W	K�����Q�X�V�a���)_:�|H�q=�,�h����e�A�n�0+o���(�c���D�o���.���uk��x�/�H50���`*����\�R�x=�{��TCM|dzC����6W[�]I?9V�PF�vH�%8�����������p�60�
t�e<0x�2��pa%~����!�ț��v������"`N^z���GS���P�߹u��}ݸ��s���fI�Y9�r�楠��c�m`J�Po�-�L����L?�?m����`^{&#�$�*1�<C�0�*����S�1c��8���`�0���aB�?���s���3�*}_���ir��A�����{[�2�F�*ǟ���Q}T��W��k�W=:U�C3���~����ӡ�';�<��� �dʹ���<�� �?���V�Ίy�0�j�V��m=9�p��EvZ^tbD���(�/���ѷg�ne/�|9US�KW晥 }���քu5��U�d�Ao�<q�+�̲�>�)�*4��TXKm�$v�	���W�eA��DFG-2�,<���`f��A#��+Ź�hXV+yP'�g#PMƂ~���~�^�~�n���^�f�~&�����t���Rߤ�ރ�x��:���W��|�.z��+V�t
&r�B�=������G�+���D3ʡ����������%+�=����<Ʉy�������7e#`����;��ǩ)��t�V�0,�r
aD�R2�h(F�Dt�g_�����Vv���|���D�E>�����ݲg���f0�����^�*?�$��gR��	0NM/��-(��#��K���ge��Z�m�����sYA��b;���d\��K��k2.��`~z	z��~�`�2�G��C0�>�[��삙��K��(�r!ėPx!�m�LH���y���m�@5�z2Y�&�6�#��̬ix/,����e������=�0�*�;�n����~��/����N�y�d%
6B�EEK{H���v��cSzp�?#��>	F�g~���6�"���Пe�x�LSq��)���
?���ʦ�}�hӄի�o尹��U�P�eEډ��<��Z�Nl�{/ͨƵ��{̢�^8��Z�/�Qv��29�O����Q�eh�J�������`�e�+�>�
4�x%y������L�˨�i%�ѥ�L2&Ѱ1ŋ7�ajPV�{�OLM�p��9�ƭ��;��6�0�v ����O��5)���k�q�����+�W=�y�/bd��������ˤ9A�8�� ��0�O)���z0�,����󁃘7�4c|��	cҿ#Q�˨�iܧ6�{�?���5���*���gaaaaaaaaaaaaaaaaa1Pq�OK�H�Psϰ&tL#�^�Rr�K�=���)�T<g6�3�0���RO��	�	+�|nm���ᣈj(a�"�#*�h�};Hm�A���+i����hO7��sT�U�Y'x!��+�<��/��?�5��i4`��0f�h�[q�� C��_ޣ�{��^eO?c���^��?ވ3V��l7��>�$��ve2Ո��7�;_�_�r�����Q~�m��=���v��v�eW*����/2^�F��M���~ �%�Q �$]��e�߇PDL��h�E=�<C����훕���w){�Z	��X#-�0&Y�V�����v����Zf�|f�l�t+u�`��s%��h/��m����G>�e����0��$�؈���|%��Pn9
��Qj��Zc��]������eD#2;�޴�-�"��2j����qc�ш��^�!�a���G�Yn�b?�������3q_|�Q��W��Z"7��Fe�/���UW_�l�<�#�<��F�����B��[>�(Q�%�nC��r{P�!�1g����gh!���u����W�����m��U݅&��|�0��)��n/2�	��aj�檢�3��&������J�O❯��x�a��ڠi��&'*j�UY��j����y~u1�k���w b��������q����A��)��O��t��a�O��+�#;���0�H�1���P���$��M��!�؉3f����:
�C�7ŝbs�,P��&��Dt�fL6������2�-_.�賰������������������z��FG)��
�}_�4QLc\A�w�F{����3���uu4_�Jhĩ$�4� �M�` �1oh��<�dp�>��p>&X\4ń	��v$�|�t��6�'�>��<5�5��x�.�GI[.$]��Q�����F���/��u|�K6[`O��#`���o���wG�X/�&�~p���y>^��gC�>����
��Z�����̦������������:�v���Z�/�T��9O_�(�y4="��=ZҾ�xޯ�Vxp���WMK/CϘxfB�A{�d�H>k�۾g����Y�������=
�ԑ.0��M'�c}-��>񇿭��vD�z�E0�2�臝$�`����_�f=�P�L��%Y�_�w<'�mh.���UK?���t���v��槕��O�iY��_ѥآD�rO�>L�Q�MȚZa�'Ҳ�\y��=��q_<��z��vw��M��;�{T�oy��1a�Qk������d�w�h�f���\f�{nx���Q����^�~��:��@��n~Y���'-���3����E>z>s�I�rH��0����%�u��Ǟ��,?5k�iѮθ�\ec���d}�kj�?�V�xf�������S���>
��Z�9P,�dU�3�o#���#%*��g�?�:�2�"�џ	C>���g�騿�a7ӕ�!�s��Ƹ�&iЉ�䫀�ޮƇ`�q��r�y��m����}�J��Qߍ1��'�}�F��y&_S�g�U6��d��ǘ��c�&���H8&��dBr�;�-9��%N^m�ǥ3;�3��;]�zՎ���{����ͱ�JZ�������t1�MD11�^��x�{nH)��ߺ"�oT�e�YXXXXXXXXXXXXXXXXXLT���6m�	�z
|a,�vuw�{2�3OMa*���:Yjӥ≷&3Q�ʍ���o�G�������c�Zy��
�x~$
���[<�zE�� ��E�s�%k�`�8����r�P�"T+0x&�'�R�C1���|�'H'#�u&3M6����ÅY��D 0�'��%��*�Z�?W{ox�E�&�`�P54&ͨ����ff���j�S�	���������l���T���+����Oٮ"����R�,��
�m���>�؃�&:�'�H@�O���k��~F� *̳4ӡ�?��}���);s)��s��G9�ڹ����|C�=��xl�M�H��t_>p3'�|Ҿ�q<���������(��ko	�������b�3��q5y�Ɨ�zcI�H
̶�Gl9�L�~ϒ��s̷�FF5&1A�['������;�,�<��C�Ǎs��g8hi�=�����-��q^.Oƣ����pSs��-W������E�%���>��5,����v��\GMG�L�T���A��I�PH2�+ѹ+uw�z�+1-B�v�i��~�y�v7Iv8�<o %_Bf]�x l�P���ީ��q�EN%N5��b�x��/�A=1g��>W���7Q��k�U5w�aL���Mk�z�kH��B?&�T.�qi���t]H!E�[Nd}¿�4�k�d6&0��I��8��\�*�5���b��as��m���P�e1w#ǎC�\�O$��l4�yw����2�,,,,,,,,,,,,,,,,,,� */�q�0��J���aF?3�����^��\6��,�F�~�����js/Z��9v+��yв���ƟN(�-�L�g��.�4^���d�i���6�p&�B �J�U�nJ!0��� *m�!5!�	����=#�����xa�uBl�`��=�~F�@5�c�3�X��R�3�}�b��]��E2��-xn�}�����8yW�At�Y3��'�h����&���j}�^�4C���0|���A/R!�HO���%׋�Y@��y`����g����3�E�a��Sձ`6�����hii-Q���"QWC�E�f��S$��_=�l-�oe��{X#����s���~�j����F�O��-Fh�ދh�q����@7�"����^,��p���rn3�O���hլ�>��o��`T�ؾ�����.2���{{Y^0���(o�t���^h
S/W s0�D���v6ԉ�����1���|��M�t�d�ݼ��J�%�9��sB�ޭ̠���k'D3n�a�̾��"��%-]I��/�J������_%�a�}X��[a�GUVS��a����<h�ғd���NǺ�iz�k}��W�I\�q�h��%�I$ek�9�������n�N�O�;#���Q���30/�2VB�H�8۸2j_�
&_���q�ok�H�P;u}�>^��a5��L?�e,�������������������b*�ꅾn��k9�`��Jb4����Z�T���.+ͅ|ޗ��#`���ʩ��?0|@)��Zoިzݨ���~�����#n0�¢���}��<�A<��?!ͷxbO�p��� �=i��0�T��1�S��D�����Vbb�S]AGi��.�
��@:�&�0�I -�5�B5&���A<����,͍G��|��o�m��s��Oğ����>�<5�Ja�}V����F���A	O��y���\̬$5����6u4L�uPd]��.$ڲ��t�ڡ�4`�x�XfiA�ϰ�d+jF��1;�d��|�����ݬ�{Ia�1c�s����h�r~�10�Z5L�$4A�u�{�+�0=�'n %�%� ��
9)7.4��?��}i��c=��t�q��5W4��lܽ}+�3(�y�#aJ�����j@1�h�����3������xl�2h[���8���k8@���3�F�1۫6��Txχ��C�&j�P��P�ڱF�¢�5�J̿a��j�����LML�	�ho�Y���L*�_�pj��H�\&#�4L4^�#�X�o��t��|㕎�X/�F�td��!el佺��d|��}�4iJ5��7U�#(G��hT�92>�y2*F�'c�J�τ̻�Eܯw�
ءR��{���<���3L����O���>�)���z{zFt�hK�iF�;z��+�;v�P�dbM�Aed2��
r#��̕`����d����x~�&\�Ig.̛L�
`���7:?N��ܫ%)��5�Y�&A��K�����k|\���J����k�pIQ#@�Aݝ��e��'�e�~��6�(�u��T*���}<�`v�(њ�]5��7J&g����q��L�.�,�)^M��5Řo7��:A�._#��b2+d�"S A�E�O�oB�g��>j��_�h��"�;8��*�|�5׎��&�H]=�O�P_������@m��x %*l4�����J��z�'���ZF�-�Z������z���?I2�{;�����2��nd���>�35�qy�т[y�[(R8�Z����å��_��x�aE�PT��������YkǢ��f����E�ۃ�I��T�ѥ]�Fi��C
��c�4j����ꫤ���Ӑ�r�g������Y6�Y'8�b̢��E[���tX��GP�>ݱ;�b2��c��Ǩ���q�T!H�b8�=
����Y�W��8�e=���$�B$'w�9>��Ή^��e��C�/��<f�^�Him�8<�y������Z�<OI���*�����n�Z/Ɲ[1^��]�;�t��Ov��u��e�YXXXXXXXXXXXXXXXXXLT����%�P׶�w��'��)QA��#�z9q��]���n��c��Mk;��h�U^��g���Ĩ3���+�%m�JZ��K9�h�&b�L���O�h?SB������y����c2�"��o]�F9�'�`BMkGT�� 2�R+�M�Q)S�J�R_7�	2��w����`�0�ȸ
�6�0�a}v�~�_�n_E"F�~q��LTnsEG4�B)��/�����q��yge�����9����fp�8H���������ZK��[{��������k���ʲ%�:)Q�(� H
H\č0�鹧g�﮻V���D!#+���{���]�Y�������y[%�Z5��c?aF+%t��?�P��{kw�8�4E��z4I{�I����"-W�3�nՙE;�JS��G}�:2��YD��f�-;�aV̈́�k�S��1Q��r�{�Bźx��3 �2]V��Hi��~*��Nz5np�ws�0v�CŌ��}G��4��5o�,��Yx�W��[�Q�E�O�������<��qL���(-.:_�ҠQ�~�78��Ԍ������'-�]�%:�㈽H��r�i�x�x���@DgWo�~����k�ڒ���z��緑v�L�k�A�즴Vow��Y����[d�Ɇ��[����u'�<��]E�n������'-��wo�O�/p�%5�:�1���N�OW����������O�x�{���e^J/$��>�
�Դ<凗��F�3gΜ9s�̙3gΜ9s�̙3g7����g����ߎ����$5cI ���+��о}��t���Ҩ��bgI��Hf��R[�:N+Æ���o{���>��g�{��)�)��Ѫ�I���,GV�w��t
�L��Ȓ�|�EY,��QF�����T��ɔVM$n��tԊ�yd�� -��"5�餶f� �m���Sk��B�|�L��ﺺA��y��yq��VILX�n�	Ѩ��h�"}*&:*R��U��"Y-��8�*��j3ȑU>_����O�sV1u>;����h��Pd���)�Llں%H���t��g*��O�lJ�����ܧ$�W��y�z�;��@ͽ�G��I��N��"���G���~W5�*|#->B�7�~�>F��ړ�m��U���L�u;?�z!)��N �=�ۋ<��8^<�on���7}xN��<փ�6��9�������U�s�8�������S��a���SD�	D3����I�N��U����L�!����=�k�qL��Qyv|<t����:�f��9�$?;���*qԢ�;
Z&��O�,?7�Џi �'h|�R�˻AI�k�������j�n6"z���j�k�P���Y��.�y��Mc���'�H����<.a������>�C;?��1�	�l񥽱H>��'B�5_�� ѧo=|��g�<F3�_���g��ϥ�)ag]�ђ5��l�~�]�b�/�a����}Μ9s�̙3gΜ9s�̙3gΜ��|���sE��V���cXC��KX�j��� ����CO-$j�H���cA�����>��pF7���E�?��W�
�.j?%��};��=�E�_{�U�p��%�Xm�p��Q��Z8�f��vy�����_� �7����Qi�๘8u��9^�BH"V"�D�C�� �r�ҙf�K@"^�4	�4I�ϵ!WuI.�QFۜ��h>�΄�_װ��E4��R,�Η����]OZ��Y�H��r�A�pC��t,�ulMJ{�f�9N�v����d#�A����,����=��I�:�ck�Yf�EE���>�oG	��99�k�ǋ}V�d�モ�VŶ���E���R��%�%2��֖6�)�ʫ(�l�"��x�E^i��ej�I��hFVu����r�x��}~ϟ)�r�.L�}�,�{a+ׯ�ё1�ѱt�25Ff��V��^ff��������lպuA�֏K�Z����U���I�ݧ�������j�ZHS��f;P�랁A旤%����sS����T?]`��=
BL�~Q��'����RT4��ڭ�CD������9����w�w�n��贡�_�9��Z%�"���e�����"�˕h����ǘ|E���5�v�kV��90�X6��0,�IjxVT���_��3������)g3Rų/d��aA��R>�c�Òo�2���_��v�Z|NxM�k��XkJ.7�Oc�i��Z��7�,�|t��k��o4"���j���)Tm�.*$�&.Q�ylC�֛��<�/��[;y�^S�u/s>�f��{}�����u�;�R��ν�v�P�^O�(l�	̚!�`g�C[�R�6��@��^E�\�{�����3�>gΜ9s�̙3gΜ9s�̙3g�nK��FK�D�Gi����
�D��h��4�����FEa0L퟾4�fp��5 0.�c�rq�¯�گ�7���A��#��s�]�I��"��jO�m��RE�=�uɢ0�1_���c'����D�h�a���'>�Ɛɿф
N��z�^sf�J֙�2��a����#�k\�	K �����"r�$�J�b(?���Z�*)/��^���� �
E���3�~Gח��G�-/&z���w�@0*��qxD�B�>$����u� �IĨ����D��9ZP(����e�6 �(O�<Q"��Sa��0�MZ�}��ij��|�$rI�^*��J����PO�H`�`�}�/�������~f�E�Q�Z�c��A:9�q�����'ʣ��jm��K�w �n��R1�d�|u�8&��Y��8�v%�8�53>���W
���oEy�ꄦHo��=�3?��q���Ɋl���d+i�u�,ۺ�� }�^����'�#�vY!�W�)*/��q˦ }��bw���928����ր�,O�Mנew����$��V����8JO�@����	�����PC4����A�P�eq���W�H�$uU�TRQ�I�A������Y i��O�N�GD��Yi�����g��d<�����}����E⯮�g¦7�xO�҈��� M�R��v	C�x��um]�[^壵���DD����e�J�(�2�3?�^c�>�"�۵��y��a��M~��z��$�t_�49��ǫo-���7c�n����W���_��x\��M�.l}m��e��tF�qFꚶ:L��MH�e��z�	��v�e:�b5^��ō7������G���Y���c"܎4o�z��ha�߇��|�JdY�c��N�evr䒘��7|������Zϱ{�~�~�7�x�����l�ݱa�F�OӔ��~b�	"�I���Gj��_kǚ=-cZ�D�#��9s�̙3gΜ9s�̙3gΜ9�	,��W�6F҇�Z�5㗰�8�+����gy~��!Ic��N�{gc# i����Kg��9è�/��r�>��c����X�W�����u;����M��H;�����S�X�Ƀ�P�I�\�6�3���gi�EEd��N�Lk�y$H<��-�Z�X�\H����,5ѦA~�2 P֮Z�����=&"�xZ�X��R��5̒t�3��y�8H�*�W���l��&���9	Lm-����{��0UH�%I�� |�����C9׍B���ZqʿO1O"._��G�p�d��(��hJ�����,���'L�da�OWʯ(��G�1&")�єa���.EE��"��
�������^<Bj`%�E�Ii�t9T��6�R�����V���h�s�q����I�Y#����̳~��z��\@9D���I�h{T�3[K0I�kn
d]����mI���x;�o Y�q�z|�z��������A}ȳy�j���$������.��Ÿ��;o����A:}Z"�N��֝;�;F���r�?�����w�֢����O��4���_@{Yq�/��#A�f�U��Q`8O����В뢇u�����|�w��Ē}"q�������%8N��T;Q���%F�݌n܏��}�� ��V��2λ��r�Z��D���K����YX����e��}� L��g~f�.�����N�����'`x"�E�S��Iz:�;��k�EK%�␾&�b߳��v r:i#��y4�57M�nK��~]j�6-��V�lMA[CW;D"�r�w�~o~q�E��p{�kƑo��/��6*�!%j�0�-j����&6o�yw�l����Z��L�L�FHW���Zi'^'��}�6��kr3��{�V��Z�7H��a�*�cK�Ү�X�X]#I�����'s���۾�g?͎	�I��� �)�x�0����Ssܑr�_�9o���� _}�� ?��
� ��Ą���#Ø/��a]KZy^�X���/a~:����F�a"���c�7������v�y����̙3gΜ9s�̙3gΜ9s���M`�D�YJ�'4ՃC����m�NDE]�/��X�O)j�m �qx�h����]�=�g������������ �ut%>�f;��_<��QCj��ۂt��J���ֆ=�&J%�.�̇Ə�B	�O��F����ݱA�����x�,���е�ڶH�F�9�8Q��)2��/��A��h��y�`<���T�|Җ�d�"E���^�T���3�v��ϼ�l�Δ@�)��,I�n�U�^Ux����she�ݏ��2ɤl��yH��n��GI�H�QS+׃���� =p��p�K � ʊ$�RI��RR�^ԛ�7�/��"���WGe��9�����v&�i�&q��ǿ�r�$�Hb�YZ�$%^y�� }}7R�H���.$��>�/��zT]~����0���j5�I�ރrSc���\ы��Y�b�n}lO�g�g��J��I�|�gO��ڝ4�L*](PG��<}�n�L�If4��p�����>���A�z �پ�A�uu⺳sh��@*�պAh�HCOڅ	j�冨Q����A�u��h��ُ�t�$��)���^\��$⊵��Ȼ�g���KϠ&�<�����[��۾ik�>��^��Zse�y�_���k�{��W����� ����������"��5^G�]KC�T)�r�z�^2�Fb��8�"q������+@0V����� g������~��Ч����}�˧�����k$���pg�!_��V��e,B*�{�g�~m׏�,�f&�y*�>�Z�����x�M��־i� �";L�|�����&�8�Oڡqb����~R�8gg�E��(?Q�.F���td�,�Q�����h���+J�Ɛ�-kJ.v�e���O���^�p��VQw�4�۬��z}�lש�^s��8b�׮���Fۍ+��EY�j1�f?{+�!��C�&x'I�m�L��ǌ�+���V��PFzj������yO�>�ㆰ�%��,+{��c��կ_��{�0�^��]"���W'9cvT�>�i�P��	8���:5{�~���o����
e��<�铎�s�̙3gΜ9s�̙3gΜ9s���3���Y�DJ�LLCCoz�>!fo���WE|�Ê�
j�:u,H��@�tQs�L�g�"���o~3H����ijm}X�f���P�gȓs �>������&�U��ߗ��/�Gi��m.�h�ً�}M�|E���0#Nu���gKQPE�e� ����� �6݅��:�Y�<��ɨ�iG"�D�L�q2Mk��(�.���] �^�ͱ[�܋��v�0�U��d
��bT�y�M����g���Vj�Id�&@&u���W�)��W�QPW0:��@T�O�?���AZd��q'�I�I3Я�=�5?�.ˌZ��^5�z�	޶�b?�ş���?����_$�Tb}�~W��x�����A����� �s�]��~���>�2�x�����V����ai�Q�L�ݧ?�� }���t�846������/�l��,��Rd?/�|����o@[��y���9i5���vta�����:5	bU�K䍤4Uw�&�ɟ���%j΍��{����B�PԪN�����a!&hS�̳_���Ǫ!���$�����{�I��A⿣���zz�O-Bi��fq��n�'H7� �Y�C�}�uj�1�C# 2+$ٲ�/57w�یr�t��H�]�v���Ǒ�y�5i^ZZcwҊN��Ɓ"åU�OY�[���c�-A�a�e~�cni�����֍�_��u�}�ud�Quw����қh	Eg=O���?:Ă��e�RV�Xz�������ej�E/��c��Gmo1$_<���,W�z����D���k��8��|�zM�SC �g�"�G�h�����5��:��Ӊ𓦬r��KWQ���ٚL^�vk�dC�$^����|�n�����]�p�g�����^/��F%ؼ�xm��jf˥-�\�k�W�˥��v�c�A������!-���waj����_,�}��ts����ǟy�w�H�?���W�o-�����c�������F��Z��'��ؑ��D� w��X��?!M���i��a����˳X��t�h�[����рJ��K��6G�9s�̙3gΜ9s�̙3gΜ9sv�Y�S4�4�c\QL*�nd�T+�+�%�$��h���YEo7���kA�L�;�ҊZ�eS��y�K�Zf������{� �fՍ�\+�um!X�Q��=߽��-ھ���$�?W�qy�Zp)���$��d�us_+�φ�:_-a-m�(f��)K��Y����S�p+����[	A��]��:���H�<5�ΜA����(_���{Qr�6B+붭 d��Q���(��O�Xs藞�
"�G4ie**��-��l]��V%9�I���?�&Ӄ�H���O�$ڥqxtnY2��QH_xZd3�JO�����т�� M�*]�����LQk�$_����}���E�c�=�� }���t��F�V�Ω9���?�q����kA���g����g�p��_��TI���Ϥ�e{U��Ʊ�gPO�[��z�u5ȪO�� �8��q�=�^Ҵ��# �e��3�@��s��<q��_����_���]�G��Rd4�a���s`�Қ�{���]�*�/V��ax���Q��SH5]Zr���z��w��-�|�t檳��}�,<��/�+��)�0_?�~��;к�9�㸚')^�g$��%�!B�7��ܹ	��)��C2�X�!ѷj��!��P�7C�o�H�50��r�'O?��|D�<�i����j�PCr�i�xG���I&�t�^r>�9J�&֍���9ksB3$���� �^@{Lp�P��8�>H�^��w���象�Iئ�Ҽ��r�94+�"�������zd-ʑ�aT��b�?�!�6�W�R>8�����
��B�ڥV{�b�qf�|F+P�E��c��sy>�:�ўg�/3_�4�g"���"�ͅ�� M���'��V8�J{R�)����,E4��l"�[��&3l-?�ͦ��V'k�;>��";��&��f+����:�u�,�1��r;q��H\n��l�ho8�h��?�D�Fi�4���s>��$ۯωw��훷�����)�Ԃ���{���-M���Jٽ��[�gA��؉�ݝ�P}���G8/��}�r��o^�����{��	����K5?�'�ӛT2���fA�|��s�̙3gΜ9s�̙3gΜ9s��&0�Зf؏4��AZY\Y� aw��mn���I.q%X$Z�+�Ҏ� ٲi-<���X9���3��(�?���i�5������?�g�<H��&x���J$H�]�����A:~
�Î];�4ɥ[I�M=���?�gf�E�O�Q8���>�r4]]7�C�U�bо��=F�H�Mf<-���p=,�j�S��C�j}�pIS��D���yY$�V�E{�x4��� �E��I��Z��^�$�T��*[=�h����c>��F=&'�/��檲�i��cQ4�T��Nh N��ga����X�|�#t�4�g���P�\���r,���� vg�AZ�yZ��e�?�2�(ǵʛ����+�2����y܇T	�����[8�e'o��j�~�кS��gq�N�A?I�:C� X~���|�駂���N�޽�iO�B0�CM8$>�ڔo#a��gi�]f��Fb�O���@{���Az��� �Ƚ��z��[X_��&@.ʳTe;�;�l��K����~�=j�I������ٮ�'�*F���D_��FQ��"����I���Y�����j�j�#��{���m�=��y������(OW�.��+q��ş���7 ����/Qf��ݽ����� �h���CV��uE ΐ�%���+A�����E(�ދ�L��78�~��j}��wqz��G���5蟧��X={�X��I���KQzQ�I�G�yw��C�^^|�Kg�.�ܽ׹�v�C�ڊs$�I��?����t��E2�T��H���4�z{��r�0��(5���������i���J��׎k}��Ik��0���M����L�yޑL��MQs����K�==Om�w�]���s������j�?fW����|;�&�6����=�r]+�ϋ��47����8�����ۑ�Ę�~�5��lqVm5j�e���4�ZU�=c[�~�c}�w4�v��'�b���ϯ�n��]n�%���/�q|Id��f���2�o�)��D�k\Q���4�\ug1/�A�7����<�7�_�{WO���b]h�f���׬8��.^�{�o��
R7��;8����v����[�u*C�Y$<k�2�5�|�����Y]#�<�gx|C�i'��"2�.���nj����}Μ9s�̙3gΜ9s�̙3gΜ�f�:XQ̊��$P]����b|h�`��� ͢�} ��Id�+z�p/H�۶a���װ��`��O~�A��@
�IV<��A�b�W��W�W�6[�[
o͓Uk��u	��ݧ���S��+�틟��Rm�{[�@P��5����IU�}�����J�ĳ�>s��zx�(���op�V���+�s*�t~�y� ]��)jM~�/�U�[iY��O�i�q4���IɳG~8H'�������V4RY�QJ��Cb�я|��a3DbPQ2GG�w����t��[KK)C䡇Uu��'خ�����ǂ�� �G��<�Ҫ����`�I$UIZv%1N���� ݱ?~����Ꮳ���A>��֟��������n�yy� }��3"O�z�ٙO���Fia�W�#�[JLEx%��U�P����w�$T���3?��;���䏃���Ӽ	k��}��4=�8�(���uy��g�@�����S�$��gHD6��85ږ�=�a�ю{����A�n�����O������V�&b��dא���.p��\�[��M\ٚ`���[q?���eD�lB+&X�Obt�뮧f��~x�4N+zs�0��w~�4�;~"t=�"f?r?H�A�ݽ�[�����α�/���|��)�n*��J�4�~��xNocT��GǙO���IVIнJ���GP�陙��zzQ�O<�� ��c�	���3A�qm����@{��g���0`4��z�?����E4B��I�3E#�|���8kFbD�]k��D[U[i��9k� �ig��!��&�l�*�E��U5�|2t��������'����'@<ws<)q��k4�2ng�=��-M��?�O����&�T�F��O����:�(4o��eT��醿��?j��k���1da��c�'���}�H�%k����H����"���n��=/S���Qk�_4���3�<���/>tQ���tq�N���d���s���އ��Gva����������>���O=�����'>�
�|8}���w��gӺM��E���������_��<晹^����[��=b�;�n�;/�èN�����5O��w��4��.�S9�ץ�X_ ��^����<:ŝ�=�}�l�~��̙3gΜ9s�̙3gΜ9s���M`&�G�>FcQtN� \aL1턇��cX��p'<�����)���J.�ɝ$���Xy~�D�<Y�
��ZD/\3���Q�:O>�� �3J�?����IQk-~�	���������o}Q]!1KR�D�/`�������IV���l�!h�e���[���n|>��hi��ω����X�y�
�5�&�%��(�@����+�"\��|�z�1����a���.W����N΀�x���� �s��.i+�ԩU����Aͼ5l��HaJl��%�@��QW�e�_�[Dg �E�Pڑ*G��DD�g�4;v@�a�Q9W��J�m�$�-M(��*��Ii\����4�h��M�c{1�l� 2j��R�Mp+��608��'m�cGA~ud����{�8���.h��d4*��E!V�D2<^JNZx",��yY;�(U��f�>B"q�ڋO?B�����0����1��o�v���ڶ	�v�ĸ�y�K��,k���NG��7Q�YO���X���$rq�����e��\���������g�A,�q���]�<t��� \wl�v�]w�:E�ӊȹ>�INk��˱�$iv�N�?���O}�Q�W�4��7A�NM��̒�ˡ��<�� o�	��[@8�Gb�D7�F�;Q��D�jQ�h�5>_���9��;��x�Q�k�R+�Gi�~�O���ӓ��9���|����]E�n�Qd�U|l�|�(�c���/�8i7&X�4�=�j1�x�|�F��:������%j%�q�pC�"bFq���`1$�E�o����>��M�V���F���ȾV�ei�V�z��7����]����'2P���Ȋ脢�aUK+�����%�k��݊��|&E"6V�,��h�<����ט�;o�Q{[�O�$_3���7L��CG~5�?q����c���~��-���oV;���ZݏY]f���i�i���s��=o����ڑ�I���ur��|��Q3��G�c�G��|��=AZY���vR	a�p16��rWV���5"�U���Ǝ�_��_�����jh�\��I�n�{c|oټ	��3?m�^���_�ߟ���{�;�X�	/�yU85}z�e:�Y���l�D_"�lh��>gΜ9s�̙3gΜ9s�̙3g�nKi���v#9x�O�b��ȕ^m��$���~�a5�l��К4�RZQ$�T^��T��PO+����S���k�@�)��~?4���t�8��^x�gﾋh���w�K���C鬖LW@-�W{����+�'�ae��g�҃$R6rE��Ǟ`y��ڒ��,���U5�Ѿ�4k��I���6"hWC�U�)����W���Q5�_�N5���7�@���f��=��GDV&��ۅ~�\o��F�t<O�D����" y�V�-���� ��9���$��]MD�H��b���y;�}Ub4Pi�������Y.��r���Dzu2L>��Q�k�JF%�� K	_Q��0�#r����P{�֮�y�?
s c׭a�� �lvvຝ��,���U��!�c	����+7���v���5[F�!L��g�X.E�D{��HZ]c+�B����-H����$�Ǆ��y�p��^y�	jHm^	�������l�i�$r+$��t?ҀK1�߁�g<|�����
�7��W���q���cH-*i!���[�E��ۏ玢`)*���:h�Y���e�Bl�����ĸ�i%��;���oل�ڛ7#�G���9x��^4��" ���d�8~�X��������My����:	���I�C�����+���j<w�ue�i���.��W^��V�=44:NfGO����kA��G?��׀�+��?��Or'��?�<��/u��K8��yeۧ����M�S$; �x��bErV��L&��96�t��f$_8?uV����уl#�ƃ�??܎�f�O���~�c6�v9ַ.t�������_3-�����I�{�e W���AΗ����v�����o�׾y^����糢_�fj���!I:�	YX-�E׷HQ��l����nK���`��¿���ڛ����f`��2����׍!e?,����m������@{g�ճ+����z�Z�Ml�Za��;!���C����y�Pü�{�<�?���4���$���R����=�
����c^��ǰ����2>����Ό3�Z��|����W�`G��泹�C%n��D�%~Q.k�~o��׿�_����@�'��p��Uxo�u��}|��n�O��i�����}Q%�w*��-/��yv��tV���|����'9��{P���c7ҍ�d���[�G�9s�̙3gΜ9s�̙3gΜ9sv�!���7B��#�S�J#����	a㊱Ȳ/?�S��+��J�#��J�E����$�~D����� &g@�m��1��3}��� =?b������� ?����g?��!2��vel�8E�y��Az��^�΃��u�� }����fW9�Lw9�����0�ZI9�Cyx��gS��WХY���K�հ֌�)�=̵&��:��(���{�֢�8���̪�^=�Ǚ������E�<�XJU��`�h��fco?<'�ٳ<��v�!3l�d����W��'�1T�}�#)�G"�ƿf�WO7<#�MH$TA$�b=T��RQ�G����Qz8(v���ӑMK�	�+*��.�}��=^�!Ϡ�)�2z���Ɏ�ᥘ�p}�1�ch�`���
��F���	��<ۙ5j���l����c��q��'��Dj�=XA�3��KdH�v���H4����.�t]�,�8Տ4�Dbg����
In͆F@��;m�AF���6�<r�_�M�"F�c��'�h["��v�E��\���ކ��� <jF3���P�N�{K����9�~�K2֯������;^���q��˳�E5��9G-�YF���N�8�WZq"㵿P�)zvg���I�­$cW2j�)��3�8>3���SK�6����gY>�0Cfr�w�f��*�H���0�?��OR{P;쨻�9h?��n�����v����}�q�	�}-.�F7��A�4Da"��c�td|��K�Z2�"|��.��8����D�����^?����$$�R�F'�"���g-�ņ��r;_�-����!�G��mmj`.Wv"�q��S�q���lx�&�Ʃi�m��*���:�bOy�S
������Kx?z� ��޷�ڞN���sT��s<���I���0/��c_�?{�O����a�:�ڹ��;�.������5��{0�c��z������c*�	����<y�w��G?�Q�j���<�=x����xO]�|HC{�����9�\Ks�K�3�S��=�Ɋ$�^~�� ��X���8OL���"��t�=E�O���q�KW�?&�c�`�J�we�����w��̙3gΜ9s�̙3gΜ9s���M`��+Q�_�� ��)��Η�V�%&����؉�˃�����4�v�D�Ǥ�B,����$+ X:�X)�c��~h��
VDO���Qj��5�����%s�8������ �E2��{�p�:���<���X�
�W��g@@��p� �?�<��+�"I��F>W�D�?�9��I��h��X�&oP!����^��>����4W����^�1��f�3�Ǭ�Q���=��$����,�)d%8֚y��L��"-�#���J~$�%s�8<~Q(mr�φ	�$=]�$x�H�LN��K�=)
e��D���"��i�HJ��*P�k����a$�/k�.y��T��W�M&�щ� �1�5�Ԇ�'Ŗlɐ'��"�Fn\�!H;H�ř�g�ʿ��ʓ�#)e�4VIS�����&T%����%R?��&���2ځƧ�+;��^}�P����զgV$L&E��"���Xft��GW�0���	ܗ��5��][`�uU��S�W����Cti��*��K�H��-(�5MZ'�L�B9}[Zlv4㩩p��>jh^�A}�NK�Q�[�ġ4��� ��_u�����aW���gKr�Շ?y�Q�4NK{2_D�K��҆L��m����5a�L��@c4~B�������屣<���z=����]^j<0D�Ph���"V���+�+��.�cGϦ�Jvؚv�����8�Ķu?"�f�z���lv�|Ɣ#��6����r��u�V�y��+�e��T�#�afǊ�h2��-��Š��Q76��hkJ /Y��y{���Z��\����]}��7����L����y��=�ʏ�t�����^�>j'Ui��wX�5�@�}��/���`]�,���\��c^��ɝ&�q�={��u�x��sO7	��_��V���Sx�;(3��[�E;X�m�N&i�^�u�,筩4*��[������j���g9o7;�����D���@ͽ7�B3��Q�o{V���2�)kH>�_���D��J���?=���"����|�&8_7Z���s�̙3gΜ9s�̙3gΜ9s��1�Ч������E��DB��Y��@i��(V_ً�[W�:>�h 1d�<��*V��><�+�Af<���A�̳?��G�����J�;��ү3���G��|��������nD�\XʇH�2I��^D{[1���>Ϳ;?�zz�=�y߽����/}	+�~Y{�a�<�� `5i��b��o��
҉<Ȓ�aF���y��D���3���+چ�#`G�1bG	���f\%�����FGj٘!:�Ԡ��#�P���Ⱥ#G��:��_�蓶��X[����A��L�Ag?H.�"�R��U���*Q#��4�|ϒL�-��8q	��Dk�`u�o��d�ˤ������I�b^&j��iEc�kU"M2���0n�[��b�����{�	�6NSorr2HEjNR{,��HXF�C����G�.�/��K���z� Ay���֭[����5��V;C���E�U�-��:�@�]�ڍo�H~<y��7H�Fi<*���g�!��1���2*�ڇ<z�6[c{��xZ䌈9OZ3�R�h�g�£�h�"�WR��hr���a��M[D���8iu�����sJݾT]'6h"�/�,�0?E��ĺ<���8�4Q�ˡ|ף/�����b;XK�i"����MЃy�Q��$_cB�ք,0��MA)� ���2��ĒW��lsb���k�"����x�/Nc�:J�]��W-�Ǖ�Z�'���ڴj��Ѩ��y�h�ٚ���"�7�}-��k�nV4Jv��W�6���<K���϶�t��-��7�5%�bƝ��hZ]��w��KM�~��M�q���k�]���x��v`JCX���^}>H׮Z��itځb�t��^��ĲH�o����b4|��gH��_���EjЍ�v��xܿD�˯�Л�Ĩ��AT��:�y�1Q}9/�|r�F�ow����V����o3�9�KB��v�Ƶ �z��^�Ǽ���c��G6f�s�����N��������V����3�w��\/���(��j����G�;w�mowtG�9s�̙3gΜ9s�̙3gΜ9sv�Y�3+�y�`&�b�����VE����m��I�g�CT�{6Qk�ZC��4��K�uRV!ٗ���D�G�~ H�dA \��J��I� �� p6n�
��ɳ�޻�w�W��	�i�eڣ-����]�
+�9��rE��9D{|�]��ڻ����� �r�F�L�`��\"�+�,m>O�$���V��5�%mb�k�1G��".���>-��d+���j*���E�m�@�?��V�ٿ�sD5sP5�|��{�����<���z�nڴ	���h�<��B��Q��׿��<�\!���w��u�~�8��O������͛���G��#���nDݲ�y�x~D��3:���;��Hd�떶`�a~Eh(*p�\ L"�L����� ���[�Q����y�6&��#G@�%����-m����K$E&�� �U���N��T5Z�"f,"�8`9���.c��a9��X+����@2���y{�a��YF�M5\G�HĔ�ٲ��V�@&|::��c;9&m�s�P�,ɼJ��d�a�fK��O��"��_ q�e�V�4:��Ez����L����	�߷0�����i�g���E�q��,r��0³o��;y��v7߲�c���\������8�t�^<�|�� =y䞢�X���7�R����vX��h�\_"���Pt��qx\E���ƍ�Tc�	Q���=��H<��9���xn����i��=;eY���ѷ2�HG����.r��ۢ�����������ɠX��Z�Q1d[]�1�dU��f���~��Y���B㾾GW�� ||��j�ő��4�jM���'P����j����e�hj��5��@�jymm7��M��"���j�F���(��%��i�[��y��K���T������}N�!����h/�<{}���+I,@�2�6k�������E��c���ǰ���^��a~?˝��Y�g� ϭ�{��8�`��%�g���� �K���u��Y_����`ټ��[o�{��u ��s����$�͐|8�Y��$��t�|� �s��h�ݜ��
�
�t�����b}g�q�a:u�5>��6�ڈ|j)/f��#��9s�̙3gΜ9s�̙3gΜ9�	,�Ч�ܷ�G��폀�;_��/�u���$r:�9������z?I���4ȧ5�Ғᥥ�g;ԓ��*" ��[�a%v�jH��X�=|�ҩ� ~��6߁�<?VD�\�����cȗ���EFQ�p����$�]��� I�U� <F��p�/��t�.y$���2�K,���(6���.�|�=�V�8c^�G'�BQ"k5����#QsY�����0�<��!'m.[�j{�����y*�gj�5��ʴ���J�ʷ�*���iIEڷ�N7��Jl_w�~G���ݶZS$�d�R*S�e��69b�Uo��~y�\g�������0;��ѣ�G�6+� ��g�g�����=���wq������>K󋄅4��A������k��K3�^z�ӧ��X��~�q�0�02J��iF:s�4����ƛ��|�+�ɾ]wa��� j�>��,ƥ�^jd�l�Vݪ��г����4}������!�����Yx���u���Ҝ�0
����E���QFoްD�/>�U<�fq�I���hμm|�ڿ�y�Ѧ==��r�}�8x�ܙP=�q�ݶQ������}��p��.�	{���]h���[X��G:L
�j��ih�X$���� ���F�����$���{���W�.�R�3�q��$��
����g?��HK;E���x��*5��4���QE�.��W��"Zw���S�{��Z �H�9��wtb��s��ڕ"aU�/|�Az��q���������njٖ��Wa��G�D���/�i[.� 3C�P�=2���֘؈�~W�4hL�5;>�m��>Qa��)(n�Zu��a���w��M�x-�Ru��ڟQ��|u����V�L��l��n}�j{^%k�d��˯|���7m}�[���L>$�U3�j��h��XQ���y��g����cwѨ}�?K��ߖ+������S���&M}�}
����� ݼ���~�������Fs�w��N��kb����>���;�����1h��8���y�LW�s)��R�����f<Σ���EK{�Z��/#����������}����S{Mf��fyA|%�S	̇_�zў#�)�1�y�4�DԚ�ί�������$ׯf.�=u���#���d8�֍wD�3gΜ9s�̙3gΜ9s�̙3g7�E4�D����'>���]͊��O�� *��H0Jaj �/�c��?D���t�n[�=�������@+Ǖ2ί�Ռ��Q�k��7	�� g�ΐP:}DH_?���1Z�5?���{Allx+�c+F�L�՞�==ub��xZ��n5���#��ϟ2H_~DI�h��3�5f)��56��G\�p�m��}����9��k�\Q��E�����NY���e20�"�(φH���~�IMM�4��_�Fc������Z�dj���� ��:H
���Ժ�m�mAz�hT5�^��S(��G3Q^��Hྷ���$H����u���)���$��]�巿���d�<)}c��M詿�>�D�������¤�ڋ4�U$ЫoA�/��g��h����^]I���Qx�.]���އ��)�������_
�� ��
�l�Qh��"��4����$Y��_���H���q��}$�C$�� �x��� �|	�覶����>��O�ix�Q��h?z	ZUj�&I����p1݁.~�-?�G��b*N}k�@Q��0�"��b5X�����zU{[C��_�9����c$����+�mW;���HfE�Ԉ+�S ��_D�!ѷ��W������D���BOZ�3$3W������{�v����ۃ����U��~?Hm��W�iӮDT"�sQ�g/��#w£�ۇ�+����[������?
�zp���I�Cd_7�=E���K�'"��Q//�-ƹ�C��,݉�r�"MkV{4�x�]���Uɪ���G^DH���Β���T��j�F���A�am��h��ב�_�hͶ�^cC5�z3�;Nfč�&�b�E5���К!�����0/f\Y�Eƛ��̖���>����T��yqLs����q�ڧ?�w��Eߟ�����ߢ�W���z�m������5#��;��=�#�S�畴��2ɾ�<vF>��?�(��]����L���b-TC�+*l�����؇��w�}d+v䜽 ��S�?�P�}r
�Y�����=VX���y���=�����h��GC|/�uv������~/��h�M�����ؙ����Q~�|������	��*�����\^������MxO�I�:"�bڧ#��9s�̙3gΜ9s�̙3gΜ9�	,�Ч�d+����� &f5ED�<J"�b����I�H�?�ޟ��y<Hw�Gԓ\����V6��j�a$�HLy� J֒��tg�ҙc:L�b�����%Msd+�qѡ��=�H�%��&z0W�k\ѭ*�(OTN�yz~��o�# <r#Xѭx�Ѕ,ə���8<Zs�=$W��(�\q6d�8x��YdҪE����h�F+&��e��Xwsߕֳ��R勏��H�n��37��4I����?E �Ҋ2FW"�uv�X�?t
d�S��3�Ȅ	8i�i�?�X����7�C+K�_xZa���`�!KBj��b�������D9/�q������*=�5��oI�ˡh�a��E��b	�p�H�'ͺ�˨��
��;�����F۽u��P�L��#�1��5���|/H��4�=��L���ø�΂DRtZcVT��ڕߋq�������I�������A�����A�P����ej:v�c��G+ً|����AZLa��p�S�]�Ov�,��H8Њ�i�����x -����۪[�\ǿ�&���<�� Udi�>P�ۆ��tp ���S����@�V!�g�w,8$���L����v�����B�Z]��ȿ�+�=(�W���	h�>���A:5����'A���G��Ǒ��4?�}"^��T�H�0�-�c��>OW@t~�e����� ]����?$��G�G��Z}_��O�¤���9����"�t�0���AT�;nҷv�L}�h��2*��h?�Զ�v˚<���َ����i�]3�6�R��M�8-���e<�1����U-|���z�[䞾7�*f�C�Hj��k�=G������aW��H�fZ}u��fhP��Z�yjS�$�2Ϸ�9k~�E�X�5.X��{x��ǐ��[����]k�.�z�d����rq�K~n��@��y�f��\�;�d��,�<�~�t ��+�����|mu�mm�y�I���z��y�������5�؉��I����lym�!�2�n�HI�c`-柕�H�|~�IcZ;Y�NiR�z^��3�8����T��_�7�K$��Ɍz<�u�%�{��y�S/�����S=80ɝ�~�"�·�V�$I�z�]}Y�+L]�������`���z�W2G�9s�̙3gΜ9s�̙3gΜ9svX���^�w�<V�Qfw����,C#��(�uҌ+�:1ɂt/Ȏ�,V"����f
ؓ������"�����E��<��l���U�}5��l��^Y���i�����0���Λ�4�|�|��U�'�����ǃ���@������I>PI262��X��XR�Eό<��h`yE^�|5�P����H�N�D��uLt�0B�{�(8��?�8�xb㎓� �w����x)HKȦ��� ������O�����>�>q%[S�gĔ��)��W���Է�4��P�!��t���х�"�2ɷ*�_G����|��G{Aڌ�@���u�u�R���<���w0
�4�|���"���K��j��;E.I�N���J����C;��(�K®���{oA{�\�����ޏC�.M ��a���1hG̑8����*�L���F{Hwg��[��:j��,�_ӝ�]�or�u�"�����_z���nh���L^�V���Jn	@�C;�}��7��O��R�R� IK����*�b�~WX��ET&���yˌJk���c�_�m��_�]���%�\�r)��5��կ�ʕ��뤦����ڹ+HM����ٮ����u���P�#R_�����t}U<j�2��L��_�������A:�}���:K���_<MbOQtU��[A4޺ڐ��l�������ct���p��?���n`H�ǡ!:��x���&���A����o�j\�W~�W���= Z��/�2�A��ħ��Ũý}�?|���ڼf�����;��0.��x����Wc$�)�a�{���8O{$j��k��ϣ�͖
�h�d��4����kv?�����v���sЏx���p����bH��<��d8�^Lk"k�1�y�l�Lt��Mu %-i�z��j-}��i�,>�st.R/��qիyВ�&�K-v@iq�������{����m�劜&�H���M����g�*�綵�̸W�W+^���l-���|7!u�:�~~i�-�O�g�����a�O}�뺡�<@�j���E�E&ء�w���� ?*�n7�s�q�:k��+�w�_'����h��B���ƛ<�m
����W�B��r��.|8.)M��AC��Ρ'�>g{b�ڍAz�}��[��{�����nb��s�̙3gΜ9s�̙3gΜ9s��&�Կ�_�E�hE��g���i��?w��(+ꮘ-!3F��+�~�����/�����3�:�5��$:2>��*Ds�B���d�ky~�i5�Q_��q	�+��ܳ�c�^WQ5��+^I��L$̟��[A�� ��rc$R��\����U��g<�q[����v5�#^�ʸ~_����j�ڸ���h��<�X 1�e�L��Z�$u��噏+PL=(_��lyƴ��h�}�4�O�lJu#Ͼ����n�e�1��R~$��y�&���v�jNR�.Oѽ��A��Yo�J��*?O2��o=�_Qz}F'��ߘ(��0�yn�����ir��ɏB�al���G�����f(�)�n��?KBM䗢��c)BUd_�t 	j�/�H��C�Ѳ�y�O� ���		�=�m��m�<\��Jbx~$�YF�>3���ȷ���D)�)�B*�i�Őjv*��e9�1Z⸱�F���I����SA�Н���Q���>��EFG~�y܏�G�e7WB���N��|���h0���ɖ�Z��25�*h��.��v�]�����Q�Ҷ{�>DΥ��*G�45&�o��������W����u�XU���4��R���q:�r��o�� -��U;Z�zXni|$Ú�?��������o�� ���+A�eH�[-{�hi(Jm~���E�ͦQ�}'�����ࡓ��q�Z���u3�R��y.X��<�#$�&���ף�
����u?� ��>�����@�~����F#M�u�+ij?��}�O0~<21E�����IJK���)��#Rcqd�=�&b,���ڞ�p��G�m��5{�Yj~�x@M�v����n2�F��17����D��f>�n=�{������z�h�Y$�1?n�Ų[��tծ"��Z��w�l�Ѭ~l��&d�9�U�	���,�M�jCZ$_�dU<�T��y���������f��-��,����q���2Y��7��b�����5&��iG1��z��\�G��jM����o};�n�<��[��h��sSUi(�3��Q|^���j��f�w��
�*xm����S^f���}��-���q�4/��2����jN�z��:Ң�<]��i�32�Wd�!(-Ĺ�x�Υ1o�}w2%�^�FϪ_���#��9s�̙3gΜ9s�̙3gΜ9�	,u`���/L00z.� !��h @��� 	3�S)E×f_X�JB��h}@E�NM ��7����#���)����M�K�Ik�w}�]�Ax��%O��}�
3Wj�G+���T���1j�o����9D�����σDY��Jn�$c�{�k	�x���9��B��5`��լ�rC&�>F�c4�*7�W���	.U$AP�_c�H*!2�d��]�\�r�D�V�D�ȒNj�I#rv��4���˒,�oH1�3J.%����P[Oc���� �j����3���d��i����)j�I���Y���y��~�ui�IEF� Q�')X^@��'����҈��?����Nڄ�Ƀ�B~
�HEϝ��~�s��{�@eR��c�(�1n�� �
�Կ��=�*l�Dx��-ϣ�NM�c��D��� �jԮ+橭�
��P��B/|9c"֔*j��S�����,���-Z�q������xD���$��~�e��� �~᧿���7�V� �W�Q�ElJK����A���|�ڱ��D{.uPc��y"�[��A�RѿE��������_����:����z,H׌"�s>�������~�'O�q���Sа[y�\��b��m�Z����P9��v�5R���n�9�a���<�٥2�ɷ~�\������w0�zOY������Al>�}Di�qܙ��c�d���s��wi��af�ʰ)@-�.0�5_�v��*^����k��_���ȣȎ�Zk�K�Qz��'r?Lȣ^���E�:���O���[q|�����ǐ(���G�mՒ�Ģl��Uc7JU�/��8k|��F/�Kk/�^���[�X^�zX&r���ǔ��h���w�]��豰�r�z/���[�����h]���nгp4�kmm���"����{w`�8�G��vܗ>�� ݹ��)j�)��M��8J�Ϟ-DF�$��'�I��m6yo���H>�ü�oE�s5h����u���@�Z$_�C�	<�A�sJ��{0>'��3����������>3Ν/�C��s����E�5���̙3gΜ9s�̙3gΜ9s���M`�{-O����+yB�ނ��,,�S�3�m�� =Ǩ��*<�U�8zf	+�F��K��*��W�Yb�����<������Ī�MI4�n4��{��Qv��6^
�Y�Y\�C.�!_���OQKp����D}��� 7�<&�Q�<e�P�Z�J�d٥\j��
+c��ǐ|�ϑ_y�b<�	]�k��<��D�u���?�C�~��O"�J$�t>E���Ֆ�J�Y+�1��y]��QI3�$+�q�+����\���5�����z�/�a-4;߉�%l��7�h���K<�7zp2j�I{��� �7}	Q�2��@$��B���	*;:�!F�K�!�*�~�OS�L�p�d��<<3��&���d(��Ɣ�5�"ָ}&cHӮy�2�?��W$�J�?	�ay-M���:�}o���4qѭ,���X�~�hă��+shwo���� O`�Di�Z|�o6l��>�d$�N�:���O���]�c�-f9�x8on����L(þ��
���I3<���f�B���ڝo����� ��IN��*��� �.��ذ"Hg+�\#	��sV��e;��c�|v��zsEy�r����C�Dii��������3(��(�� ��[�[s%z���>��y�+����;~�x�����q��S$q˜'�W�����D܍B@\�|,�䋳�a{ZV���a��z�]]��|�D�����$�y��93ϲ4�ⴳ�Z~�Ί��o�_c��kB85?A䄋;O���i�t��b��K�1ˮ���<f��2���	���f'lv��'�'���_V���}����v5�d~3����C���mG�?]���69M��G�A��	1u�-�IFZ������\�ˎ`��呟ﾈ_�@�ݱZ.�����%V;�L����F�O��A:=9��  #�IDAT���f��z8�~?�;�t��āY� ;5����Ob��� �;1Ov�=��_;���&��9��%�yt��늲;���g�~��1�^�7�zP�,.
�#��9s�̙3gΜ9s�̙3gΜ9�	,�?�O�C���$�7��=���A��d.�&6@[ο�� }� �pְ2:_���gY�	/~�T�S"��j�]����O!�ߺU�>�e�� �}�� �%��\wĆW|��t`��x�s����DU�>$�Hg��蝗@9u,HO��r�ܩ ��d�HS{O�O�Z�9��"J���Z	�@ǟ�5�/���hx�����:��X��A�.?ׄ�kfM<�Ƴ ���)�R���,�&"���ۚ��0����z���}(��Q��)1���5P�(ʭ-א��w^��"�|C���7�ăW_*�Mp�<���#I���\(_&L������.��w#�_��k�:˓k<̼n��]��t����y�YiL@W�j?�5�6��ex���4ј�t?km	��䇄�Ϩ�jW�.j:��7�,���_��s$�2Ԁ�<Z�R*T^�n����T;L)�8NQ��giw%�U�ۭ��b�R$��YF���V,S�э�ffNi�p!TNC����G���\��8�۪���n&�!Mmԡ�Q��ѼT�y�����T��:�*ʓ�F�h�C�M�@i�K$������U�,�@�u��u������O^�y�X.j�·�ˮ���+,�lV�T-�V�X�j��ƈoTc)��f�����D�6�H�8d�cGv�I�l	ز<�V����)�g}��ku��ʏ��6Q���c�+W+����2��mGc�?�I�x�(��l>��q�f�i���K$[$�]e��h�gq;J���c~��ڶ��]�M�oz�Z}?���JD���a��ޕ�˵�c�k睭�h=�u@ˠ(��ֳ�͝G԰~��A��>�m^�1H��qg���zQZ;����
{��~[�zB�<P$"��eF��sХ�S���Ƒ�ǃ��,v�$���t��1|�L��3DZ�)��W|Ԇ�l
��N���<|�k0H'/06����;�ҕ������.hb�Z�tD�3gΜ9s�̙3gΜ9s�̙3g7�5]�Y%Ӻ7c�&��b���m����/i��F5�tV��H+�F��,�
u��Y��n�����&��W���{�ҡn��,���`�����.h� �3 :I؉(�#�t��`�����9͡3�|��^�������Vn�V`���5�0kj�Dm
����\Z��V^l6���=#�y�2o%�����z�ca��.�u mۣQ�<1V'(�yN�+'���"�j1�/�����D�CS"�+3�5�r��	=ޏ�S�{E�G��u��ʈ��x�x�,�̷�XEi�q��!��=[�-FS)BdD�`v[�Ȧw�y���GN�ʣ�����|:��3Ѭŷ*�ϪO�Ƥ���j����E�&�%��C����bN�N�����65[kD�ke��������T�d�	�e���5Ltڤ��1fR^�t(H��HȑP���a��u��"ޒ]8o�d�}����ى�ڪ���]�|}��ߪ��Az�(4���~>��p?��p�+a>i�iܜ��\�_J&�2>�#�I��f��8O�jj�����y��V�	�s'A��L�{�ĉp>�N,-��u���^���i׈p0�EC���5���V��`!�<a�3����.�x�c�y>�	@�l|���lש�,6*�5�Ef����q��1��YgY������k�ē�>�Ԯn;[�(ŉe���+nxZdu�����?h�|���ڵy��ڎf{���V�١�8��f}���wZL�D�咴憣� �>���P7ȵm��U�4G-xi�ur�&C�M��Z��1P�U�;,���i2����<w�L\�����ns�,�Q�;��a�j�ۚ�No�����E�q�!��F���_=L��$֣.��N�LR$�=A:��6�H>��m�ӎ�s�̙3gΜ9s�̙3gΜ9s��&��B_���%��JҊ�������n�����@�>�Z3UxT�kԄJR�(#��}�c�="��4���0�,`�6A)7�H$3X������]�o�cǰ���;�k~��:�i�t�֋���d>�-��虆 ��ɜ���갢������#T�l��F���{vt�&.C&���q������U�b�������L�SS���GG��:��]�|$�R�G��'����Y�\oO�a1�#�l-=z`,M;�\���"��h�����@����}���F�m�r�]�};�d�&U���LT�p9��
��7�#����L������4��&)���ʣ�#�ԌO����}��6D�:|� ���Ҧ3ڃ�6c��yV�oϐ���[�ʿg�n�ي�cT�jϫyCJ�`d9:��Q�&&*}>�<�O�ƕZ�Ԑ��'�o��i���o$�԰�P0����]4D·�����q���0ݲZ�s��ʱ>Yݥ<���*��Ο17�č������KQ�뚥ab�f�@�-΁�k��umɆVI�Xb��k5wi�I�7������ꆶ��S��Le��k���~���s�؏��t5f��vw�h�Ɓ�H����2�w��=(��uZ�]������4�-��/�pk��W�A.[{4�~u��"�]�f�!2�%�fq׳߿Z���V;���fQ�o����q��K쏶ı^�D�O�U��p�� }q?R�����|u���� v�����!̫;�Sh��>Ʊ���� ���}g�d�|��,n2M�_h'J�}��J��y3�d��Pk[1 z���;��ꕜ�w�b�ӸN_�u�� ]��N����M�ӿ���2���'��]�v��wD�3gΜ9s�̙3gΜ9s�̙3g7�E���۪���hCi��Ⱦ�}X��� ���o�9h�M.iI�%�bi!�hJV��4�:IrX���t"��jb��M!��x{= 	�|F}L�4 8��&tl�����%k��G�3��������D��t��і]d�MzarF�<[���D�S%���n��E�Q�#/rH�e��R��vA�X�C��DG��9j[v@]�Tl�й�g*�9`��6|^C��j���ڄ[�$k�Y�����I��3���%i��0�c�)� ij1c�<N+!-Rǅ5�QT��O���ۑ�j�߶��vnH[�?M?K�O���)��OOّ�{y�01f�5L���K�h���Q�=��p�ZYR��Z��s���b��O��h��j~D	K�����gϷ�q�p�E��E<�D�1-��9<6��%|�v*���;���}�H_8��,���<ۋ��M�j����^-3��5��[�Q�^��YF_���Ͽ�۷i� �����^eeF���hֵ��%���:`��n���~Cd�;�hBN�Qw�m������+�z�z~$,24���x�j4X�z�E����*�����b��}��|i�Q�l�\\��?Oآ�h\��%�9�Y����dZ��k�����e�-k��iM����|M���϶�/��������g�o�k��;���ޡ֌���`R_'h<�z��=�>�/��к������%���w���p��[����О~��;A:S�<�1j�n�8��mVZ5��H�
���b�b�S�����|�/�}ة�S�uWv!V�(��g��� ����!�n���&_�%{��WB�z衆�9�ϙ3g�_{W��q����DJr�Ny�+��*�r�%�C�n*���,U>��8��X�,Q"ERC����@�o��P2�� ���������`0��`0��B��\� J�h {����o����
��h�}���*\�qEu�̓WP���22ȋ!3L��`!C�4��sb���]d6�^�b'��S��I�JhH	�������b�i+��r�|�j	�k�bq�r�O0����̷(\mb�H��7�3�cӧ��	z��DƶN=o���Ntzm��}y���.�`TĂ�|�����3m�ƨ/�0�9D���UxԸDK��ܠd%����yc�E��������;������7V��=�'c��2���+�i��5�{J�^�@�D�"d�ª�>i��Z���'�i���)]b�b���n����z���|�~�#�O��8)�|u���;�p�|4�"���X0�K���ASe�-����M~�O��ן�v�w߀�.y�.�������O���嗘�Љ��v���S�c	��{Me�h�P��!���.ߋ�r��5eŸ��7pǛ��<���s�WR�9C���p(�uu�o>/���C��c�lf:f��}2C榉u��m@��3�%�y����b>�y�,۵w������z����^:3PC��3r�E,s�+�f��W��
b��"��r����]x�2/0m��<8��R����#��;aJq?��y�`
���7_]b|_q�| L��.��������I�������kQOF�S�!�{�[Kg9̯w����`��`���|�������= �=r�,K�����`0��`0����u7�r!;x����N��3����V@���t.�A���5��.�;+��dY�K�"F	I9e���[i��������=��N�\z^Q&�`��H��Pz�r`~E�V_�?��pś#43�Jq��7��P���=\Q���B�\x��0�13��j����Y\Cz�9��(�9(�j�j/5	B�R�����^h��t�H�X�M��Y,U�R����T˖��T
 ����i2�V���ߍ������G��*��C缴dJ'��C�w�%��m,�7�/���6�hQ��tF��cо�����~��{h\��������ϓW�d�}�����X>�\]�w�l�-��SH�|S�|5G�福M��w�GF8�Ly��y�y�:�v����ĥ�A�{'�Acy�n$`�A�h3Im�\�n���0��{����4�7
�/�k�Ӟ�;����{H�R>�)GƋ�W�d��М|��]�i�2*���Z�5�%�p]w,����g�o��P�V�:�Z2쵄�yd|7D�<����1(�LAq��i|���	���p8���('��ސ��J��S`�s\�!���z�w@�j��a��?����>>iL�����k3�n7F��`0��`0��p��Ч2x����%�?�`%�w���
?<~X����*|t
�B�� �/�&i\�Eo���7`/��9Ǆ3\���N�8�vѣ��D/�ٰ�A�{�+�.Q�fHd�+���\�R�Y\ꋶ���B�I'ƞ�����uzݨ��il,���N����4/�g��P�gs~Q��=�w{�� 9{ޟ����7�n��RX6�������cZv��2�������e��0(�f����5�E�B��&*��k�ٳ��BI��ݝ�����X��b(C������:1��8��G�b�\RH�tqo,�/�^T��.h�]_]�7{^v��c��e�g�0|�ǧK���0�r���ާS��W�%0�ǣ�Zwi(O����	����h�Tꝛ�_O���MS}<Q.#�ti�W�	�
�W�0﻾�����|䕛M�ގ��V����k7�n���=}�L����T��h��I>�D��$�Q=�)=5��q�'��B�mPK7�ĝ"�L�p���R�Z}��eםnu}h���Y�Ԣ��m�O�� ���QH�����,P��Wqkf|3�Ne�3Z��؋	DX��p5���+X�x�w�v��}�P�]M;g0>ͷ'� ������wwzX���ۛ@x�̾�=�7�Ol=(��ٮ0F��`0��`0��p�~�/���C0���J�}Y	�}��*�������i~��*���GUxr
�,�Xt��u�dF��*<�|����''U��?�ʋL�|D�ʱ���R]�E�)͐+�mni��Hs����d�%P��S�/&Z����3nE���������8�p�����ZD��g9��³���~v�|?�v�Og�&�^��(������uKVWM�HX`ˎ���/9=Q�����53k��]����hp-=����D04�b�[�����߶�]�HFb�m�Ƒ�U����P��Z�%s�!�|8j��Č.H�V����I+���_3�ƅ�b���ӗUx� �HV+�R�xO?�BzGw_K��⽏Z{+d���������غ���������}�y&3���:����lЈDfl�Po�k�f��fܸ�QoK�G� 4� i�������y�7��0NX�iܿ����%\�� ���tӎ�B���|�t�Z3˽!��#��Mn��8�$���
�^��ݦ��m���YT��i_Nh�	����>|D��?9�P&@Zu�����ۙBw�ō���t���fhJ�z/^Z=�~Ov��]&6<o��Wu?\������������r���E��K���ԌO�~���/����8���U8E������f�w"��w�c�Z9A-�0���0����xZ��wg�s�������u�̿�@h{���0���3��`0��`0n����-\��1z/�Lpto��
���'��ɗOaE��	h�}���]�b��샀��,�J�9K���B8�p�"��Ș(Wtӣ��e�5��>Q�JZBj�¢�2��(�M���4Jee�$K}�9]b�Bs��U���Ox���]��`$Ҟ}yg����"/ϝR���[�jx�My�o
�W.�Ѡ
c_P�i���m@�N��Aj543J$T�̖C����Ζ���[_3����7���85� ���R�,�P��L�����3K���K'����ǌF*R�����s7��鉓wےIG�-zY{�ã���yJ�4���ڣ���=s��큖���Ec���q�ᎃ]�M#ϳ��f$�i�!�L~f�IF]�̠�,�ܲ��L2!J��9���>�|��\J��@J����1�Z�ls�IeF����?.�& �vL��^Mc�:a�`���-.^��1x��z*��
zc�����/"�!&s��T�S�{5�O=)U��͛�qP�X�X����m�S��A4ߐ+�=�u�;u��͹�O+�}ܘq���Q[�j��<���4?�;S`��o��#���0I������T���"��|������G�֎}3�w��g0��`0��`0���B_H�bH�X����}K4���W��DM�5�'��>H�-Wx���2��q赐{��.\����/��� PL��Ch�y�"�̑���P�3���^֜����Z�w#���8G^�C�S(�1��K�'���t��!���zp�e�LVժ��c�1���Kb���wVI�i�
4�޽�s��?�;.�AK��{���իy�8�*�V'G�c��7�f/ۿ8�/�?���y탘�J��7��$�����|�J�c�"��Yalˊ�)�koq��)�|!/\d���#�h6{�/$1���_���EY�W/ĸ��l�X̠b�'���n�g$�Nk��'����]7F1Ƨ��Z.����箆,���ܵ��C�K�;-�/�f�ύ9y��� Ӧ/6s+gCLtԂ,�z��)B3�@��-��G�	�����K�����n�u>^�mw?�-�*�+f(�Xm���K1�4�B�xZz���Ӌ��3
�,�L��w�<���Z��!�\�i�̡�<����A<���i�|�Xd�9׵�G�U�V�e�e�L?9~�U�R!�?��?*�ϛ?k�T��g�p���u���Vmd����p��>��`�'S�~��G�yJ馛�Yc|����P�Oοi'c��x?��37c���`0��`0� �/���cB���K{9y1�%��kl*w�1�rn�>��HY�DTq̌��B���4�s,��j�����X����u>�%i�⒘t<�K2f
���o	���Y�őL8��%��4j����ƈ"1w(�b�g�QLb�wELo�r�����ӛ�A����.��X#���T*�"(�D���i2-7]m(����Վ�<��5�*��^da��޽w����^G �Ǝ�^_́�z�4���@�9��Č�(Z4��z����$u�7j��ި�-��Bwi+	ONQ������R�gCI�wD�k�=���y.��@ۑ��'(���g"�Ux�-�����#��G����Q��^N��#hw��p:�9�%K�Z^. �_3|���$��;s�	m����H���D��p}]�g��_�?�m���&��e�%3�D��b��mO[P�� �T���,����4Q�0�=�2�4o�Z�<2�l�� Z����x�zَ�x!Q�p�fv�_��.#�z(�{ƽ��@c��s㕛�����3�s!ǻ�ko�����Jq^[/�~�K/k<�k,��ӦT�rg�y��0E�7F~$��g0��`0��`0����'���v
P[��c���)+���P2 ��򬌘�u�c8H��4��q���%���j�S��gtW�^����v�:��+�J�!F�@^�a��fK�n��,%.��-fR�l-��
"��	�����֕Y�Cj�45�2}=-˵��L������[N������G����1~Q�
���{U�Fo�Kd6���ez�V��[\#p��v�b	�1��y��I�Ϟ��t\��t
���aNf��[`��?���
��z��_Т�D��+˥��+��5�݅�1�0�C��g�D�~=�8Q�R���Gs<�P&=<�����G�������.|�Z]C}<<���L���7�ыn��A���!}���%�<�Py���z�75���Ưx�͇��#���q���k�5���o譾v�R-A߉ص�moIynkE��и��tM.���R73�Z3õ�j�J�6�`%'xA��@�-�%g�>��`0��`0�����I'��N�    IEND�B`�PK
     mdZ�=;��s  �s  /   images/446f47db-f7ac-4e06-8ce0-bf970f803875.png�PNG

   IHDR   d   J   MD�  0�iCCPICC Profile  x��||eE���6�G��y�]�$�{�R�f�IvC�]�%�lv7��l��.  ]�4\�R��4������I���̝�x����/�}�Mδ3�|Ϲ�^��3��¹��I2o����)����gu�W���o]��z����-]]	~���{,i��G�i����gݙ����a1~���a����_��B��'���u��Dc���!z��G�w<9�����n��oե��w�vI2n���ŋ�d�.�4���`��Ҽ�\ ��3�͜�$�B"��K��>�Ɯ7���9I2����ó�d-���׽G�5{���69�L\Z��~���ӻ��ĮU�2֜�ff����[��?8<4�u�d%Ӵ)KӁ��X���L˅M�M=M��K��n�ٻ{�e�'+��IW��d��5��N�˒f�J���֎�5��׭���`2���P2�l�4�]�3�M�^��ɼ��gI�Ԯ��T'~{\�s	�Y�ѶA{oR,���g����u��e�C��,��@����jM$=	�Bos�8}l���-!���Ƕ3/L�����}l3%�&�ڗǶ�:IV_;Ink���6��+%�%[&�a������S�s�K�k�ے�'�W�ViؼA4�Ұw��g4\��P�k�V���>�Q��zbte����|�3c6�;��1O��t�̱W���8;�q���J�W�����/���W��ʏUX������\叫v�z�j-�ݲ�^��5�X��5�\�{k~���k}����[��u�X�����{e�C����ڠm�?o��F�lt��{n2f�k7����=��1��/&_����/�N?����b`�m�|m�k����[|��m.n�ӼCm��{_�Kzov��� �s�^z��Ӷ��������x���h�lҭ��N��N�l�s[��׏�咎�:ߚ�aW�K�/�y~��sv�f�{N���|��S���덽w8e�s�����<�O��s7�/|zx�E�.����6Xv�A�|�w�<����:��#�?ꜣ's���vܣ'�{⸓.<����O?⌉g���Y�t�%�w^��Oλ���.��+/?�ʽ~�r��k>���q�~9���o�����x�7O�y�]��s�}'>pȃxd�/|��O6=}�3>���S_������.�m�Ƥ�v|[����}������bE�W��h��(�v%&6�6\7j�Q��zc�L��^c^{�u�ݸҬ���/�|s�U�]���[��5N[�µ�^��u\��뽶�����č��x�M�lz�f?����ˍɗ�0�ib�ӷ��ղ����Y�\�ts�ǿ�B�f�o��j=����6n��W���~��w��k[�tj�E��k�s�Ǧ���;_��&�sש��u���v��;~��3v�m��G���=��G��ʷV����V���=u�o���E�����9��p���z������7~2�ʢ�7-�n�.��y�вesЙ_򝛾{�!����Q=R5�{�=�%�������?a��:�ړ~q�\u��]z�O��3�=�̳N=�?:��#�=�����%?^�����h���t��Y��v�˶�|�+��������磯�\�ε�]��/��-7tܸ�M���yѯ��[O����/���_��7w���;����w�q���|p��{���x���=��C�=|�n}��G��叝���8�O�=�詽�����gv�v��6���ϯ�¸G�4��[��^]���4������xs�['���|�w?����o�����}t��ϭ�������5�0j�QG�zg����������m:��f�?W��r�*��z�jǯ~��y�Z7�}�:����zoa��m��F;n��&�mz�f�l~G��/���q6�شŎ[N�j��~��mNn�q��k�|�����9�*[�[5��*v�m�����m��ܡeǩ_�v˂I���<��m����)���|�;�T:���թ��v���e�w��4}̌��M�}�=��o\��_�O�~c�����͜1�?kh��9G�����^?��yO�}a��Û/b�ۖ�t��pܲs���~�;���CW>l���mG�vԜ���Qǜr�y߿��k��儻�ȉO����ϟ�ҩ�����o���3�=��?��}x��~pއ�t��?^q!�xqr�'?}o��.�å7\v��'\q䕇]u�ώ��)W�uͅ�^y������nx��'oz��/���_�}��5�^�c�_o��-�ݹ��������̾w�}s��灹�~���y��?��	����S;��S�8�O�򐧖<=�������.���\�����~a������}������m�^�����ז����K޼�k�y3���w����Z��ZN�����㙟��H~���0�ἆ�G�5���j��c��d���4n�qo�t��+o��߭r��v��g�q����u�ڷ�s��O����W@���ԍnrڦ7m�Lu��l��K�&>��-n��^���m�mڦyRm�������������y��m�w���:;L�Q��e椃[O�|Yۯw�Ӕ���~}�]L�n�˦�h�-]�u���;y���#v�h����ܞ+���䷧������3��b���>1���/�ys�}W�����;,�Zؿ�~Ç-:m��%�\z��>�����>x�w�w�~HߡK;��K����Ǐz��c�=v���q-�w���N�wҒ�:��S�sڡ��ã�8��c�:��ct�9'�{�yg��?��U?����/���?�����K{��.?���<��~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW��U�Y��U�w������s����`����������cW?~����'�{괧�������ß=���z��G��������ۥ�\���{��7�zs˷��g����s軧���_7��������[��W 9,��Y^��$����]�bŎo'�Ӯ<��wW�x}��a��r�I�����I2�KI"�a��g�lq:0Ǫ9.͹�g�G��1���)Ã����&��8p�C'�]2���Z�ޕv�[�$#��j��::��&��F�$�޽�{_3�m��u�:�����W���u/�� ���};0{�^o����+r�����)E�=�?�Ư�8>=����z&^�3�"����F�6�������п?Ϳ�~��W�zF?�W�3&w�o+��9�v2� ���z��3��i/VJ����e�hq�>�[�P�"p,HH%8�����/����\�� �����p�e
�Ҝ.p�j�����n]	��%��o��?I怚���W[25iǘ���|�}��n����&��[S�p,B�2�:�L8�=Ȁ�Au��z�c&8���!O��e���7�} �s�;�5-�:��g��?�?�2�\�M#V���+i��A��"N��pmS@w���$%31����Bf$#:W������S�7i�D�� ����?�!� s?�4�@;��J�:�-��SX����e��|�I|�?o:��0� $�)sd���2���K�E�gC�vs������l�g��A�s�"��m��j�R��������;����2<{�ܹ����C{�/Z0���?<{pqu`N������Y������i��Sڧ���:sh���������޶��ƞ�����eUf���V�m%sՁFL=�����������8�����e��JO��)m}��;�zzۺ�'��uv�M�nۣh� ��;z��;�u�u�uU��L�n���tOi��k����=��mjo�q���Ńա�:K�ۿ�kxAS�u��ÝK��;���|]}�{t�aܝ��zv�6N����Lj�i�k�~��J�(�[OW[kowKGޭcz'�6;���Z'w�j�5�eƤUkk�k��j��Z��e��2uZwgKG��m��z���ї�i�q����ʌ��m��:�����aRwKo���}]�zz�'u�y�ʤ6�TİGGGD��=m'z�Si^Zm�oN�����܊.���D�ڊ�\<8�����9A"���k�fk��?f5?��Ξ*�e5�Xm��a�������K�L����=���Y���H�C��:ZZw��!?:���=nW~3��sw7d���������8��I��3��z �jc3���sڴޝG0u������Ӷ��6K�qZWo{'���	c��iS�4�T�2uz礶�>ld�����=U�E<����o':��JOKgW�S
��n�����I������������#��i��fZ����A?�c��V�2���'[�F�
+a�ҽ�U�jt�W���^U�ƅIU�����~�������8���R-2�YiҊ�����~�f��k�q����O�����2��~�	f��ʚf�[�O0�
Q1Qz��8(���8:���'%�JM��=����&2�9�Ei)h�V)�T���c�e�k<�R��<2Z�Hוl�����AGͳ*�]��(4�M%�2����*�)�s]iMs�Y4�q����u�r+5�`�Iiy5n�E�م�Y-�)�@g�٪�%�#�%�_������Ό��Ԡ<F�J�J��X�05e��T�B�)����U%�%�1rנ�*Nf$3T/�i%C8ľS�v�Y��̬#�J�F�-6bY�܎>K�MX�6�1�HJ�H�U��&�2l�p�4[��M-5�$*���NA�� �Ժ#��e�F���ƪ�fRn����I�2G.�R�H��
<P�C�G%�Lf��5!�$��j�x�י��5��56��@���0�)l�8�z�k��~��R�Sk+p
��Q�:��Ƥ�ր�{� ��)�T�[��^G0��$��e�TY�#f��p0ZV��dXOp�T�9��@H7�R)�F+s�u���I)@�����r�
$�tMH:�z��mKx��ž�K@�p�D�G�%���ʩ�%]C��T�
ǲ�Gs�Q6+SN�����~*���L���p�8w�9iwRA#�5f��	%�AX���K�uRKK�uk3if=�Fa���K��*\U��y��#2���"�'����&�q4�xMl�i���'~D�T���@+G�$ͬ'������ ���B�%�ZU8|,ܣ%ͬ'�/����;�m��>�"���N���a�dA�t����,U�YUX�ι�:�^��#��0�	`��FA�֕�0�j�:~(+L	��CU�q	Q��u�Dq,����p���?CGQ�h������?�>�����=PH�?C�_�?�*L���ʩE��;�:��*J���+58��Iޖ��	�LC�d/n6�FC��� \��_1�?�$U��N)"�(�4����@���#&��I]�)U�6�2�)p
P{سդ�������z��� ��
�C����{*qR�JM1�T�� �42�U�hB�TJ*t��b5,���h;0�\��Z�F���*p�Z�!�:�t�jx		,��a�`�FT`)��| �#$9bFhf���Q�ë�R��%ͬ'$ia9Eq˒$�TFp\W��a�_G�,Q��$�#�Ru怈�HS5�@)���76�R�Zҹ 2�,�R:J����4��pE���$"��(���p�_G���r��>��P����j�PX��zB�n�w��0#�8y���(�؎$�'�0��C
cB�"�R�iA3R�z�0	�o� $CZ�f̠�p�v�u�!p}�5�#݃[� �Z(|���	x�a�����G��j ,*J�d1����%!�B,a9�8�]E钬!Be��'&���2� h�LI�gD`E��Q����.8 9�([����
�Ԡ�O"e*O%� ��d:EG��e:PFX�i�s�a
���X!�F$�.}0�P�9e,��c}G�U!(kd�FƁ�C&������ܭ�#�i��)�%�j���QĎ��8 ��A�=9X�/ WS���wD<Eg9X�?	��=�ȭ�;

� ,���{���P �K��x�@*�@� Dq��<+֋l�>Y�R�g�C���	r�W �b���A`��SN���D૘+��()���@�vd)*�������� ��)���BN<YuT�Рd�Ry��Dq�jd8��)2��(J9��*3*�0#I�p�BW�,�(���)�T�j2�3G�tQ ��W��(�G,U��bV!����?C �A"�/�-wE�k�b��d�qF p�d�>0� 5����%�*V(��F�RR�wK�;�O��g� "wnX4�T��R��1+���[0��+#sQ��+p���W�@(�"ׁsd��Y�G&+��x�(@ #C^N³!X��
�W��3"��yXE�3tP��U��)����������TE���U%�R)�g�	�����
�е��=�T ,�ܣL��(��q��5 aԹGC�F���pl�{,:
�r�F�s:P�I�-�J������Pmi8a8��Sa���f%=�bIU��gR���TH�>����mZ�6��"���'��DO^�[���"�g�[����� ��(q�Q�3
v�%��(��:��eU�b`���� 	E>��C��YVG.z"�d 䒪3���u�3����w�(���Ѯ~(]-����YVK.zr��T�#+�����jmy�񫥴�CH)ὔs͚`z%+-'�@��`(�%���%�	;��e��ؓ���M�@�=m��=Y�(4�� �1�p�䝡�����KL$J�����մ(u^2@��)�T���2r`K���fN�3.d;��\�I:~$=��@�{�~��*�5z��t�S�V��9�jڧ.q�q���s��"�	U6��eSY���}�eS��)�f�)0�iKzFϔR�I �`��J�+S���@ rZ6�D�ŠU~8��L#��� -���/!o�ی��-[Pi�ϴq��2�Ig��D\���j�yY��y ���%=#A���i��Ǩ"CePڧ,�q�������T3��%
�SOU�5�& ����kAu*�Жt���U���dÆd��	dwH�H��Z=�Z�QIy*�Q0�&+���%^3���q�yBR��w*qpNz�KӘ��`S���K2��Pt��A�����OQ�_S�q�z�(iNV�M�$&H	��1
WlDO	� ��L�Qqr�Ty
��H���cJ��D�7��(�J�¸K�0�0�
=Ed�?'���4��\������`t�L%(9�qZ˭��P�3���� �!����U�'�g��g��=�}�f�P���L�H�EO[�f�����J�r���0�(sy�@���Y�t<�aj�9EV�

M��)���r=YfiNF�G�A�c��KI���I����U�HV��q�Tw�u�J'WyOn4��(K�cOzPĀ%H��H�)a��\�,���B֨W��j��J
o���Y���+�g�łzl��i�S�`���p�����e��}Ҝ��g�'��	�h
���.
�V�;r�p�6��fȊ���,3��	�
���~��C����2+�QT��/zR%�S>'Ҹ~H�����V ��* ����J	�J^�o�O���(��;�×t�R��ۢ'E�T@[2*S�(�I�"�0���#f�̸���P>MZ=DOU�3n�����:=Z�甔��2?�Isfy��V���<�8z�{R�R����K�?�ׄ��ZP}Or 1:F��q�TR��cq����A*0��W�e`��SGeR5��%�z䚹�^=�.iĞP�Y�F��SN�9�O�}~ڛ }̃7K]D�H}��J���(!��P�	 ń�"]D"l�dIt��Đg�(Rq�Q\d�V�ʒ�BfX[
���1����)\�t�����vȅQ.H�o�,�Ӕ��� ���'J�����)[�
MȨX.�#(�ڼgF�L�9�x��=�|�t=��BBz�������&�bR���a��F��q��PyM
�i��!�	I��F����pʤ���<O=	�iQr�q�����N(���)�)���Y&�
27�dqѮB7?�����C���
۳����ڭ�O�[��Mb�rÕMVm�o^�y��Ӽ��c�y6�u�yVF���mD�̪��]6���EP� ���!������&z�Dw�4E�j���9-��`�o��yCs��1��%s�-j�6��=�r�VYrIR�\�����$��uH����!��-�G:^�g\DR���ݓWJ:^M7��+i�Ƚ礥��@�x���8�Z�*����ע��b6�K��缔���$2c�tňx��G{�UѩOZ�	��2�-����Ll�HCT�=�����jEh1:��N�|T��2�EhE`t��������9�@��9^ZB��rFO�s[�/�uG��J@�@��Μ��;��?1��N=���%u��RbǫSzt�Zm�]x+��At����n��A� �����,�W�7;���D�I��'qX��E��}+��n
�:W#�V�zU~��x��|H�HԎ�~rAѵM/�@��٬���Đo�n�1�I�9?��x^�$�Z�6�df�r��B�疛�k�I�
z��0������9�L�d<�D��Gb�\�	"o58='��|7�e���,#_$] �����ߦ�3"�d�9��7$��V�$�~�5Г%��*52�Y�u�6�p����,_B� ���U�nЄn��x�Q䭈�~��":Jߍ*z9�SIתa�<�$��|~!��f�i�Pf<)����s��]�kuY�$N%t�����Bb�0y�I-�9�)�r^�?^�V���Ҧ*��X.3�^��`��ZA�����r�_�s��z�Z��yu~������a�s]�ru��_A�xA7a�v�㕩7H�D~�#'�)4]��ym�g��iH�Ck��Y�n2o��o��S(RɜW��H|84�TOB�r��(Z�V#�
$g~�ty]z^�_�r��MV� 	�)��&�F�DM�9'�nN�y�5�\!�N�<
��<	��K* 3HV&��|Λ�f�ji	��6���r�Z%z�@ʠ%�J���7����I
���`o�\+�_�� �K����V1(�w��/�$�c��"ZAx�J2+F��+ϋ�٠.ጵ��S9�k=/9k�j�)�u� (�t�d^��N&2?B�+���
}��a��;F:Mu���v�c�tN�:��PQ&���E� �˱��@������q/�\x���>P+saϓ�z�D��܏�è�U3��PH��IN�]�[\�g��=L��K�)q��0�g�,�"��|	�X�j��_I����\�X�\+�i�z�5{O 2�^�"��­	�2V��~��� �e�_:�˯��7�y�,d�ݵ��D��e�C���r�*@�6tC����C9�*0DAfE�������'����ޠ�{2]|��I�HH��
�L���{��/�� p Y�ܤ�j�N!�d�y��t��n2��0L���u [ɘ�![|΂yO����������0Z"���D��x��0�W��đ����0p�և[�ڛ4'o�<bfl���OhE��yC�@��Z�'��1�GC�8
��{.FW��-0�7�HN�7��Uy_�#��Ⱦ�C:������EuӬ yȬ8��a8D�'��&�V�}��d�0}7�9��1�#	���p~ǰ�=o�a�՟0���1CF��/���{�2{�~܈ahZ�Ρ�2�Z��1��7&�T|���6�WO��er�Y<���_ʲ0��>BrJB��"��xx���ӄ���[`(��a
S!i���+)��H�׳�a���%G���$6ă�D�)Y�D��8A�q#��p�ޭ�L�ԑ���[`��F�{؁��WD�i$�QyI�g�y��g>nR&�]7�����Na96+��n=o�0X:��v�]<� 恷�0Xm�r��y3�yC��T�%|�IY�1t�� �t�6�,b��=�a��>��F�\[�#$��I��ﱧ�BR�UP���h���-0��2��T��c1��[r�S�1kU1�i��R��I���1}އ$��U�5���ɽS �¹�"�z#����,���eIoC"b����Z:pR���E#$���J��] x�*"��y=�T������[`,'�E�	gA7e3�[`,�ER#汧�F�'D �O�;�֟E�0��4��U����ED�� w�n\i)�-0]m�NL�B��)��F��X��_*��AF#�_xCY�&z��-0�>�f�e����GɈa����̼��TH��AF��2���T�j_ޗȈa$2'�}���|��g2b$����&�t����0HWT*�$���1��a\��x�g�"#������0U���x��H�UэPYNbX��2b�n�R�Rg���0�"������K
�y�)�O�%9J����YDC�\�NC7�9D#	q�@j���F��
�xT��XЇ�a��yX$\E8!����1"w�- m�:�ce1��Oɛ@Zx�9��FRu1LL���I�fàՆq�����~܈a�¸D���G����d�0hաbZ�:ݤ�k��R�nP�2�𵷋�a0��A Ï(�㐊FR���`��i�3�[`��S���5ؼJ�x����JB��`��U�0��/sOʀ�1�J��-0ZC�H���С�i=o�a��m`���%�>��������-�'��W�u(�[`�����w�i�k
*bŘ�ABk��MK_�P�(�Wo�
*�}*=��511}ZW�����*b�L�+�����n��T�0���+}���	0��uZ1�E�U�;���>`�y�(�{�!z݁��>�Q�(�[�ިXx����1���?�ʐK��k�y�`AA� |�Qt���Y�0��3�a�*t=bEwȳ� |ȧ:��Q�F�9}(�=F�1�k}~���xo�ȭx�F�3�!X��Ǫ�a�e!��A�@�P�V� �����҆ڕ��ޗ�A�p��V|mEG�+}D媠}p+��a���ح�礦˙��FY�@א��R��ۦ���D�=�?71��k�{���)�C�atV$m��R+��:b
�,�&�&���ǩ:bڭwx��T���WG�黩�s�9i����a�d�^B^�C�<>��h�SAPT��"���k�x���`��l��?�À�{��X�Ky݉F#��O�#���5D�"|2K�T 9=�p��`
�Y<��O�Hn�`
��%@g��@執�a0��nE+���Iz^��FCS���B�J��a�
5��M~M��sވa0E𓚤Zu�Y:bLa}�Hw��,��5DC_�ࡄ�¹�}~�#�q�گ�(N����y7T3<���lz�c"���)'?�:���8d"�A�

Co�2C�R¸�Ak�{����5�bW�G��5T$	�E]��-�뺉�Z�Ã��89o�a���!�׀��͛�a�5���-OZ���Z=ޡ'����%��1�� a�n����/��a{5�C��X@Z_G4��W���W0o"���~oàU�:�!�/H�k�&bËg�=4T������pև(�:i"�!��^ʇ�� �L�0`Pa�z� ^7à5�>�X�¸:�L�0��Z�;��ri��Ɛ����4�<7À�P�pB*?,�[`����-��GHz��kL&b��3���6X<��g&b�{Á��C��x�D�PP!'�q5�k�&b0dv�CӰc��#�1�e� ��]<\��+11��Z!���b#o�a� ���z�J2��[`C�)�Y��z��o�0�M�c f�&�k��+ۈa,}Q^�fC}�����1P�!��.Z��f=o�a�V�<�����]�����{Ɲ3�!7����E1��a�p��`0�c�����Bɹ��l�0"!B
̛��/����0����o����(��2�����xa	��q��_o�0��*�W�����<o�a,U�Āj^�ع�b#���)��R�y%���җn�7@��Oڈa0��
2@*��5R1��uK��wA��<o�a�G%����K�d��-b�3��ᰃ�4�x�-0����n:⃔<&���%�;pt�͇qrPao�XCߐ�I�t֕�r��Xz�x���[��Iϲ��w�Z,]��֥��Rw�$�XRP�Ȟ�   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �    �  ��    x       ASCII   Screenshot7�o  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>946</exif:PixelYDimension>
         <exif:PixelXDimension>1274</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
�g.  @_IDATx�}�W�d�u&�]��Vey��NO���1p$8 (�� �B�Jz�V!)B+E�e!=*b_V��c#6�z���$  �8`L��������MVz��w�of�4V�SSUY�y�{�w�c��܀���h{m~g���?�'��C,�c��o|>��}}^ܶ���������w����^x�t���B<�������[���s�0Y��
�����o}��X�9x����k�>����!���ue���7�5]dc)8�*��}O�⇫�����>���'�G�ɕ�u�8v���G�#��D2�F������!�Lb}k��]�t�UO��T\#+���l��<∌�'��ӟz<�p�o�6ޫ�E�P���&w�eT�*lG��l<�:�z�E�tTP�d	1
��j��7ηuLL��i�p��{X���L.���=��Q��^��mܾAL�P�6����C��F�����A@Ax��q
'�j��u�)|[<�ʡ=�!i;H�1�_��4��6\~�����o%%�4z~^��GW`gS37Q�v7��7�La���{o�SwP&��?���$�?�"V{h�}$b4���G9vI>&���G��?P���(p����)�c��c3b2#��im��A�-���<�=���������m|Ը��������_ާBxa�Y�Uk���9,L�Q!����q����^xS��Q�"����<d�f���v�7f�sZvA����q��ϥ�����`QеnW��A���^�Bs�~��k�WY�f���Y��X�ΣK#����ФR��>�c�K/��=$'m4�������}t�����Ǹ��Vh��-��-z},.�"p-<�X�ks�h 	���U�{-�4�P�T<��N^U}�	l��.�dn	i*�I���Xŝ�+��_�3��,��Z��c�y,�)|���v����)�%|������7w��iu��
��Q�
%MZ�O���D!^�F��y"\�����]�j�*V�â�Y��^����'h�%|�����]4�]���.=�CH2R�,6�\KN:a��������'�y��7ϷG�
��|$	���Դ��v�%}�[U�UL�3�F~�%��u��zx,N��]�Q½� V�I��{Ԛ-d�	���*�:j.�_�O�C���=p�4@B<��>u��I�{|��r��'�/���û��8iM�2
q��xf?���`!�U��}��x�W�����<ї7߮v�Q8���_>��:�����nuM-��<�r	's(䒄��żZ�E�&�i���87���4�o��U{Ml�v�Xi���"����>���4Ob�M8l�s$�X�PQ�n�T��%L�Vۻ����3����v�B�a���l�G�k�X���o��|��|��1b+M��x��+��&~��W��x�>>��`'�X=���Nfd��%r�����\j�23���u��ZDa�4?��_��=�������46��:W�x�SA��0��W�:0Ӆ��*R��$1գu��D�V��*�F����h��| G��(N��q��|����%�a�Mf\�ѭ�no���#H���)��}����u�bxs���֖p�4�]�D�[���l�Ԥ�">p5����ė~��϶��^�>a��h���=f�/eP���g��q��`�Tx���f��+�q�Ә���`�9�w�mSy�Ӏ1,��xK`��qm��@c�x����*�8�ps�Y���^B堁�����2n24�z��P����M'#:5$�D
J���@/j�xA����%��+,�a��i׵v�Ytz�l���ԙyB���Q��z�=>�F���d)zL�śH�b Ϧs|<�1D��B!����j�6㏐�  ��;%��[1�*۩w�<4�M�<(��\,�{X�q��^�B���⍵Z�MGN/#Up1;}i����@�O�A�7�|�����T\��HY�|�K�&�Q.�~(_���������R"�-�������F�^@67AK�!E���&a ��+l�� c%�B�ZiRX�%.s��c���I�~�2�Db<{������a������G���������oQ��p�����F����ACH�3�_B0�Q$�^>���ߣ\? ��^P?��	���-Ɵ6�'Jo�ڽx_Ԥ��kwq47�����&�E�'ۊ���.ag��������_�3����du�~��w=Y"6A�K�����A�;�ޣ�Vj��㧒c�j�4^����6��‬/GF1�F�����}�W��p��9���w�WO���ZUy�K#��G+���Z�����C���&rd*m�T�T�0�z^�:���M_\�D!����wn�G�a����;��;?��ӧ��?�C�P�k���G�˿���/���i�.��������o�.]��D2�b,��pЫ��.2R�A.�A��@HŒ��1����Iƒ�ē_���S'0�榲T\;��$�Z����Y{q��>�� ���k��D˧����ZB_��^9q'r3J���;ॢ�#����'��铤��k5�;��ԥ��K���[��J�dE��ܻ��f��. M��{�j<�[ױ7��-	M��b��"�:����>z�K$w�%	d������_�
.�x���@٥��3Id�p^��^�h2�1�u:m�<ݚL�̀���y����A��xy��`��b<2�@�j?0�!��%�OP�\{�l��G �?J��XGy��c�gq��Q�_���9_��3H��˟�:xxe�Z@O}k[(d��#����_��9� LV���d����.~g�V��!4�;KS%�d��ʘ%�I����2���vw�F�!�-��o���]��|J�!	T.���Sӭ)^<�˷p�� ���ng���B,�P�����zl�I!+.b�Uׅx�y��|S�9�u���8��T���GYP��ĵ5�",����6���ːxc����6��]'_|W7o�|������&�]8I��l�m��H}{�eS��7o��bp#�$g_���Fsd�ro�F��tVi�%:�Սq�@��'�¿|�&��f���I�^i�j��MZ%2���)?��ν��Z�����iy3Q�`�'Y.���b�����]����\\d�y���$��I�H�2�}21╍�0����s�4�c�9��B&GV�1���-�x�8�\k���řܲ�V�uQ�on^+@\�>n�|$�����
��&T� ��6���0'������I�:��1f�d�$��[\g�H��Ĺ�0Ո���+�!;�o�Fc��I�R�+�$%R|TB�+��cr��S�� �CK�!���ƛ�f�$�%�^��3�Z�X#10Ƥ'�MRI�v�7RmW��.o`���+��գؘ��1���z��ܴXs~:��lT�u�E�pHFE�� ݋�IA�B2lE��+�;z˖��@YM�
	JE!�� ��Յ��	B+�2�U����������[�N�A>����O7�
Aph��W�-�49����|�FQ���sM�4Pi�^e��54Dp��Yq�|��V�Q����X�f��N�n�b�t�f�˙��:�2,�Yo"�J�{�P�@��H���6����3�*j�J�\�^����3�O��O���<-N��4��b o3��M�0�1�@N�h�"\Z�ͬ܎���XH[BC�h�®��@�Ē�����G����b��|�<Wr&Ɓ��$vo#�89�4Gف��u���zs��0��uY��pR�C���8��-��8T�5<̊�<�D��(�&J��F$�xr��U���X�d �q)�u��0*j21��WE��avb��WUe��Q9I,,-a�4�ϕU'�Q"͌�Z^}��c'N�gT����@��Ҍf�"�q��B'�
���"o`z-q�Y>�G`N>��'y	s�?s��if���m���?)2ڟX:������4fK3(��#�\���Ɩxv�E�ɴM�J3H�x_�n�|����%�e���0�a��3't �!R{�B\6���������l�M)�F�d!5yB&�����kJ���}���"�`�]�����`3��V�D��Z*ļZ_K�iH^9���
��z�J�٤�M�%��k�ۡc�1��@���%h^w�vM�yK��c7�w%���dJ�@+�B���
y,PB��m2´���4io�t:�D�F�9|��&��$���qE�D,N㑌���0�_[�\]���SS�8,&�0�H����M�[n`R}.L�n�V���F������"��V�Uy��������C��u�G�`"U��{��)�L�t�̇�3x%D�N�$v�x��t�������烃�\��B�O��L�v�.��a)G�����ʴ���$5�(ӓZ
�2���K�6}�_�'X�2�~�B���ҙ82�n��"�11���C82
�ds�3GK1���]d�Q�6���e�Ba-�"۵�<z/Re��Hz&�,�E�C��yq,�*�vIaӤ|���
Lz	m���i[ۛ8�>	�顗hc���<�Q!�D��]��@�z�X���f|Ɯ��	H�#M��y����R#bC¯�zR!"ۂ��e�K��-3su�.���5��//Q!T>/���q'��k �af�}�q�F)hL������HEI^3cT�����'�9�b ����(2v����5Z�1��K�H�$T�6��(h8�J����2k���b:lG)H���~z"k��&
k�&�9�萇�6uZy��Çw�`�H�mf�́V9i_h2^$��(�I�}��=�㣄�~v��1<�� :Y\�9���>_�hk��$�3�����d�P�����8�'�Z�c��A������㏑?2��?ff��U��@PA��b���+2�L*8�ص��B%S�dJ��s$�vJ-�|(�������d�#�������L�M�5&4_�j0�*J<S�l��EQ��M���!r���b��K,�R�`�<q����ÑL		Z�������X>{�w� ����e@�&E���"-m����E��rbas�%<�^���<�I��J����V�q�p1����0�\�w���{������6�����o�*X����]���G���������3--c�JzK�����P!뫐�w�LE�;�͑�[&��S�q���}���1^��d:�,�����o��;8}r�P����5�*����eX�� oZ�.��Q.ò��>�>W����\G�6�?Mz+�q��@=��W�}�Aw��*���>�������"f�q&vFc@�V%�Cܻϯ1.��mkI<9�;'��$�e5����k����`zI��%�Bn]XSs��7��.l<K��ˋ�����xa�\�9���� ���7�!S*efqz�b�����!���}��i�t~1�C�����la�17��=?h�pn(�#�u�z�s�*�0��F�^6W���ʚ�>R�(Â���R
�B٥��1y�^����:���k�Pˠq���M$�Smr�k�M������=<٭�`���t�;ث���\�U/�D�3�iQ�!M�5��ui5.ȯcXw��h�^?y�(�2x�hvh0-����Q�1	��圫kP�h�=��-L+�'>��T�^K�$��\W��;� �sg��ٹ�k:�tQ�٢⤚�p�C�#�[b\���S�/��n���!̥����^cG�G�f@�P]3���Hs�������]��� 
9����%���qS$�ܰ�1{���<��N�zx�]���[�.�#<�ɸ�(ӣ$�91I�|�x��&P1����aP뛲�HE�!��~?P"���˂���v[�xQ�1�*KKSJ,�0F3�:�Tp{�R1x-4�^C6�0�Č�H
��a� !=Q=#F�,e�Y*j�'�!<��z��j��aỉ;Z�`ZG��6's<��q�
T��1�8),���<|�ڊ����bvf��.vW��Ǚ4�\V�I�`��N�mj�\�R�ٍ�6�`� K|}b�DEm���3���EE�.ֶ��h�p��-�i��2�5# ORӽ�
&�*��C�q\���ZSӉ��ް�eFpQT�K+crT"�o�`u�I��Fk�U��C^ݣ�̜��K�>����O�I�i�z_>K���TY|��T���D����ɺ嚉=B9�B�dR-.�z��J����4RL���B{�&�w��P���Ɠu��mL���9��WI�]��?����A�Y��I,���*���#����H��`�C�4�Iq���4�i�<�Ԡ����v��-�(4����Z-��"�v����LX�&> T�<O'_Ua:*|�}���a�V�.�z�耂��]
���FhG��B#�bF�Ol�uZ�uL:jls'��hA�q̢�=C�MǊ�oۄ:�n�"<�i���^��䯄~n�fW[�R��H����q��\���>��?��An�7ص�fHݬl���2�L��7�ʦMZ��&�pWjT�daS�
�)�B���(��Z�t��[},,,h.��'�#�R-��X_�Ќ{̴1����|Z�������B6��z�%~v:Ml�<���C�r�9�uuI�Wk����6��s�E�?�w�y��H�\��2fffAD��]�pے�ŧI�p���!_�TN#����p�f�B�2��<ʕ�N�u�5���ϜD�U�5�;�6�3YU��aâ��GE%�i����`���LȘ�w��Iz])m3LQ��%E6gESeD�>V��d��S��,)+�S��qh
���mp����*���ߤwvq��9�g�0�u:=�$;�F)���Y*co���cg�/���;��	V�o��k���g�������&lϕ@{����n�`M��bvq�PՅ��5hE�S����
�Lu��laS8%*1A�������9��j�#\G���r��@멵�htdK-e52,�%D6�,�1�mni9čŴg!�"4Q��F� �H��	S����y<�$�������F��҂��<A"e��Q�yn�]�^[Z���i����˸4�@�I�����?�������L���j�93�!�rR7�e\̽0�^���nSN=D?���&1"�� �t�6^��+�<�����8i�jy�q�6�,�1�O�8�Bid�F�Z�lw�F�2�A�*	�Đ�/IB\]��	J?#X	.$D:�R����(j<�^QcB8�ǚ�2��)& �'K>"-���&inWe���'� ɽ��i�1��\��_���TT_{��15y��?�����c�?IG����Bv͠\�8o;L��B�HI)���)k[�h�R�y�ˢeb��C���^u���c�է�v50�D��f��W2�fÂ���1���Q&Ŭ��w��V*u��G)!C� ?�|=3��TF��Z3#��V�^4�)�&���dT�Á��ɦ�����s�+����o��@��b�fUɌ�8�F��뿂�I"1;���6�����.����U�����Ft�D��R�lml"a3+-�HO扅�
�e�������{^�2�깴ĸY�2$�ގ��e^�kM�Đ@!#j�8a=�ěb��E{�Q�;[�cp5� p���g(�|>��K�y'����j�u�"ƭ_�c��@�I���aK(�<yL*��\���C����%B�&*P�4}>��k�x�yl��0x�q�
S��Ͻ���v��x:	?4R�hW\�Z���ﾇ�_�]�=���y���/�FV�ŕ���H�E��
Sڽ2ǚHkkmd����m�D�Z0�d�z�UF8
�x����N8� �K��܁�I�K<W�O$4>���Z��X,�G�;��L�Ɗ��X��h���Dϋ{�as���A�	�C3)�L!$�^3Y_���q�����˳3��_Ǒţ�W��s�����3�6� ��Wr��~v�cHǳ��`5�������tǢŘ����.:�rt�t1��a[1�2�軄��-#��m��:��Z�0�>aΣ�ų	���pBC� 51�uv|�7���5�����Q��I��L�$�H0w]G�J&+dB�����	!RE{F���=���y���0s�n���?wϾpQ��u�����*�P�UPJ�"?�\#�?~����t�|�G�Eq9��/���S �ଆ���b�rɼb�%S}��h�F>n�Fp+��`��>�����7�"�+0�_\8���oj� BpRn(K[��a�&��k?�2S&L����%EL��U�A8���'8ҟ����p����oP�!E�:��D�x�T�f{�����q�D	;Ovq��o��^��`"TW�=�Z����b����gZpo����ۿ��Xi���u-�Ǒ4p�W�c*���ͧ�%S9�d�B'�Y@��M�?�l{r.�l�����S�8�T�4=�5�!���5��O;��sF��C�S4=�+$�dE�E�۸�����z�PXgB��I�����(1BEew��2�ѨƿZ�4�p��E���:F�Eoh�e��z���h��!A��hѸ��c~�cin;�
�./��&���e��6�	Y��ZS�w[85�ڃ�^NG�\�yRƜ�ɏX��d��P�aj~�F]-Q��;ثul��>]:�vC�0�� �nQ��9J��(LH��
�4;�J���PY�^���i��p����(��֡�Ŷ�;�q�3��DA]<�d0���n��S����Y0����^��u4�5�s�9�,ˀ�&�f��^8������P�.đ=���q�'�96�٣���It%�oHcK��)�4�K��u<���T�-�)�nZ\�}#�$R^�h�R:|�Z���:w�REB�
)���6'da�y\�v�Z=7>��F��a��y\8b�a�R�K�u��">=�M�6��0n0��/�~��&��$	� `��׵>/P�#�#�Ne�]暚V�P�R
K���&{��^��Z��~a�_�	���]�@�6	� ����0���f,O��)k6�t��CƿF���4TEA_��	��)�z�V0*`j��%LI'z����!�Q�\J'���E�-����l8�!B�i1t���Z����2���͌�ny �O2���R�t]7�A#SK�������2��Z��*^KQ/��*o����C�x�=*�D����!�*��+3�Ӈ�2��*��a:�s
$ 2[6=����6��o"!B&"e�%��^W���HVI��x�*&SH1c/��Ê� Wh�29(Z�I�:VXV����[]�3�6�}�L�z	t�-�1�:9�?��������z�J��IY'�Ǉ�I����8	v�2��"/W��W�>����=�V�*�|���5X/�e������|��7��8��3������,�4^"r�`�Y���ѯ��+���h1q�"�~�F�D�̭��b�ޥp�dfIdb�m����#�Ǳ�:����g5�&�0�&E�=�~�Զ���w�b�����lX,6�쐙�X*�6cE�����G����G�G�q/8T�W\��轌� ��iO���
/���\���@�����;ؼ[A���3'.�l��?�ɹ~�'O#U��CdkAc}��?��Vh�����l+�D��1�׏����Cڙ�7���W��}׳�Y]���b9�@�	3d�Vօ4��� �`�=�i�v�`�1�k{�(ʸ�(�|ԧ��m���p~���:�����x�+��|w��bg��Cp�h���[(�%�,`�^��&:RaN;�鎳��mlbj�2f2G�5d�N*�q��"�H�	��}:��4隌���]�BIQ�2A�Ig�)ft?�X�$5��U;lW��mvp��w��ų�����Rpt�S�%x���-jv[�6 ����r�=L��1sae�t#Bd�6�)��8��CY�~�"��?��qp(���~Ȋ��B
7~u�
�8����-i�m�����\~�>X�~����!j��c��;�x
7�װ�x{�Q�.ȝ����Y�ʓU���R��V� ��mt�����r��i;2�i�Pz�;ڴ�V��խ�Op,W��_y.����g��yĪ��j���Mgp��)|r��|x��_dBi��'����n(��F�A�������O{F�J��?����-�	��t:i��3TC0�r���Ej4�$��6	zx2�G�	e*�ѱV!F����ʛ]��Y���S�q��U��G|���Y`�y�,����X>3�,J:}�����x���]�����˧�����z��7����0�'�x\7Ô�et�=���<����;�­2	��땇�:�`=E��� l�V�S���=/�:�#?GJ)�W)���
G2�1N<������~Af�Ssh�~Wnczf6ߴYoaaq�o�8�A>?�S2�&���,
�P߮��0��:Z�u�(���p�*CNZ��3	���gN�n:�)ۀc�xh�N�k��3�TQ4_�������`[��ŗ_~���ã�+�.AM+�9�,.D��M��~����p*e���0Y������71C���Nz������˙-�.�ΖP:x�p"�V����I���6N���$��jL.��"�\,�`�Ԥ.��k�4"JQء@̉:�$5'���C>���ܺ��k��rj]Yҿ���8��å0��wr��LJ�Eh�{e�����xu����)��nc��`'�1V�<���ǟJCh�0�(y�X��#W�!7�Bi!G���f$7���-j�`���Un7�����kz:�����]�k_��s��#n�F'����B)=�fǥr�%����Es�a��L�9�%�l�Eq]�1�Bo�]�}7o��W��e�ʍj_�o���[�3�*٭`����)����M�j��[x���􎢶K��ёK�E�I�X��H���Ct�S
gij�R��N�ā,/1Us���@��k��l��H!,�y͊�j��NP�W��e�8����$�"��i�.rUk���?���G.a��B�a�s��r검9oJ�~���#�64V�d-rVz:�N������|��W���T��@<J\Y�h&4ȶzbrLK'�������c�.p��Q<?sI7�y�m��q�M�G��d���,a�����L�6�3#^�T��H�&4�([�l��hfi��J����v\E9A�<G�,0fH|l�177��/!u���	s}��z��b~r���Z]��z�.����жҘ,N¯�q��([�=��}ْO+_��	���_�0���}����UHM`&7�t<���Wq����z�	V~U�"�%I�W�'�'���k��J���i2Xoo�I�
T��N���;�R�e���f�X�m3��	s�s�V<���`s��Q���O�Rd��+��,��i��B����%��#R��	��#g��7��{��\*�4�X;�a�^P�$Z�NF\�_P>@<Hb�0�2��:2�C��-	(a]�L�.,A\&�S
祐dL(�Kx�� -�I�hWpug�I��.Zl$A��ԇZ���+�ۼ�^�j�$|�μ.ʽ�ER����v���C= @�yh?E����7'�+���ATz�8Q�Vۜ�Be������]s���w(̮���]C�k��H�.s��^�3��t�~'�)�i'T�5\��;h�r��gf/���2��#k���sKs���R���@�Ykh�)���������Fs�Ԡ'�/�x�;ĒVAG` ��H,/�*w*؆�i�m�f���ݤ��ѧ��	���Q[^��\�-E��Es��(0�֧���L?z�9P@�]gXɕgn�k�����&��d{F�C��0�����k�����Do�+Iʜ*&��l�G��%�ݩi2���6qt��r�:�����X�٠�G��_������O��	��?=͉���RY�y�\9���͝1m�H�*;W����қN�M�]�ݾ�˧��{^W��B�����g�]��ҫ�Axs�8�2YT�%Yڑ��ߨ졵@�
��>E�R�F2,XF�t�L�jNؽ�N3O���$��b���5���4qH��M����C�r�9�n�~�/b��cT�-,_���cKhdwLfV"�0�ҤeF�8`��W��=,K�%zO�������l��Ca��~��l�����o`23��3+`�`[^b	��5��TL� �+�#��c"]@mP��`��Sx��	������A�l*�B0�Lj{f�z8���p�b 4w��B�,$I�x��ܵ��<nqQ�8�FD׵Ʈa��X9��a���$Ce�{夦�/x�&-7nr��[�ǎ7٨v�����=د���fJ�Pi5�	�5���7W���%ME�=����8�<R�X6��j9�b�M�� ��
f���&��� ��6*�}&U�̘tc��=3����C��;�pk̢C���Q�$�-s��3�Y� F�� pt=+�YG,.�;of�^Ɖ<v쒁�3E�qݩ������9.	Z�w�-�_����{���@���h��vQ��E~��#1�b�[�8=u�y��FL��ѯb"5����R���:6�1W�a�O��c�������Y&h���r��+Tdգ��(bI�����-L�r�؇T;�B��G�2��`�1L
�v̼��� ��ѳ%#�lv~=���D!g�9���K��ww�[x��N��tv��ֻ�����K'��O�|��nU�-F�}K&�8��7^��nZ��r�*�4FL�'�T��E{�*��;(�X�����q���u���}.�e@��@C�	�&YL1��¶��CZ=Lf����.o�h �St �2�bߊN��=�7o�ְ$a���K-=$�}D0c^f�%4A�k��h���C�FP������P}p�]���K��x�,�ݕ�qdj�.,b���G������%�}��'۶�������P��¤S���X�%�\Y����'V�Z^Ň��eӜ�3��#:$�G�WOW2hw���uS7��vv��H��0|'�N����h(.�mG�<k��!�X��/"�FĮ�@l�E}�PE�0��F�x���2��YW�q�|��MfR��1�p�&v�p�`Ug�>�Y�c�^�Q:�*��&�����C,pqdv
�����6�[�A���M�zC:*g&��<��8uc��]0@�Q�WN��=a"y�t���Fu����7�'d,�3��굕"�|���_a[�k�ox��*�6A��!0��rHֈ)ET}��o�sX��Y{��
;� U������X������ʥq��ed݌�]��&��ԙ3� 3ɣ8w�y�����mR��X�>��k��q�����"�{���6j	���h��lhL�����*�

Tj�b"K!�����j�<��c���I�~��_kF�)G����&8�0���ǢlE����.��މ�&����V�2)�
�1�uQ�����=CfA�p��5T�zk��0AG.����v��^���$y�2x1SPl��˺ 9#d���4}T�Qs�<!CNJ���j���lM=ɰ��s�vGI�G����]2��9���I����Q���^>�|��rK8\�ę�'\��f�qG�sϜ�}�8�P!IGc��=����1��,8�t+��~8-c��0�D�$���a�v��BlR�;��h�ՙOȩ:f(a�`�����Gd�N�ږ�j���m��h���<ʌ�},旰��י.i	BkI�e�ըFj�f�AG"�X��E��ꤤ]����MqP�3��7�W�p��@Sx��N�$��E��B���CZa�{�Y>���,,��X�(�K�H��sQ����C`����Q�t��H"���TW'?tۀ���@������]�8��~19A�����ki��g�=:@��������@J�1/�e��	2�[�7�B��s�!�Q�rRV�ef�a�mp�ƛM����
��i��3!2Yc�1�	I���-��p�^k|b��qd��E!S�1+�U2��6�f�C��-��П�L�(��U�5��ᖱ>���lc�B��{� E���ps�	�)m�t99MN
�2}!A��$Q i2^4;�ҏ��z"�����*;~�C��յ��;����,����*��(����R��$�x �3��l<��G����:��"�tx�uIEW�`sɌ�\��&j<�|��[Kc_%e�S����_A!���S|~x�����w�G�:f�;�K��j���������R~����_9vY��7����3�g�PZ�o�T=m�P�N�lJ�����uKõ�t'�ੜ�޲n��Lܐ�����o�e�7�|9�{��Xc�	���P�~3�=E�G��굁=��9��U��.��W.~3�)}�F}�m�l=F�Tе�R�;S<�o]�C\���5�(&����>��~��O����H !o:r0���=K���RƆ��&%p9�W��W��2d-eg��Rh�&zZ��1�hy?����4pk�9����:�Z��BF��(|x�Z��M�"���! ��FЃp|��C�0~����P��|<�2�1�}��̜���o���*��Sf��$�g��c�������#}��cx��e|p�W�������w�ѽ��ʅ/���O�w�j@Փ$x�D6�[�����vW��t��@S������E��׸0��-�Dc���	ǔ&���s�Gpk�紐]�Tr
W7���#���)�X! 2;�aČ���9H���p$|3�pHs�^02k��:;�?��U\�{��q��s��_��&nt_=�%|��>םLM ���ѓ�������dr\x�T���Q�W�L���*56�O��㤵]��{�_�A^7a��fwS��9U6G맘�l77� T�_�jǘ�K%U*�-i0�B�7HZ݆z��ĥ�[��g�p�ٓ8
҆%i�_�����Qa�0ꡏ<!�A�)��1�.��#E��L?�-UG'��˩����_���o�%�]�D�;�-^���^��g����1>����Cz���z�D�T�c�D�	�'�^�9��ʍ&z%�'���m=�˖)F���+7�Kd��
r�W�`���7-Y���G�G�P�4u��*iz3�-K�/���esR�y��/%"�~T���Їm�~7*���-����'�Β��d"�.1��=���e25I���^C�O���x�ݷ�7���E��Q���nk�l�'�7@Ŭ-�M�KG>���7�>D����˗ �M��~�D�?�v�5|�{y'���el����o�KK/�k�d�!���+�_տ5���n����z�>�|�쬭:��{#��]:��t隣���(Ǭ5���%�#��&Co>E"�wF*����(�G�3�ia���s;����ⱄ����+�N�1+��xy�����?��_����o��w����c(MN���
6��$Wi���f�&K�M_��Ĥ�[�+t�:�s�V?��D��IܱR��יA�L�V[�X,-�li	;[�(��ج�0O�,��N、|&Ƞޯ)������+4x&y=\�)���;t��5�íp��b�10lR!L��8D�ǼaF�А���i"��^+�x�����~��t	�X�|�?��o���&�M�e�(Ϗ�X;�Wx�����=hl:����*�ꣿ���*�9���������}�j�Q���5���_�B<O����dAO���%%ǐ/NM�u5��h��wI��E<��E�ob�W���>�Y����P�1�e�.��0d�HX� ��)yWU�����=L
���a�8c?D:�F�	�!ED0�ׇ��e� ���i�����'�\~�llo�虓�^�G�x{�m\,�y��rf_8��{���[��Ӆ#H;9ܺ+TH��\j��^ۗS��@}'���k@CB����^��BX,E��xxG~/t.��_\x�vM���/�5�7�7[mW���f��Z}-�SDo\�#U���l1e�'Ԛ��4�4ӣ�Am��Ɏ`'�C>��Pԣ�G�%�%kL!Q����XQr=7�Q�O9!�k�ww��3����Y=��/�~��u��f��X��8�N�jg.�m�`�-Ghw���0'V�c0�:�����fvX��u����,��!F~�X�P��׆�%�ۙ�k��+�Q~r��@`IO�5�r��C::FB��n�ДB��O�X2�'U��$m�A�9�U���=�T6bhV;,�c�	��v�m�ʰW�k�vt^�LaǏ��S����|��u�rQ-7��*    IEND�B`�PK
     mdZ�?���� �� /   images/ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.png�PNG

   IHDR  �  �   ��ߊ   	pHYs  �  ��+  ��IDATx��w�$�u�2�|����n�����`a���!R�/��D]('��E�#���H(�(�D��5�`�ߝ�ٙٱ;����._���~/�U}�S(n0���hTU���2�&ϿYXXXXXX�7K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�} K�}��/��l�v���O���A��'tB�\
(p�s�?{��N�p��z����@^��MA��1V��'���My�Y�����8��j��<&�㺉u����~ �`�tڥf3h���)�3tpX#���V�w�������y�`��%z߃ �j�T��kwe�A��styN|����݉�v���!֕J��h=������8�t:�}��y�`����{גc3���k���ͦ?P�Q(l9�N|�3�Xv��X�~�-�}�{ΐ�E���E_����ݯ�����L&��t6��[�W&c~�w�V���D,��K`	��0ީ�`;����@D �@��}����4�a��Q��@������d|�}�����u�=� yb��~�s������aǇ�}�}+�����t�{�;����W!~ܿ���qpp_!�x t�έ����ƣ{�q���sC0��N���{���sXB��+�ر�Ɋ�d�<�ө�<�O�*Vb�n��~�6��e"�|����@�J 1�vz6��y��#�o6�r>ޛD�����3���c�$��'ק��g=G�S	V�ѱ�Y�b�W��y��Γ�\�:�o�X#@��z��Žp�b�ɤ�5����Ϲl�Z<��G��\3)sV���$�� ��-�
۶mss����~
���8�V�D�z��w�9"���k��MM�$Js?�h4ۄ����B@����u�sd����.��&	]I_5^S 0��q8W��4�� :6��V��"n7�ɴ�)D��FLa��_I�������&�
)�c�vR�͑�X�h�B��T��5�Mx/�8�v�i��󱞬ݡ�\�	�,�S%�� ��-�
o��&�C�Z~D 6�/^�ط�ti�
%'�����$��J�&���l}��0�S24�V��x�]M��yH�O�7�I�:o���ti�IWaC��s�u�e�Qo��Ѽ��~y��uB���x���������1��e�^�S��w͇���-���
`	ݢ�0::�� (���5&8'6�2)D�Y���T��ik���8��k��X��0R��빬����Jrј�:������.~r����y}��>GHԧ��.Z~�!�B7�ϸ�k��&m��)/Zy�Ga��FkRb��I�X��E�r:�mh�B�L�<kL�:��̕����͠i���\�.���{��~���O��*x��L$XP(|��K��q�8�¢�a	ݢ� �j~�תն&R�g��uM���2��d���$}��qj6WM�Ԣ�sA�
S�U7�� 9=�Ԅ��;����K��浘~�fm�aj��8�$t 1x�d�ڴ�Ztz�i����{�{���W׉�ˉ�A���,,�XB��;d�������֌L�Jp�*��	�U4T~��(�XaM��EJ�I0��P�1��Z:2��%I��.C�j���h̖ߠk�A�̱��륅����J��@1���A XZ�5N;b>����&�V	0�~fO�Ұ��}�y��DZp&��{��V�ږ���=���Ծ���N��!��y�S�U����hPL�_GZ���B��e����5����3l�w���ϸ>.+���{��إ����4�[�⪀%t�>D(>r<�W�Ҏ�:��_I�Lj��|o�=y��y�ڮ�2f�EAgݩe��=�6��z�fZ2*���͠>SCO�����ܷR$��ϜS}牴�����c����T"�s�t�Nxdaq��E_a������6a�@�I"6�I�W:�~6��z�%�L�O�e��㨙�\�I��y�L庆�~]�����AS�1�ｮ�m�0R�z]���M�n&R��cZ5�u&3�׫�0�\�a�O:��>�%t����ÇQ4�5I�$�K��K�{�ٮ���ģ�lS36���)p I2�yH^��kF�����^�WMZ5x �O�y����f,A�8S0��G��Ma���k�)0�����j�W,�[�6n�2�0I�!*�I-7i�N�}����2כ&m3�m���fn7䒚t�s��z�4/i��
o�z�� �^�	S��%8�{s���	�1�L���b���2���=d!8N�}
K�}�R�BwL�Wp��!��րI���f
S�6�Q(�h���'��L�:�J&~��^�JHj�J��y�cA���$f���L�ݯs'�G���b��'�!zY:�L'f%e���*�%t��B>�g2ܤ��4���\B��gi����ܟԐMa!�}��'�H��)D��s暓dk�g�Ԏ�yMS}/S�y��l�mf0[����^�Y^5sL�\� %�@���[���K�}30ʉ5P� "߬���E�� �K��Tq3�p%�{R�OoF����ڬ�)�����f~��vS�W�5�0�#)�$�����:�Y�=�i�=�c�����h4$}O��g3'�g�Vp�Xha�ϰ�nяp�����iJǫ?A�P�ВZ�I\fڕ�J�G�HS�S�2���L��s�(�����d�m����fJ�kZ)�H�~}ՊU�u�)�hs���rYۦ�z��I���k��ΡתB��-�ߝ�>�Z��/�z[�/��u�����E?"lkn+�]ajW�XI�dPC�7��^ڥ�&�v�wl�ӕ�A@͘�L�9v2 .�='���O��z��n�=�\�i�WB6]�
�Z�k5����}��5��Ke�sGd߹�����b���XB��Ctjw'	3������g��+O�i���/IȪu+)���{	���oc�isIj�*�$��^s{w�P4h��(y�\K�{��Wб�?s,�C�Y���oaq5��E�!�i�A)�DD�f�K��MB�yAq�`��&��m�@B#Nj��f�c��^��伽�_�q�(v���An��k�e�0��}/��y0��o6o��<�4�;�9��UK�}�j�
2��9+H2�L2O�%M�I�wR[7�bj�J�@2�,y��ħ�oݧ�'���|���kKV�K�;H�j���n��\�`j���n���4oS�#�|�q�8�|���XX�,�[�%��\��Y���)Tz�y��8?�d�v�;ԏ�����s���\��;7��L[3Mٺ�x�3�����\}S�6�4�`��{U��1�
uZ �߼�$�'�yL���ߟ��p�;G���j�%t��C��<]j��e���� -E����׶�f���nf���d���)ᙑ�Ir6߯t=�޼�=�Ǜ�j��u��B��\�@�K�Q�]����H�O^�)����sӱ=���W��-,���-�
(,Cq�Z2.�W���"Ϥ_���m��U`0	�<i\���}f��Ntv�NT	]I����c J�f�[2�[��t\S�7���Ӽ��J�I��YF�߼��4:�ό�7��4��u�U�0���ёV�-�Ě�kX��Mw,,���-�
�����0�\�$ɋ��ME�饻�+�K�(�@Rm�ok�8?ʝ^\^�"�v�yLr+}���X��?OZL���RM�T!�R��s�V�>L�{&�Cy��a���z�?1[��?�����V��1�C|�" �Ѱ\8�hΔr��dE|�h�H��x�qw廤�^��'),ɼ��NL��r�>����֪i�2��UK�}�\.'O��/<i~�m��)Ԣ�͂+���L�I�:��0��^��Nj15V=�Ft��ڦk��t���do��u�͆ߥ�'�Vi����3mM��$������$)��i1�������RX����=��]��*`	ݢ� ������h��7i��Y����Nw������y�߂�$�D	���$�^�ufZ]�y�f�2h��E�����YtP7��7��4�'�l�>'���O�$o��H�73������X3���NW,�[����=ÚM�҂&��nՄ�c����=y�JQ��D����D���'5i3���k+A�f�l"c��z�W���U_?�^��u-����o
-�y�ޘ�R�sMa-���}�nkaq5��E_ap��e[�E��p���&LS�y���)��dzi�I�Z5P9��+�� ����k�R��f]w��nf�q�\�+խW��^C����j����˥�k�e���?�Yά��$yS�����K7�u��>�,���E_��f{��;�&�&I&	阝 3���M�p�Ji�:D�6���箔{�$N�)��J��N���Z�׹Yo=�G�g�t����7�L�[i��i�H
1fj�f�g�}[�r;��yOL���YX\��n�wH������yI��Ip�q�W-qڝW����Z��r;fh���ڹ��S�@PZ��L��p�.�����J�*0���L����'s���d��%s����o]�8'9�y�3e�����a��Rַ��CXB��K���gS�"m�&��0Ћ�ԗ��i6�˽	lS�79�,P��K�V��[��XL�5�j�}i2�MM����qfN{���v�����Z��I��n=7i�75�.�>�mz{����U�C��;�����q`��Fdpip[ˈ87����X:ik�N�фI�KK�2�w��U@�ք?佇�>㈤��=��|f����d�`���_��U�@Q�rǫ(�L�Kj�j��͸o9�S>��9_���9�g�W(⌂t� #.�T���O�V�x�>���w��kXB��+,//;�\&�n��������`1=���WҲ���^�q�c�ڭ��s���I��&י4�'�K�Sm�;���Z�j�7I�k֏7ה����BLK��;3��,W���8������/�¢`	ݢ��ʝ	$	D����I�O���Ju�M�p/B7}�&��2�'}��b z���[�%�s��W,Ar���a^W2ݭ����KV�3K�&�h�A�_޼~�;�Z	!I	�+0α�e,�XB��+d2!��4�$a�)S�����@���v�}���I����<W�LRF�դ��l�b�W�k�uӥ`oF��z�e�W2N�%y?LkC2��,V
������Z��g9���'XB��+��eX��!{��M-�$nӴ�̱z��u�����"�䚺���� f��&�^Z{b�����f��b$z�zz�]�馀b�t�T��ۮ���t���2�4��w��=^i��K�}h��j�d���1�;� /}�$mF��>[=�q���t���s�}�ꘫ���8VR�0���T*�E潄��9&4�ݴ"`��iu9��M���^Z30����t�V"uK�W,�[���ti��P�r��I�+������i��`��_/�r� ����6��X��\��d�x��J���$�꘽�{լW�H
�1Ɍ��1�T��a��dݖ�-�XB��?J���q��<�L��N!�d�\�z�k��u���I֦��js��CۖV�2�+�!`��6o��t�N�J������aV"� lI!ڣ����en(�N[~��S�H	���"f\Z��qh���V��+������f��g�U��|NJ�������u�J�-ʈ���S$/�Jl[t��k���c�(`�q��?�O��ZG��UK�}�t:%�sdm�I�h�	�t��"�Zq�Y�I! '�O+�u�x����)Z�f���^�����lt�Wa�3���m||}֝8}N�	�s෰TE�W�O�֠~�Z��Պ�-;·����l���0s�3�N�i��抇QP����n��F�V�5�=�J�B�?�P�B�T/��P�V�B!UKU�R}уHi�j�I{����U��)2}����E�-��R�
A���>��������|^ڍםY \Yz�cl�,�e��XX�+,�[�2�l�Je���)��K���V�&Ȕ��n����-�f���^���d"��L�J�}���z č�i�5u����MEm��af6��������Io����8|"-^k£xKT`^.�)�I����*	9�J%*�Ã���@��Dk׌���{�J��o�W_}�^x�-:p|�Za��l�R|]A|ߵ�k�Ր�X1gy�D���Ѓ���D���:z
f�4�B:����D�����E��ܨC�r�l	�⪀%t��B�\��Z����U��cvbӺ���B�j�u�v�6 f�<#͜��nD�EQL�ql��q���
��N5�P��Hg�5\���P�O�6F�D��"y����J����4�� �c�Gb� Y��:�-���ȴ����NJ�\*S._�|�z��c6h�5�������ߣ|�.��0��`�@�c�#\�,x��W�b�_�i5=���ߜ�5#c���_�1��[4<R�K�T�\�[+�.�)h�`�`���,,�XB��+3��Z����^C�p��>�	�r2M�$#ֻ�źs�M����������
�Z��]]�!(ཎ���^�\��n�%�D�a��f���t_L�Yָ;�p�O�:��ځ������ƨ֨�u4��m|�R�JK�
��hv�D˵���g
��]&��3,8��\s�V���C�Y/���T�A�p%�^�
E
�)��X��P�f�zT�=���������mh�E���E_Q�Z�K�*P�)��D$�|����р�(����G��u7�͎��˂�(]l�Ƌ�EWG� W�{"C����FW�N���f�K�����Q�������T�\k+luڸR�޹#�	���@��t���0��!l�����Hí�ᫎ���^�U��ȧa�Vå}���y����i�oҁ�g��=*�D�g�L�͆��QCn|���c��0E����n��~�����4::Fs�x% ����ɨ�熱��F�� ��Ld����sXB��"@.8Q;I�ڥӍC;���N����vF�X����ir�2��'��j�3�'���h*��ł�ܡ�5�f(�j&2QÇ�iEѪY+�&+�%���p*�
�t��f��ٱ�Q�Q�xM"���ic�<p%zm�\GD�:,푲�lϏWD�gXcF�X
AcL� T�����h�"�Ʃf�:�>4F�=�w���iZ^�g��јCLʭ����Wޒ�JerÔ����\��C�R���礩R�Q&�s�Y���_��S���Sgg(�_�c7��"�Ǔ����n$lx�}���D���5[��S.�p���J��,���w�K5��[g����\��������fɩ�h���9�5��?H,��X	�t:8��pj�#�����Vgf&�;wR�q+LX��K��0����ݻy���������|advv6�{Y�ó6�l�����PK�-U�ײL�^~�X�	wa~>�R�L&�+�l�^O�Ŵ�h��a3�O�S-V�s-r!kh.�@֓��s���2?�'��`
�2�����(�y�n@F�j������ips5�- �(�L�C;�K�v��E�eQiV���=Z2h�ȝD����mȐ|R�S��%-4C�����{PEǴ�hӑ����|��U�4���Uن�8```@�aqq^�g�)>�M���L���]/G��\wD{wιB�ѽE*_4���0��/0��dm33s��!Uj.�8���3O�C�X8qe칅<�G�֮�E>BY��N�I��v�����^}�����˭R��e��=�
�T�Qw�0pW�s����ń�.//�f3�T+Ԫ���e�l:I0l�e���7�h�Z�l�a��[�u˖����<�o�㖟�?}���7Α���%t�_�DR_��W?���/gg�o*����`���<�V:l�j��j3�fD�*0I�X\51^s�5t�ܔ35s֩T*��/:͖�A�R?-ϑ������@�F�F��o4kN�Q�/�N19��Q��Q7ަ���du�dP�%�zR��Z����Ȫ��W[V=Ό�שּׂ=Cl�oɵi#�N�t���N{b.���(��IQ�h}�l�5��D�C3�g�EU�"|*]���q~C�%��Z-S:���%r�1�W�5�K��-&v����han�i�.��;����04�������|�D�BN���y��)�gs���S��S�8 [��N��=i�`�aÆ���ݻ~�;{�ԩ����D�O粴��D�LZ~K.\!�-��$� ��B*��w������8i1�|?��gY(��-�n�k�mEv>�[�N���ۻ�9�C����>����{�}�j�W��-.�J�����_�����o7m^�%�Ĳ���޻����˃�Vk��Ç��7ަsS(�C؊���hhp�>��Oҷ��=�8;G���/��Ç�<�����ݷ���=x���?���q�ںu����QYfBt�/
����5/*��o6�`��NLL�g>�iڴa�U�Z��]��뻄��������5��{U�&
.��4�]�4�j�u
�t���q-�q�U�U�?44$D�F�x��Tg��TH0��}]p%���ۣX&f���^K9�A���+�^�㮑�Qt4nl� Yz�=Ք�sI�k�9-:�,QA��!t\�8Co��=�܋b����L�% ��q]�ˋ4�����͛��:S,�s&�Eڽ�M*��Ԭ7dm��ħ������w��G���y�ۿ�=��s|^��[5F��y�q�t�M�Ҫ������7Y�*��~�T)��_�����|�����
���e���������'�x��䲙�L���u'�����h=(R��r���M�������h=!knkdЌ�]s��`��y�c�c�.:x� ���˃��B�A:��r+�uW$0,�Ͳ�U&�Ə?�]>�B�9�0�TE���C}��m�F�'��n�i'��_��K2܌x凌���j{��O(�+��Jј��۩t����Jh���D{Ǖ��C����I�yt�qp žy�\(��Q�$�u�S� ���(y�D��$�>{S�ǝ���^�!���2��B9;���v*��G�����ٟ��-�*�**��Pe��$��[n�����ru�,7D-�q�`�;�w;���,|�ŗ��ޓ�>�K�L~�C�g�^:{�<�v�&V��;n��>��O�\���Q�Q���>�ڵk=�ܳk�;�|��?8s���ƿ�Y�����nqY8y��-_���y�s6��ڝ��M���g��x?TG��ZPah�Z��z�-4:2D����^}}��0Cc<z��<<?���S�\eMr����@;v�$��3�����<�����ӧ�+_�
;v��l�@�K�L�e~���􅳔�2��K�3���C��(�S��n�k�X|��QE.Y����&���
��Dn�µЋ�bf����+���U�� b��I���j��~�+h��#�x�D�~�|�v��|\��k�s6^u^���D@�5@�5�k�fs7R�d<�7@�a��zT/.�C�����8��h�>�9��������o�[L�c��#��)��_�_�JR����!�n~v���[ߤY���B9ֺ�h���q�]�];I>k���~���o�����|?�bá�z�F��|x��b�|rr�F�
�?7z�������뮻Nι8u��1A��Y���V�O��o�C�?��/�ȗ�"YX\XB�����?���W�U6��n���GŔ��ˬ���k6��Ke�"���8�{�t��?qQ��a����!�r�z���l�fm�:�����C3~�=tp�>~̷(�"�j���}�O��H�ť}��ߣ%�Ρ��� !d��� &�������!�]N��.^R>���;Z��sz���i$}L�N\n�UK���H�zܰ�#Iq��s㠳N�}5�������\�5棂4��;7��S�}*�SZʮƝ�P�i��y��H?G�X�HQ����]���@J�j�_*T�A�O,��_`���v��X�r�5��C�}��ͤ�BX6%���2�o��*�*U^kF=�A����{$�vn�FG�i�I�|��w9�2z���k���S�������i��8U��|�g������-�h�����j�Ž�e�ڳg�Щ��7�%t�+K��w~a~�5�T�Y��۶�y<oϞ9Os�%��k��)��-P�	iͺ49���ZXb�g! ��_z�&&����,����>�0]�փ�������O���'�_�":�.��?�ڼa���Fu���{�~�W?K3����=.F�ZgͿ��K�+K��&@d��L��mT��T+��Z�s����(֢eH]-��&�N~{;-�h�jZ�m�N��Nnz`��ŏtJ��K�2���t��9�ɵ��VJ�cAC2��H�v�ֳ6�H�	�4���AT//Z�A} �����?=��E�OE5[���}\wމ��E�zq�G��v�S!��5k&Ă��ذ��7nZO����X8ˊV��Ǟ��Y��>��Gi����_�2����������{���a!a`�Ν4}a�^~�Uq��Y�\3N�6��B�s���*��
y!�j���c�bt���;�����N�<}-YX\!XB��,d�A�p�V49�Z�_M۽g/�izf��߸�Xk�h�+��ã��)�3��r�
�"���Y/���گ�>�OБ#G�'O��.^�(5$�UJK44X��w�Z�2�>q����x��5�5I-C�q��`F���
�g2XM� ��t��>C�Er����/���+���۝h���&}�S��oF�'�# N3p��n
,�@�s�~|V�]4�0�J���"_|�.vH'#�W {?N���	5\^|���#�#�-pR���;Q���b7�fw���[�{^B1���
��D@��w,8����#�<Ĥ��V�^M��������&�Q�C>���5����+L�ȴ��ߪ���wA��8���0/YUG���M��c�{�Mڰi3i���q!���XK����'>��o��;ＳI�`XB��8L�^ݯ�p~����4����H^����j:q�I�e������(�?}�ff�X;_�i��(&����ߣ]�n�����ǿ�=���t���={���̌P�ǆ�}qq1�o�|ʤ������b����<���ùV�R��#�G����j��ٺS�M���� &K�M�H<*�ڹAȏ6{|���9�c:R�NsӐv%��n��Ea�c�y�hpD�k��(�k����t��.Ĺ�@*�}��*�Ǯ�hR^�]��5��ڰG��q���^ؔ���[AJ����5E���@�X�`���T��,���}.����]w�6���� _�"a�#��S�@���D�j�����o�a�b.u�)7��N�?�<MOO�w��g��jV����m�x������歛�ο��𨔞��F����X(��b,�[��a	��r��H*�ɤ��a�\\\�%kRn]����o���h��u�����Kn��)B�ޏh�]7G�p���i!�\.Kֶ�Q�Y�.��\�.��
�*�9-:�,�49���_��s���������Y&��Z���;�hJ��a��p����'��JQ'�V�a���U�5S�L��m�6����tk�:>`j�浙Z}Tƶ�ϸyMf�^�|������y�%�,1��TA�7ڙzq�3���FCo��iA���q��
�BC���r�"h�ș�}�X?N$Dէ�v9�.@xy�j0�Zx����������f�I)�@���Ay�Z�*�T�[^*��=I/�D��̧D �����'��O��x��yI��K���z��H�#E	�k����_����ΑQ��AD�#���n*5��]����������VKLLn�����Ҧ�[�Y��'
�H@?�.^��B2p��:s�^۽�j�
���K�� �k��=�Z�n=���!?����+/��}O�x����KD<L��st�軴qӇhna�G�i��[�!;L�|��(D�q����\�j����!���:��N�Q�? �̀2�L����bQ���A�J�~���6���l �  �&k�n[����x��<"�V�%�ZjǤ�ׄ��K�hPՋk�C���+`օW�@�-�����t,�(`N4�x�������(�)���X��m+���R���6�F�~"H��ި�b�H-M�	9�u�y��Gr$�Eoh��B��p���%*�x�t�}GKL���7R��=��T����c���� �ѱ!j��;t� :�.-�i`x��Yh=r�(��{�n޹�ҙ�r�Mt��ד�ɓ���t6*���tgN�����4<>�F|[\������ }�̅��� �����EZ�Zs�0?؊��5X�L����G�й�)��":Ҏ��\�����/��بhF�3������%-�ԅ�%�����OĜ�;"φX���2�+t�u���Ҳ �6�f���ԕ�l�\��U�k73q�+ZG�6���u*���Y��v����њ������L����;C��v���|���k���\�Kݯ0-m~#Q�q�^wg�-�E�s���y�8XωL�QZ]��RD�5�q�h{�`a�Z�ڨ�'��/./���b/�Tw��qZ3����RL�Y&�\#2&J�������|\U/-�Ňze��@N�U�� �w����7ߤ?��?����!=���i������c4W������|9�<_W�K�`���oұc'����䚍�b6둅��%t�ˁ�Tj�o� �Ӌ��K/��r���:�$����iqa��ܳ��.�H5�lf��&?�Y�	tp4Gy��,E��3���o�IkV���jZZ*��e֐�D�?�O�^GY~����8B��~����\~@�Eg�>eͺ�KS�8��9��_�7�BSr35֨tjK�H㾴�j�&�'��a��@�8�^� z��o�~U?=���f���J�/�'o��5�O] ���ܟ��L�ױM�4�I�����y�%��M.�rw�.�v�~�f�)"S-��`V�B.G9�N;J����4><A�����iav����_b����>Agϝ�7��w�yGb3�x�	Z�jU�KT*-��ci�7�z���P�{n~����O鞻o����(M��S.�%e����O?K_�җh�5�K����ykn��b��nqY(�S�Ԑ|m�.�����w%O;@����ť
k�5~��)�
J���$�/��昨���O�{�?AϿ��<�gYs�,���G%b��AP��͛7�>�j������{��s���j~��x��u(3�E~�CQ��!�9�qw
����Y�!�n��ܮ��ĪdMv�oj�Jت�*�����?S�0k�����rş
"��c�<�w�����v�w���5�N�����։��<�fԒO���Q�zJ��-f)��2"/�`����L����T,��ԉ����O���sHS�s�GUC�*���ɓ"��_����.),��kX���p͠ ,;��!`�����[X��ﾃ����^{�mB����oӳO?%��쀜;2<�6j5��[\XB��,�M/�*g)��d�e�D{�6Y.W��K6�c�J>0JgJ%�zI��a�_D:D�������}�8@��� k���*��U���v�9�����4>4F��������>A7�x��� ���s~��	�n��T^�*k  Dg7�N�SC�?M���XK�cU�N��e�A7S�T��t^ՔM�TI�$^@ק�����?�j�f�_����յ@�2�Y��ټ~��c�V����JۓA�f|�nBפ�)k(�vʦ"w���0kη3����|U*�yg�MASoI&,<�y҅e��۷�Ν;��k��4��[�I���7閛o��o��^x�%:��ij�>��I�{s����[��>��������>*�	���3��7_M�����\�����nq9pʵ����tAc-�^�֋6�.--.	A��Y,���d��$�P�֨H�mDIW�ZbM禛n�����=�Kj9s��L��}o%��^���w���Z*f|)f��I�g#2x�7�����w�:d��%Q��"nq��^}o���ҝ��h3�]�G%t3^��$�9?W(��:��c��Uc7���@�K[�y��9�x]�I��i�4y�>��M�B��k\>f�8=6ſ�g��Gz���ׇp�V�J�����7�=�8�Nж5�d�w�c������4;v^��y�ݴc�.z���rƄ`�9a~G�·�~��G�h-�ޖ��Z��*�\�m�M!P�w��K:ύ�,̣]+���S��F�f	������ ��f��M�F��%��Ղ���|.�J�Z���>{�5�j�$>�@����T�'�|���o��hHo��:?~�6m�D����<T׭�������t��Yj�pL#������n��.ҩS�����t��m��d�噶��1h���'|�(�ˌk�t��L�6I��6S���J�R�<&�������@&:�j�*$$S�ig��6�h�H�dCRy\-b���/���q��՜K	zK��D��ս�׉�@�Ѽ�5�;�j:iu���tM$c�(���I��D�T�tu��(��rs��/�G>�(��y*U�S��W�H��Eɜ���.����򒔃E5B�֟~�iz����W��Ⱥ�=h�R�h��$-.�Q>���4�;�Q�_ST��PXf���i��i�P�����K���r���f��?�
�<!��Zm�$�F��(0�7#?6?�)��j��ޥ�j�F�/�?���?���\��ڨ�m�R�0N���:M��H�^���MN��\���A!{�ߕ�83	y=h�)I���X�M�֓�x@�H��S;6���sӇ׈W+�F�d��e��a�+�w6�&�(H�ى���4JQ� /lG��K�Լ��c���v�w �A�Z��5XOץ�xd.`.�R��@@P��N:���8��M�o�{���
�܍�Gz"\n:N���b��$�:���A&f�{���c�������~�Q���3�o|C*���� �w�&2)�kKT��k؊�ԛ���7C|�Աu�p``�,,�,�[\�t�s�ߜ�����/�F�N��9��J���P�8 Z�~QTU�2�䙤�9L�z���!�:�u&X͛(\���%k~y~@S�lzf��� 06:�дDʧ2i��Y����H3OE�A�ބL6�A�Z� ���I� �B4�.�	���y��ZA�J� �7J��4�q��	!E�����:��<����"�A�v�F�ϝ;'D��@4�V#pD���U�5������/�q�et�=66&���־�~s#�{�ڵm�u����h�؎�D;[��d�ǅ� �m�و
������̸��d�A;�I�ZC��!j�[b�q(*��Nli����ђ������-��Q�M�@Θ5	�z�����J����\+� ���K���:��XM�c#�,�����a�rr�e���@��*��UT͑�A���?jǚ�-�,�[\�V���C1ۦ��*���L ~`��B����9y�#��4hphH���Yj^A[���S��pP$��Q?�=�V6:s�>e>�J��L��ǩ�l	��P�̉�n��D]�🙶%ד����0���)aj�N�x�	Z��	�*�$-O�zzZ�� Q*]���2D�si=55%�A ��8-ca����T����ܸ�07��5a�J��hq� b�T��c��:u�|iÊ��>����Y>k���z�F��ɀC5�'�Z;L�)�]��޸����a���~�xO�/y���D����o5
D�C�y&�3g�IC*�u�t�
�'Ȣ�h}�kb|�D�#���io@R��>��2��|���NU(��r�a��~��W#ԪלFʳ�nqE`	����='�af̗��&��TC�(�_+ʬ-�g��͖�ة��c3�ѡq��Qʨ���gL��:�hA
hԂҚ p����L�\���OKO�ŅY�[UZX���N��w]��ב��x��U|�N�J����,f���)A�I��krE��� a��2�k��3�L����眅v;P��Ql���=^�ԥ�InkA*n��?�a>�h�<>��PFB��&˿�X�d�&v@��T�Q��A�P��0�G��p�0?����l�f e��@�Pī����c���[9;Qe:���j���9Z3���p7�� ��*�6�d�������ȉ@�, ]*�a>M^�y���f<����s5J�4�j-�_��V���:��Ei�[a�gق����|�5��nqE`	���X�E�O�����kV���~ ���^�6hfv�*���F4<��.ʀBkG��t���T�7��s�hQ�ҍ�m�`.���Ξ��'�={߈}�q�r��Nd�ad�w"���|�hC����L�e�`s)�i7Hfp��uJ�І�E���8l�x 5]�O��j׾���\�,������A@J�.�8؇��t��bN���|-�P��=qC��~# ���5��>�|����{�-0���A]Q���fLI�us�̵����0�[o�A�Px�&��'��,���O��@�
����
W����Y�� 7@Y�m[�R>�e��<mݲI�ɞ;{��:�{�=416B��N�!��I��R�AS���w�����+�Hi�L��|�ZB��"��nq��a�dL-�C���m��o�Nk׮���k����1Gg�]��}��x�mr򞔇-H-�r���ڲek[+s��[�J� ��w�#-]��ffifz���g�'��cߣ�'�������[��v�����r�)�r������2�$u]��_a��i����A�0���N����Y&΋g�T-��`����6�����p�q�@dW�Uv�1j��l��x/�&��T0��pm 
�b��64{�?�y\�~xh�H�i��a+�\%�F�@] �R��9
��v����W�y�5n������6�K��,��R�����4u�<]<�B>w�,=��3K����ܢ��M�
,X6�-�� ���K��)�����k�;��X^Z���c��~ ~�jy��n^ς�(ҺM�%�"��"����i��h��j��^۽O���	�����/��-.(��6��26�_G�����k�F���t��������}���kߢ��T(HC�Rm����v�Z�0�!:s�Ů��襗^�`&�亵�jb5eL��)�������f�y����O=B�Z��8L�N<.9�R|5�Z�Jz}I'�D*��ǭ�ps���G�ڦFʃ�����-U��h4;� ��B ��ASq����G�Ž�`<��#]��J��G��k��\��1>ǂ��'�F�s�.Y��A��g�e���5�j��=��0�[Ҁ4UH���=ւ��K#�;Y�J}�I�s�/��, ��,4�<��������O��o�7���˥�T���	*��Wb�ugffN�;o��~��TZ\����Ī���3��*ּ|�A����|?.�y}��t��Qz�чYx�#Gܸc��AӧM7\O��ۿM'��UX��-�[\1XB��,��ړ6�c���|��%���1�X����J��ŧx'k>��[�A�g�����qǪ�IIW{ꩧi�����O~�^�)D���,~���"�D���?7S���I�|^_g�E���6m��[n�I��O���-I�#R�OjJ�I�F{ϰC&f�RӏnV@��r�|����g�-�F��6h��Î�a;7[���A�J����@z�m�#����T�q��u=��q���! ��p.��8>dh���T��k��-�o[��+�;�\��5��L+�����������{k��;�a����${��e�,HF�wO�Q�@��ч?� e�<�w�,m�ϨP�֮R��0�m!��ý��;����sld5}��_��?�Q��_�R~����/�0B�ëijvA������[��i�P$�5�ֻ�{ﾇ��ē�d����[\)XB��,�~#@��T� f�뮻��P��	f�]�yW�!�?�SL>6��>p?��o?J��6
b9@��v"@�
A�m�-c,J.���j������>�0?�ΈFU(f�_���~ݒ��3��bM@Z
�:A�Љj�JJx����daw59�L���n5��XA� ��; ������&@��Zs]�� lc�
x�ڹ��q�@�8�4j|/�z�{ Q�0�C��ZtM��@7��������CP�!@hl���Ƽ��콶��,/�ף�Lw���	ݗ�Jt]C �7��T)U��/��mظ���/�kHf�\Y��G������Q��ځ{X'~{�j<��gŢ�,h�t��i�p�>��l�W�"=� �a�&Z31��E���y�vA~���(��W���;�S����tϿK�W��-.�ۅO;�j����p�a���;y����8��a���i~(�u���7�l��y���K�=K�s��e��wv�&�?$���#D1>2*�#C�Tbr+�1�j����'z�]�b>C�����\������S������P���u@��X�C�<�5�ڌ�6K���u�C��~5�G)_n;X�
�D>�����|��LJ��&'W�M�����NS��#�t�*U� P+#�e���9���j; �0bR�3H�a���"�]5��S���Z���q�q� n�^��0&���@����v+VM�����oetz��v��YS�\7�T��ϑo4ɑ�y5��j���'U�a�r�]��8ZAnUP�J��9���^3A�֮�����ݽ����>�c�:���������]���֭��k@ϝ��o�E��:�o=�m�|=}�#S�筣�L��]K��"F�EK�W��-.���M?d�7*��o�;IN��~�cZ̈́�<u������r�J�ũ!�|~��e��i��7� �ѣG%5m`t�����.^8O�s����5{����ڠ���;?M�cC�/S˯K[SO��衝��{��}�ș����؜lV�k_���,5W�� m5f�5�fv�ݮUڎ9��gMV�i���,�6@	O�X��j� t)��s?�� [	*�ׅlUyC�W�Z�~���ڵƹ��5� �jAP6֤�5>k����jzZϴ��=�֫Do���:������F8�ʆ
���'L�0����R�X�_�T���Ւ�x��)p��6:q�\?���5kh�����7_�u�ޭ�\E��O���G�Ϝ�\6ł�z��2EI�sR�D�� N$�8����2��nq9�0��>�úh4s3Ӕ�f��i~n�����W�v��H�=.��{���{N����;?po��vz�#QU�� �l�N�<A�����4xߪ�	�������THj��{龻��kT]�r{�R���(&�$ȇ響���*�'��-G��VJ�J�J� *(H�y���Ą�𑛕��͠)s:�Lˁ�X�y�puΤY۬O/y���k���OS��":j	��e��v-���ɼ}�,�+��ldd2�.���G�q(��tM��dHd�iO���j�s3�4;=G�rC�06�+�y���O���&��^x�9jv��N���"��5"�$�mh(GC������X0am��p�dYhh6+b�A/��:�l��ŕ�%t��B%Y����A��C�R�jҵ�ma���C٣ֈ	�a ���4�Q6����T�:�Ľ�����7�1ڪ´>5}A4*͡_�J�������5�Il�|��!�f]W��)I8����x�Bk��m��SWR2���6�dj�i7����?��>-���m�u�p�����M��W�h{\�V�L�V���L.۾^5�kKU��לs��߁��ֺ�f�{uAh�\�oj�0�c�9�ɪrz�B�fTX'��a����rÕJY*��9�=���Ϻ�&f�q�֭_O�B���c�i�:�A�/������<���iB*杓 �y&s�\�����}��>x��ZIA\@t��*);\��(ǯ�������8�?�^�y�W��-.!���-��=�p�"�~�ڤ��"?<S�.�6<X@TuY���/��>!�a�ggh`hLH���)����h��v��Z\��k0��S��|���.��C�i���X�g�@�s�Q�V3�������v�Ͱ��	C5Z��}�g���kf[O���������[�ӂ1J�z������4`ѹ�R��6A*�뼺~�P���qJ��5JT;k�:�j�07��R�M6�QAF��,��^�������"���%����ϝ?E?���Ig��>D���,d�0�T*-{��v1���[XZ��������F�~�3�,�4���
�Kљ������m�l�M[�Q~p��<VynAH��{�ї��Uq	�Z=B~˵ڹ��%t��B.����`N|�G��'����LHn0�����f����Nh���rl�T%�3��v��@w�q����K:}�,}�_�Gy�����~���Lsm"D!2����9:��~*//҉��ӻ�f-~��9�̜X�4R� ��҇�'JBJ(&�i'3���\͈�6��A�2�R�v-{��ƫ��U��:U�4��j%�>��5�P��V�3�T+٩6�&6*��Ĭ�T�f��ݠ�ٙN��o��Bh�>����V��R��1�G��:�n�4�G��ƂD���ر�t���t͍7�Λn��3�,���_�N?E�\A��B�K�B��z�6	�3ʝw��g����e�R����G���Sg���i�Y��3�ghͺM�~�VB~�=����<L7n�L��l�,,�,�[\�t*̡�K&E��(Uʋt�0k��52$���k9>�=3EKK%r�R!Ҋ
Ei��t��{,�&�=��o��vj�:��P$��������@���?��?��2���@7��ɚI��D�ݔ�W�Z�ҭ�:Z��+LӹYM.�+����T�ǘ�]�ES�9�i���ꀮI���J�:��6�s�pH��Û�f�5@����(���>j�[�b1�=�*8��L�[����9ӭ���s��"s7|t:�Ha��^qh�Y;A'O�����j� ��A~��%��J :��ZPX�RZ���Y:r�yL�CC#r/~���s?MK��~/�f�;�����ȱA��cg@���\%?D	ڷi͚��v�F���%8ך�-�,�[\�AC*���$ZD�܉���S347��O�:/��+�:kDc��f�R#Ҭ���i�y(0S*W蕗_�W_y���,�2��V�i~|{���r�e�yRK:���˴cǍ����o�C�N/�������471Ӻ(V�J�VikI�&Uͫ�4[	�]�5y�Шn����怦�Z���k�9�'nV�ӆ)J�j���7���樫`���y���ZLBo�Ꙅ-�E`L��G�m�{���G�7��Y]	����Jz��c,M�S��4�K�b�M��K��w�}7}��XGN��<'��V+�4�����bA�_z��bxp@����-,�.�K	Y�I��D[MH�N]��jm�̖�iN�ފ;�W1�Wh|<z�;;eM�W��-.��v3�Ji$��VA
~��S���d�
��Rn����Ayx�3^�i�5p���Jb19(,S��Y=d�
�먴���(>NM�Z5:H�l�D�X+CT�7��5z����=!����FZ9��T3����oZ��a�V2Өm�L�7"A�ۡYc�kQL�МAjp5�@� :́kX�ł�Ħ&t��!L���	փhl)��k�l?t�́�i@� �k�Z4?��k�mWn���j�܎f�k��B��@l(J��(�1�U*���P��D�z���6$����nk��a�o�!��q�tmS��8��L�?q3 =��ãm���:\wq�(������)����±���ޢt� �3�?��~E���؂T��� �2����x��{4�.�p�,,��	�w��?!���>\�]�q��nq�`	��P���VMM��� �W���7�I�S����LL��z���8
�t�J�=i�(�&J��>kU)j�q9Ҍ�Z���m�y�[�_��I��G��g���ޒ�ѕ-��&1â&����a�w��(��+H�Asz<��ig4G�� ;h� q�F��xt@���^���A�C���65_c-*ས�i�=lG����b2 �믿^�}������8�����W\���=!kT�{g��v�2�6Ղ��o���Ր���!��Q�Ns�a�Fj�j�X/����XG�]P��ZF�"(��U� �7��dh�+ҧ>������Q���Q�D����?��,���Z���i�8 Č@�k��fM�N]8����� 0:A_�S�EZZ���6G�`)I;n�V���2��nq9pJ�E�٪3�c��+AO��e���.�������Zk٥%֦KT���\Y�q�)1a"�=�Ht<:�As,2���}�v����O=��>+���	�@���!rR^L~~T��Sm$�&o�<��S�9A�V�7֏B/hJ"u�y;��Z.���F�s���;w
Qj�t����j*W39̿خ)e �� dmӪ٠c�Y��0���\��� ym�o߾vԻ
X�
50��:!L`-����Z������k�=�ڱ>3E��x��uaM�>��u�b>�W�U���^�(���>�~3 /���S:��X��k�;�q�@긞��X���Y?��5I]k֣�>D薗�J�bz��� �Ш�4p���t�a���؀�Nb���/��-.��8�Y-�JMʬ��y1�%W������Z}�&�ի&����� vRQ1�N��ÜJ{L	6���@����.=��T�B�oP��xH#�	������ԝ��=f��܌�ƫvR3�TۡjG4̩����5�\���?҆6��7HS΀<p<�h���p��õ'���A, S�w��@�IA#��0���b)��p��C�W�-�}�Av�
�q��z�5��}hyX-^a �n-=������=ý��m�*�l�sDeg�m�J�7S[��ie�P,<�]-�jTp��e��G�V|p�T�45=E��%vׅ�������v�tj�r�ynn&"�'�y��+�{T�z�"��"� �2�K�����ϝ���Mkaq`	��rf3� ���ԯ7(�e(�� ��يs�s�e�N�Q�K|�yt[.EiWu&M�	OKe-T`�����b���V��fMxl|"����СF�I��}br�F���%���ȡX�t5�}��ԗ7+�)��Q��eL5{��j��󎘒�l�B�7l2��q�|aI�(�DM	I+!�O#�A�Ђ�>:��8�w�Y�� _�	��1 V ����~Y���1��QA@��U�6۰�� D,�mFq}���\?������!ta��������
0؎���p�l�d���;�[�.�v�K��-|ϑfL:�e������xL�˕�\����]���y����@�L6O�f�*s5�f:�G����-���-Q���k�Ã!�:�[X��%�sb�Z� +V*�8�Ҭ5�[\XB��<�|֩=�,��-��Bl��.Q&���ay�H���<?TYE���&�x����Ai��mq�F�6�˃�R�Iz��ML�w���z|O�{����?BǏ��#��VщS�������ж�ү��7z�fW3=��íU�T[�A{��)O U�����V�ѐA8^���Xq��Kƹ�r��� Z�v��{=����\4- yb=�����5 �hx��CH@y]uC@[׊y*d`N������u�ݻ7n5��8B�^��z1�F΃�!X`��b�;�x��c��N��1�M-*L�i�F�ߝY{�y.W�1�������hb5:�-��h�����ߒҷ舶a�&t���o����JK�|�}�Ek��ťYZ31)�t|�^�uӵ��{"�LL��S'�ҋ/�Lo��UYXE/�ln@\@W
��-.i/�_�ү�A��W�Ѻ��Yc]ÚtdF*ϱ�NҾ�(���R�.~uԿ��3� F�w�����n��&��^{�5:y�x��y7�&���)��_��^}����~`��m��T�2�P��3ڦ��Xة߮~t�N5�J{xk5���OM� 1�!�����YM� U<����4�P3�F�ئ��Ad �(�)�kBۧ����؏��G��o���:@P'N�'�	"�g�a>��B����{F�u]g��r���� f 3�,��g{�3۲G~�=�c�zoyyf����i4��%Y�5%���H1@�ȡ�:wu�������/h�������]U��{���m�7��p����1~0>��x�
�yC��a>��1����x=���<�_[���؏���
����WߐB�!���5r��{F������{$��Y�~�u.�t��
@ٛ��r��1����6g��Ћ{6v�O6oZ/7ݼJzz���d�9Y�f��F�����ߨ�^�����x(�Ē@Y 	 =��}��6�\&%����Z�T����5�e���j�$�vJ�0,�8n�>/����8yZ�z-�n�L�,�i�,W  a���k2|��Z�M�-�d�҈m�ss�����%��?��n�enZ�@7��iɤ���w�QL{>kIT�J���O�B���-x ��HaQ��� �q<,b?:c�8�mT���qt��`�ê�2^�Lp\k�� �� �x3�`Ȓ.$�a��F���kIx�7]�q�q�9"k׮��t@�A���((��c�V����3��7 󇲀yc>�s�3y�Ix,q�' c:w|��t�໭꺀�?d~d���ZU�o �ݿH����}��N���Ke��Z�i��`=O�:&��.�����e߃U�-Y��7�~ʵ�����&}�yY����Mal�L�D�c|ܚ����ӑͥ#�n��  z 7"���c�!�bHDK+`-��W7ָ�Q�-��ͷ�*����;����c#j�'�@?Rm6䓟���~�!k��M������铧�i��;���j��Ւ�N������wQ>���䳿��5f���Q�/��H]��G�s�6�P�%���pOs�S�����t,`�2��x �� 4 {�8�:���}�k�=W�6�d��1q�J�o�}��	[x2��q.Y��j�y�`,($��� ~�-�� �
l59��{6v����=�n�]�9p�P���g��kbܸ7�5�T�j�wIE��x(�����'�W�$�u�|�-�$F��3T/�$�M���-j9o��n��Cr��ai5U�ץ�Dc]�I�}�z����m��f�������/��ݻ���9L�]��>7s�Y��ee��AY��_�z:�83�ٴq@��تKT�t߮j���u.�I �܈��h�bc[������%C�A��$��k�����+�m�WR-�n��&���'��ذϟ�`�NLM˥+W�.��
v.��X��1���VT�����m9�ǫ�t��(0p�����%.��F�r��g&�o���d�lȊ �;�����LI�1���>�����u`�B�ą9aL�;�.g΁ӵ���̝D,�����b�Z� [ 9�Ͼ���91�৪�S�����-R��������<�~�<R�r,�^��� !OD�1U8�^5B�Q3R��n�*�rSj���w�]�<Yn�������i�ve�`ӫ��:��x���b	���>����MOMH�<'�|F+�o�}��\o4��Lܼ�&�*X���l�B�}��e�&yg�>I�s��TK	d$ �@nHԊj[[�Hȸ�S��Y��v�:��<kVؑ#�$��I:�77������v;$_���dz�h	I���ߖ�}�s�A�g��w��׍��ʞz�r��I��ްf���o��*!�xaX^~����;��V�r��%�)��BT;�i4e�Gbr��]�~��N�����y��OK�#�@����Ke-�?���8��e&�Y�g	�=�1vk�X�����R�F�rB��{����f]=�_��gC�X�Z ���[��dcQ�y��k��1�����ll]o�����r
g?�*� JW�=K��-˷���Y������I�'N���B�fJ�{a�U���ܼVR��?����MYkU|���\�T�ɤ#�N�F:s����eb� �p\z�ݺ>I��j�/�g������@dA$ �@nHb��'�1�eŦ�z�J�hԞp#6����� �b�ڡ&�$�K� 6�3u����~����,f�?{N��OI<��.���{g����EK��=��#�X�2�K�)�F�$ �V��Ao4��}�a��u���Bv@c{M��!(�rn�k��3��{�{E�P�k
C�f'ر�8A�.�LK�O��gR㘘k�	��f�cl 8��������@���Z��7���M��̇2曼0�nt��r֫3��z?s��T$�� %��fے%��tF�i��rIx��a,}��{�op��L.o���vx2�9n �w��=�>�x�_�IG�oH<��M�2c�j�WGep�r��u=��(����:��YK���,��ȍ�1 ���c�`j�\R�>uB-�W;�֗/_�%�VJ_�"�\�R�+;r���e��2�]��G>"1��''��z\w��^2U�2�a�:(a��{h�
7�����+�!��1W�\�u��>PDM�Y�`�� ��d8Z�tZ�x�aV53�	��o�����-�Ы��gĉi�����N�8���<���L�|q9��9�dXF淎	�t�3>��+̪��2C��n-����{+��p]�\�:���ߐ�)J�k���XƼ&0�rP �#����H�(�kj���9 >���)�#�ױ�M���qDF�4�8x#�� n���+��A����>|D^~�e���;e��-�ç�r�}��?=|R�/��3�N�[��Z�h&�0 ��[�D`,��u =�� ��!i6��rI-�j�a�uɉ'��Zg�Р%�V���&��-��sH��}8�$ m�m������#H��hK�9l	_ ���|O��%����\�s��4��p�6붏��\tk��Ɇt�G��m$5����/����mk
�;���4��\j@f:c�l@��76���c���8��0��3�� �� ��M�y$͑U�$4L@ñ�Nz���D)��A�;��?�JIg�S��;����:בY�%�|\���;�1��/��w[���3Ш����|�N�
[.��RѶ�� �QW�N��qIe�v}xmp�'N����[>(��ה�}��V�0::"��w�����ټ*ӳ�t�m�t��ZWn�*<Q�_W�����w�~c��f2��` z 7$�x�����hN7躹`���Ro�d�-[�"X$K��^�S0k+����l�Y���>�������-[�X��p�
Ӎ�1ʫP��|I��W�l�`�ks��e��$:�d7�Qʺ���9W�|�pƐ��q������;��߅?�F@Cf9����Ը����\�.q =>�Ŏ�  �>$�A	]�T2�99�i�C��@�"�5f�c|�nn��ٞ��q?����c���y���8A�>C
�0n�����\����� ���"�M�{%cW��t�2I���F�*�j]�كb�g	J' ��	�&��߿h�w�_�x�	+���e�0s.�Hw�¨��Cv}$š���
�f۔�}�|�w�����س�@=�� ��i�&��F��lr�`1}�y��2vuʁ_;b�@~jz�]��Ue�c=��o�T�}��5�ڹk���~���G���~���p�������G�J���՗���~X"��D�I��B���xC�q\��<��T� ]&k�"��&�ӥ>11f`�dt%�w��~�qҳ���ZHR�83�r ��f�o�����w\c:��O_˄/(:P&��F�<2�� Б��'�aKV���(=�>��^�U�)[�g�3�pe���a�����~�3-u6��_5��0K^�r��q���^��G��D�m"t<+�u�<t�Ø�0&B9Pn�xg�S09*��+�"w�q��A��K$e�P����c���-rX��|wV6nܬk�Te2,���S�"�/���~����#4Mc���@D@�%���m$.�V-��2Z�V�!S����Ε,�<��r<���F�o*�5���]����1�W�25>�m���'�w��]i7ʖ���d4�.Q��m�v2��*�u���0g��ē��mvs��-.�����@�Ns؁�<0�n���}^�2����ܯX��g}�K�,u�ϡ,@8_�3,K(2$g���|�;�	�������yr��2G<cB� �+�0��{�"��-��Y�w��>���<�)>_���̥jqg(p�Ƈ�B�7&X���f�SI�wc
���V�,�B��C ;jȹ�g�L�"�W��3g���}�h�z7�Z�%�d�˭I;�I����կ|�~�a������ܹӔ34���܁��9yg�!���%K�t����V�����,@����i)(�������P�a��//�rC+��H(j���*hI�27S�M|�I)V\��H4nq�t������h����*@��7�f�M�,)	5��mboZs&~�ܯ�뺙7䞻�Ƀ>(��#�j�d��K|�t��5����puG:q\��b&&�@�% ӵ6~`J6=k��C�=d��e�밾��n��Ų�=��q���,Py�+�1~(� ���)j���*+�L0M���"U->��
�u�s;s挍��*�}*��:!.���.�����L�u�]az5�h�K�h�`����2*0_�W*���b,������e�ݯ��J�e��e�ۗ��+6�?��tqN���)�֌��{�]w�}N�]��c��SO�Z�;ԕ4Z����5̤Ҧ�@у��ʌ�O�șs#�R�$��Y�v���{{��Ϋ2��	��Z�Պ'�{ "�r#�N$�usѪ��?��u�n
Ec��D�`��?��mVzċM�JE�z�M�l^"��T�������Ę���*	U�(�R�������Z�N���ruΔ�_��_V�	ɾ��ɏ~���n��w��KtC{W�x�ǵ����~��>�W��T B�^ԫ�F 2����pX��i� ��=X�lU�>��&�>���L�3B=��t�x1�6�{f6==�Y��B	��NkCQ@> ���Oy�^�����r�0������ �Cс�Ƀp�j�`��ݿq�FU欋M����׌+aH��6�����ܶm�ʣ��P%�c]��eK��E��w	��;����K��F*�����F�}�ګF"��'��Q�R-��,����^`�.�ٌ~�j�GR,U��j��"��  z 7"�ݡ&-��Y+�A�1)K��ܒ����H��;V/���u�ι�bu �(w��"H�R�R�X�cPn��;�Ⱥ�vE�򕿑��iqUk�j%i���=weW�N����3#,@��nn���x.��:3:oX����܆� �{ƹ 
(%d�㸴�	���c�lU��������X A�ɘ5���|�L���39�1_$�qc=�1m۶m��p��rW��}�L��~�^+T֔����{G ����� ��q߬�'3�{p��x�3��y�)��U��2)�e�T���&"���Ay��J�A> ���:gxQ�!�r���Gh�!.�3,Ux���ǭ��,����7�(�I�Y�^�_���ju&h�ȂH �܈�ڭf���jy��F�2�K�<zOXU��M,>��>��,؄��0�F�q�S)�f��U�Y�< �;sХ��~�������P�|�%�P(ֹ���[:NS7��3��]�b��@��0�nm��
�T*�bf�O)X����0hwR�B*��5O���nu�����0���2�O��̰|͟�NN|�� �iUc^p��2߲e��+z׮]�����{g���sz"0&ѰU+����w�m�u���<P ����~B�s�:�����c^���FA�zUb�9AC6�%��~!!K2��q�6z�SO='��3
�.\���!��s�e��%օ���9b��Gd�����m�L��G��q͚Ԑ�����Gm�Y�������&��=�� ��!���nj ?P�:��%B��w���b���־��^]7�e2�? �.M`n�ľx1-�P2b�VK������\�l�s+Ќ\�h;J߆���:�%2?g��,%�H�X��1sl�$���i��}  ���K�E`��L�c���K�3���V��q���� ��x��O����
�6�,7�1Xg���F&�: ׄR��qx�Y��2`~��֠�)W���a%�����G��p
��>�ϵ��]?ֲ��}o�z6��(q��H�B�	)�N�2�x�hX�W�,���rU^R�w�{�'����L�x�]y��1'��9.�X$���g�	oB��G�s�êςXG/�����O׫o�@dA$ �@nHP���,�����z>w�PXM��X2e �%�B�5��Ջ7-�)�Hw Y�`�{�jV&�{!  ��,�a��*��ry�6f9v������<d1t�p����� a�.,QX|���6��Z	��W/��E�Y��'\i{ �D5 ,E���i��|��� 4�B�>���f�6@nn?�K�pM2����5��I�2�kǬ{��������`��&s ��qP"�tH%����p���?k�}�y<��4��yT�:�x²��N�d��K�;�����XN�"�mR�.��;l�!b�/�����ׯ]k��{�3x��)8{�`5�΃ԒJ��VwK���)!ɤ8�d���e�G$�Ey�[m�ld����H �܈�"�1H
����zvnF�
3V�R�V�����4tS��֗ؤ#)�����aZ��j˭��*"ⵦ���{�ڐ�&�zuī��X./��\�����n�Q$l���ߪ���d;b@l|�!�&7oYH lY�	�Z���m�9D:n^d�3+��bdCR�2V!�� Fp��#��	`$�A�5�� $8����j����!P$�����3���@@b�=���������w�m�I�,X1���i�צ�zN{�~�ܫ?�MJXZ�lC��x����j��N 4*#ȋ(��V�<X�A��i��E�I)*�cL��o�v�d�z��v���RG�s^�ŋ�����$�k<��xĞ��*��ƿ�v�Ʉd��JyF-���������g �ʤ�[S�G�}&W%�$�le�ʁ -.�� ��1	�"q�v�V,�dnZ�c��Q$����vX6��d�'����%�8�j�q9y���1�4�Ɠ�!���U�+�!�-�M)�;Ћ���;�+�\Z��5����A������%9�?��p�����4C� ��
Y�,^u/��;��V{	�8X�Q��=F��W����p�Z�^�ޞ�Y^ ) +Y�HL���^č#Q׻�e�Í��t���2nt  �M.�cǎ��ڡ0�4�"�ΘX���u��q|��� OX�P*��^���v{�ӝ�7eF���<��{�^|Φ.��*�M]�Nh8��L��,tT�<��<·��-x�6G#i"L�b����Qɥ�妍i]ǜY�]�܁����bU���굫������ҿh��úB�K�҉����%ƕНW+�ՖjqZ��d��[eǎ{<NF���R-�e�Ҩ<���r��1��G�:<A���C`��  z 7"!݌�a���z|¬�M7�$�<��mr�W,���dSS3rn���>uF���2%s����RP��j�X����W6/^�
�}������eI��M��qyG�Z�=o﵍��Z����$#M��@�(�˚]h�k�
�����k�3����ns��G�@��[�۫2� �5�c��zV��[�2��T�<�Z�#�ֲ���
���`�^� ����l�0�`�kAA�g�6�L07��+wc�>)OI��BC �^��gB��\��}!��N76���e�+�@ؕϽ�w����,S������{g\�b*j
f���Pq<!Ըߴ�f�7���d�Z���.����7�/��/JR���菌ܨ:;'+W,�����g5m�n�V�z,�3��߬�˖�~�c9q��>�)*��3� �=�� ��!A�˄��@���ˮ�Joo�%S�O�˲��-k�;�+5Ś'N9װ�b�Ē��%��_�n�&۷o�\&kn��G�S0��ʫ�)�M�☉�N˟����Jڣ��W*�	c���V���7��k��,;����E����'A���҄D���Mm4�
L�����ݘ��R/��4����IX��c�&�k&�Y�;�T��y�|2�AQ`,�}���N>Ƿ�k����|k�P�w���'���I�k��֕�̮kTh\��\�T�8f�������@`�q���@��җ�Ƶ�M��kEdr�(�m1b����[�����L��M���o}KJ�9UP����|�F�8�O�G��0Z��c���t&-K��e�ΝR,�dbrZʵZ{62 z "�r#J(�����,��v�27;\�o����X��6�7��)�޷��^�z�%_�ˋ���-�O~�礻��Z��ٳGf�&m�5zX� �l%��X+�⬺�_�<*�ZQ~ᗞ����G�<;.Ǐ�������%W��5�罝a5���l�J��\�,iMCX~:Y[X jZ�T���^Z�y�%�b��N'�cM� �{B���l���M�5�&��X?P�Z̔�y8��{8�|�O^�k��h����MNvZ���w�˼B���Ƶ��`en�������+�HR��f�sn�����{V�0?l���$��V'~�ƺ�>|L~��v�	�CV�^��CN/^�
D�*W$��Qp�����Mټ�V�|e\�{�'�yP����	�_P@䆤���!w�H@ʁͮ��L.��M����\�s��m�h.�^�D�Z�f���MĥZ���!=�K&�&��r8l���WezzYnF:>ɒ�˥V-�~��1��M���,O�,����Z��� �������?x�~t/��Y�����.c�N�1s���鍀n$%��I%p�}Ҥ�u�e���s��K_����޹o�ܜ'�J���W����:P��{6��*����خmϊ��E���v�:�_���ӧ�c=$����jed����쳯�L�"S��23W�R7�)�NUkW>/gΞ�����lݺU��r����}J��_������+�}�23]�u�6HF-ytxCr��+�B$jc�m0�H�U =�� ��!i�Z�L2%]9P\v  )����$��F�]�r�!g�]47(2��ݎ�� ���O���d͆u�s�n��޻,�{f��|����Ȩ���8nKϫ�*���5�W_���t�d��=��/ɢ>��b�y����{:�4�QZ��en�Z�v���K�4�q���`�r'�o{pL�c�9�[[���9-{ �fX�αI�J��9@,ݳ��!���5�������&8mO��+5�h��)������? �v�����\�|�T
�s���X��zP<b �����+Wʊ՛���J(ڒ.�sϽ�Q��2�%��G���ey�'��������o����XR#捱9'�5�iB�,}<S�Tښ���KT����lC���9K "�rC�I$[a	u6������C�Y����SO_6�r��1g����|ONƧ�e�P��n��
�g�]��֮���~H��g�IY�d�ter�� �dF��� ���!�j�`ԯ�z�q�(���f�w_����G���x63ȩ �-)��a�G�
�k�Ę�m��c�cӺ���� <�ms��x��d��ǚ���_^fY�
���B�bֵ̚����+���!�]����$7R�
k��Y�9
�'����NǇ
I&Ҧ0!1͟�N$�	/Fԍa��J�z�ócme��ԂK�Z1&Cx��;j�~��IX�HzO�?n4��JQ����UI$ch~.SS��<m����>!�\�)8����Zy�\�~�ȑ �=�� ��1э�ZS+��8�]}q�6I��!��slt��g�Gy�!��mF�l��;v�{w�h��)��%Ṑ����W���d;0w!��d<e.�Ҝc ���R�e��C�Z�.�5�;��	�>8��	��l��E`' ���=xz[�0�qg$��	^t�C`Aܘ��O�[�$�����Gv�����ieS��F��)pq=��2~N.v��~�<=��>��D{Ν�Dyd,�0=Ҙw���mU�V��k����|���ԅ�G�o��O��rd�r��QS���VW�d�R;����y�*Cc
�a9y�\�4*��K�d�a@�d�xQ��� ��H(T�'=�� ��	UJ���hQ`GF�a�n���{O���Z��*R*��
y�q=vb�'7ܓ錁4ܝZl��l�"K<��^x�UZu�����KV�w=z��m+�~-쑣GN�~jnY4�Al?�t�qK��qG3��O�J!(S 0HDù /�yY�F+�Ie��v&��"z�����!L�q�>�����O% �\��	�d��x�� �	[~���}�u�x=�m֯��~πt�[k�j��Oy�������Ð�?��c��2��|��tA�n������jX�h'�u�'��<���P�M���۶�鑳z?I��r��)yg�^�:!�xҔ�|~�LM^�����m�����Ľ�y�w�B�Z��ͮ\�
���@D@�E7�h<͖Jsw3, Q�Sӟ�ZБZ[ʥ�̖x�U�_��]R�%X�T)X�n�ܼy��<qBΫ%�������:26\4y�wd����~,�����lp��墠�0�c��-s��=����TU)w��B : $�x�4�Ԧ��F��&���% �]স�\Ҵr;�\=뗠B�9 �-u��<	� P�=��L~�R���úy�۟R�1�>o�d�#�,�3��U(����?��*2�eg};�
��;D�����i�ܑ	B���$RU��],��B8"�\��
�U����:�:�\��2Ni�Y6o�f	�}�������^�{�q�g_��G�������k��hCu�*�G��o�;�%n�B��H $�rݢuJ����~�6WfN&���𑣶9�&�V�J`Uk�1E+*�͕�ZrXͳs�d�Gy�J�V�[c���/�,o��g�06�F�f�K�Б#�b�,]l�h���?+��)�oK2��Ř��<dt�訆�%4׀�*b��F���'�	�c�l������U'���vfB{����Bi���O:�1�mM���t���	!���]�֝�	dh����E���0����b��+WL����(�S2��J
y�I{�W�Y� Q�ÄJ�?	x�y����p���n����'.I.�+�>�aXak���[�f]�=�~���9I�X!}=������K/�D2�ݒ��<f欳x�3�2j�Wt�Uٳg��^�T�H��XF;�.�<g��r��q��׾.}�P.K�v�|���H �,���u���pR7����/����x�X�s�.8���X�P��R�ძM4�6W`Ŋ���d��ҕ�Ys�tcQ��7����1˵���c�'��/|�jWe�p�Y��sR��Z��F��^�x�m�(p��K�s�ò��FL�uQs�v��&�A����B���G}�w�7����L����aZ���[��]ی�CY0�#����fn��毯qM�G���G5k ��lK�,�����{����LuT,����qY����X��{>컃��^_=;���^�(gϝ�e+V��U���'`�͖���J���� �V7���蕗_�W^yU���%�]85l<+V��z�j�	��r�ʌ�d�^�V�cQE�-Zb-W���g���Ĕ�X�R�,[V�����$�@H@�e`��vq�B=��.������Y��y+;��v�w$�%����ų���w��I�~,�C�)�ŋ獄���'O9�pl��ܺE���o�q���?&�HM��q�|���ܤې��ۧu�W�PK\ˬ: �mZ��g�p��%Z������2'�]�ן�g�&&$��!��v��)~	W(?Ph�J< q�[�҂gR�f$~�dͲ�Zu4��B�F8T:���F��\J ��ֆ�w�7���|'�<�6|���1q��S@�xԭg3��X��G�|H��e����e��we���>��'de�%=?b��P/��������>�=�n��W,l�Օ7v���]����T�!9y���:="=}�z��3W�nqb���Y�S��j��rOO.h�ȂI �\�lܸ��z��c��������n�`����-j��ikl���a\X芮�!�: ���h2j@4=S0p/��u`f��e�֔�\�%5�u���X{z�2;}�6�}胲f��<xD���3R��N\�uز~렁e�5~���G�LFR� A�����g�ӍN��ߘ���R/&~1I׶v�^"]��d4ƞI��o��X7掵#�2���j��L�w�e29�9�Z�ʬp��M7�dǃK>�3���@~���.�9�#�cx؁���0g��h[������N��ݮǾGO�x�>U���fd׮]v��K����a}.ڲt�?�i%�h7��"�͸v���Ti@��fOy$����z#d������i������_�'R��ߡ���WM	d�$ �@n@��=�|�Ѭ���%us$1��ql�
B���m۲Neјsz[yW�%�՛`ө��L�yW6��W cc�d� rY�U����o��@�?}H����N>��}�Ld,���R���0�m���.Ѹ��B����b>P �	����uZ�.A*g��3�����{u�dkc�PaM�� ��8����� <b��.�50w @��q/`:�yȴ��m��==v�^������J�1O$b|��#�w�^���;��Iu p]/��{�O���DB4�Pc�'���1(l�:6v��m_����c�0G�t �֬ ��<Y?z/Y0ߝ�9v������<W�U[��~���)�Vi�8$����)wͺ��LI2�-]��۬�Z˱��Ui�e,�3�sJ�rj��Ԋ�gA����q�-�Ta�E3����I �\�\�x"}�ԩX7�x�k.�=P�F8g��1�!o5:�*:b��
�H	K����d�d,n�¨!��s4b�C��A�Z�VU6�ʢZ.��{�n�RmV&�/v��},��M �b��ə���p? R�(���5�g�8 �p�{<��3�� ��d�10/��a��� �p��@ɸ4:�a���( %������xw�y���dp�Dǡc���+W��� �x���߶y�g߾}66�w����5"�����o�`=ùf,�}a�p>k�Q�����1�kb9>��%���Z���DG{�Z������A8�n��  ��\E.�\�w���� �2W*���fC��<.5뉎�'�~���#�
YXTp�==U�$>pėJe�/!����A��*��p���u5�,���u˹s#Y�l2 ߸nn%l���Y$!�xf����ǣ�)�!ȩ�B\��'�B��Z�n���M-��s� Ĵ5�X�l�\<F��q�DI�8{�%���L�޲,w@��rw��P(fqZ�R��۾V���h�1==i�4��`���?��Y�u�P8`�www)8��2&ē��:�$�J]���]��Ӯ`�/͕���F�cd'�u��x���R��1�(��)�;�j(� ���~��	ٹs����o��в�r4��7l���O�ִ>�X 8���u�"��-��v-r��.�����IqH"`�\(ǎ픎�U�yb|(P`�t�s�}����/(�G�@���r1�sg.I>�չ;�ZW�60��Rv��0ȁ!U���ͪwt��k#4���x�c��dUq��+�l�Ue�����+juW����{hV�(%���
lY�S˧@�#rt�{�{�yX�k���WoRc$�� ��nQk)��S�66��Y$	��8˹m�rc+W%�-3��+�r�p���}m$���d��v�U��m�.!���:}���X�j �eKMQ�4rN⺹'uXm�Zs^����A��7q|�r����X�e�~/q+�e�E��`8�1&6u��I�q R,cc��J�� x R|���pGC�����a����D;\���P$p_PDz�! 
@����`��q����N�~�r�x�2�y<K�`�3s�sa|���pX� �T&ic�f�a�f�X�g|�!�$ r]�t�ul���hl�Q�e�O�?���[z~�8273� �3k:Wqyx2����̸Ta��u��yG�
�mbbJuw<�S^|�Y���仩�+��k�T�;�8}s��*F��H�q�Q��@Y 	 =���t��T*^lVebr\&��S9����ݭ�
�	#p!{�lqN�j� F:11��j)I�%��SI뺆%pk'�	�� �;���C�3��X>�����X�~��2��[�X|��cACB��xv�u)	A
�y�f�T?Ʃa�> �� �$)!��7�h9.����_�Z���c����)��q�bZ���]�ܗ����:�*�5yq�73�-�R�^��*Ir����9�ea|����"��(\���~�F��5���t��nq 7 �c]`��PlȜ�o��z�B��9��"�+��,�0��ón>���P��ʰ.�r�T�J��)]��P��{ǽ��[�n��yɀ��s-�=	fh�'s�Λ7�bkQ)��̙�239!w�u�>t�'��������5+l��#W����d�MuV���v�2���` z �-�����mg��
O{=��d���V�ˀ�kZ6��EX<�l��Nh��n���MNy�t%��m7��Z^���%Y���u@�8�\�g����ޑd�%�xK���k��XU�z͖%�E<�`Cf��.h�6� �c�ԅ���� ]�:~MkPX� w�FM{�kx �l<����������j Tzp,�hc=!�Ƨb���⺸R���h]c\�O��#��`�����(:d����~X� %�ω����!,��l���X�渞��<����e��s��iP��7��|��W���G?�
A��9��X[���@��np�.���6d��p�8u��n�LZ>��O[ܾ=���s�R�L���7��;v��@�*~��8�NϠ��M˳Ͻ"g�/Z餮m���SY0	 =��[n�>^�9v����a��3��:Y�n���eK�e���S���g��+����j�a/]�B7Ҷ�� +VW<��V�N)x�<R2������ZZ��%�:�t%�����l"�kzp�C�-aCG� 9|���]����@��L�93�]ɕHWW�8�!T\Mu�C�j�ݨ�`��9횜 @���!�d0XǬ��ۜ$4<�sc���bﱔ®m,�㹬��u���tHa/��`�2� �����?�n��;���+��{���V��j�s�Oz��:�?�j�zM&�+���8 o����Z�V6n�"{�~F:��6|朼��ٱ�~ٺ�V�Pa�_,��W��~Y��6���|��Ƈ�כ����Z�Ǣ�����}V�_8-s3�2пL���Fi�jGdp(/���j��O_���x섍p8 z &�r�244T�8}**�LRڡ^ku�b�2Y�a�.R@_n�f(}�����:�K���i�h��Oʡ�G�^P�x�$����ǭ�ŗ~bV;Z]|�ֆ�����D�Y�f�1ε�3f�ێ��˵���b�ՎՈ� ` k��ᮆ[`�"; 	1s����醕뱆���wT�F\�V,^g��N�;�h�����5�x�����`��Ď׆�=��ٹ�j�$7~֡��]�7��*��&�a����� T��ٌ��z�]�x	o��\���R,V�dɈ[�V��sK��9J������|G�茗�IA�\YH��?�яX~ �5��^}>��>����zT*e9t쐼������Y�EC���6�O_zQz�{��|H��)�pnR���d	�PT��;�ܮ��1}�.��x�rd�$ �@�[t�O��L��N���Euc\���-2�x����K|����ɶl�jq���.Z=1b�5/�	<6td�ߴq��ڽS����RR�����e�u,9�FaŧR	�+8]�<*����?�a�4Jr�¨��o�G��Y��<��%�K�q���N�{@Ʋ4v#�)�\�~O$B�)�q���=+�Խ�[�ڮ���KNc�0�KzW '�A����1G(��م)��5������7�����0>���V8���&t�s\�'������
����r��mx�3&&=�:�p�[�P����DZW�v(T��s��}�vi5u�H�rFu�0.������� ����<����>=�۔Zܡ�E=?,������lU-�?���`�#�y�Ǥ��C�A9e[�K�Y��^����.�u�Mr��H4$��p z �-cc#='N��FP@���U˥+�gnb�V��$��� {d3���=]��cǏ���JR7dl�=�}��������>�8���;f�3>���|Dz{�2S��g�yF>����cPRD~ts��[>�m�� AluҘ'{w3k�y�� #h�Ӗ�wW#w8��G�4�g?u(  k^��2�*$~^t��A	�O�=	���f|Bk��8~c^8���h��}��G�6�-��S��������f�k��hv�	��P@�̀�

�
�p	�;��xM�\2�%��w����Z('�����W����/-�r�����q�l���<����:tH>��#���~V~�3��?�O�I�x�e٢
'J��w�t���jO��Ы����W%�EW7]�\Jڍ��(��33���I �\����%k�Zʲ���4���O�W�j�ܾ�N�8э-�����e���/yQ )�D�[����^��g�e�-�e��=r��!��c�4rnXĔ�wW����G�|_�{�{G�+p�תu��%�p]�ב������SB$�ML��K<�k�Z*K"3k2�θ�����������wgR�sfF=A�nhr��}M���@`'�,���H�B�X�m��n�M�T6�A<��%(B"����=�A���ϰ���n�Ƽh�۽�g��#�c1���JG������WJH�=~�\(��t�,�G$��J�&ɌKP̴Br�w��F_�4Zu	�5�P����7���lܗ_zA{�ay�]����4��hJ�7�$�����㦀.�M�6��1����K,��[�z &�r݂��l��n�q#�@�o��icJF.]��j��1L˰n;�2� 0�}iw����O~�Iټ�9|�e]��֛�yP��2	��@lC+%f����@k6iY�X�ŎA͉x��V�Y	�ȋ��k~+� `b�V�T�u,V6�|�+��s�<��MR ̂'�+���"f�~H�J+��Qix�9c�8�B'C1"H�����L���6X�ZP����?a͟���#��A�c��s�r`����~W{��/(�Oy�{k�,yS
J:�T���V��ho�C�dL(b�<���w\�;v쐷�z����/#�=�ݼW�P�$�ٙ�]�w�ޣ�="��=��7��:���27[oU*� �ȂI �\���]չ�R5	YF���+2vuB��u������ʩ����o�&���g`4v媵1-Ѭ���s��=���e݆�FGZ�+X�t�k��d6f���.u��u���Pp�[Ʊ�wܵufX��y������N� x�jua3�;x�J�ܨ��� P�G��\��َ��@��V4���.i�t����v{u�a��"&�q�0���	�ժƔj��lLMMwJ��f�	�<��B�z�֟�tf�3��@��Ѝ�D>�,=���,�q}79f�3���<U���N�׋�"F�~n��bE�}I��4����9@���I�n��x'D�I�e�=w˧~�gT�k�3���U�;��.#gϪBАt&+c�S�W%���˺H��*�O�G��+�8��	)L�HN����\C�L �,���u˚��S�l�z�ȑ���e�d���	9y�e��|��ec3{��'����r�d@V�7a#������/�(����EX� ������	@/�Z�hw�w���L1E�ɒv��$�1���86�pM�@IU (��N:�3��qM6���H ���x�T����,�d-��u��uZ��|���
X;����Er�f�20���M�6��@B�>K� ^8kˤ�ŋ�ll��u���Ӂs0 7k�Y��$rSy�9���b�_���i���#T��~e��#d4��{���\.R���$Pâa
B?�r�*��!D>##-�������w�� =)�:�	!��<~X��-�l��~샦��&%K�|�	���M��j�b� �Y0	 =����`���oT��m�HWk]A�nh%��M\ڰT��k�(��$��[W��Z�i1T ʇ :p�c������Ԅ,ZX�,�Z�e�d�9y晧;�@�^����N��*����u˴��女'^�_��\� p s������@?k�{�36 ���Sp]d8��(�x�{h|�A�j�s��Y� ga�c� U$e���h�.bf��ݍ��lx:�l�b��1�Q��ZC��w��Ļ�k����/�y@9@i���3���߽���zsZ�,9�1%����+rMN ��5��w`ߴ�7� 2��?�V���)$l�6vRj͒�'����S�WFj���I�K֟ ���*��~~�ay���ezr�>ǳ���{���q�r��������f��1���U����K9=|D�d�X������/ �rR�MM��"�0tg��X<)g�8�w8�,`X� K�g�Z�T�u�+�Z�ZE���a�Fs�Y�H��80�A��ܳ�C
�5ːA��^p�|o�����t�i�� B��7��ޞ'jq<���MA�-� o 1��Lq�I�Z�����j����4�P�`f9�C( ɫW/v�d &;�AQ��ǚ����ze�>�0��˖�i����X3zC��H�:ָC�H���*�����=�����5![�����z��A���w�L����^�Kj�˝?�/Q����7B�Y������y��	Y4�\r�^>s���l��j^y��Չq`x|z�����D�)4ᱜ�\���g�b�9U��?�g'"�ʬ>tJn۶Y�j��ߒ���;T)������ޓ_|Ir]ݺ�N�C �,���u�ٳ9�ޢ���K�D��ȥ+
 �$�rɎ([?�pL2�Y�)��J���*���믿.1��j}>���f5V+e;r"��:�m���B���F��f\�zL؀���%sybo�"�R�yв3+��\��L� i0��@���ذ|���c�8�IW����zZ�H�B9�z?p�33O���u*� �ġP�=0��p��v�ڇ�vw>�k�u�8������ȅ��PV ���AY�8*ޢ zP�c<\nv�-�`sܫ?��9�ԧۛ?t�3߀.w��X�^��>�f<_C:���BjE�M�[?r^��M}ޒ���jbvvN���LN���ԬT�g
s�~�=2g�e=�;��v��c'Ny5����>iá�
li�)�gd��>U�e��9z䄌^�Q�?0:zY-��=���Ҵ�Ѡ}j '�r�2>>��|�R²���q[\�V�Ѡbs���9 �\,�1�DJ]A ����?3+�����82�!�i��hHbu�^�3]ΰh��Ǐ����{v�!���W����o��C�27]� "��2N0Ľ��(�`IP;v�X���&^�QXڈ�C�ׄ�N:�U`��C�v��h��x���%llH~��W�s���J� ����}�(^X���qk�q���d�o��a��P��	ڬ]g;��[���h�Ӻ��h�Ǳ�˵�m]g�����8���m�!:H���7�r��ҕ햁�k`��+��Ɏ�hd=P�9Em�׿�5=~���|V�^��Z3����N�g9��K�ҔH<'�G&�̅Q	GZ��X�;A�}J"Ś>�����{ &�r݂ͩ\��Dcm���k-�[�����Xn�m���M?�0�W�$+O�N�z�aQ
rI��XK�[w���]ͱ����ҕ�KW�d߻�����B�,_��6�������+��YT�C,!O�	o��찣!�,���JΊ���`	CG�9��َ�aL�j�Ξ$1"q����A�!�;���;��(�C��f�,��Y�%�tw��5\Ӑ�)��񃃋�7��/��@�,U?˚����X5�蘝N�4��1�� ��i�3s�ʀ�h�!�d����sn�!��)s�ԴܵB�%nc�t�c��0z���<8��q���ǑL�䓟�Y��(H42�з��s�^��Q��T�m����e�e��,s<;|N����ӕ�+�t.u�����j�l��U��0�8��	��Rm5�<[�L_�D�Qi���r��@Y 	 =��T*�T˹�2�����BqI�Q*��ȓ�z�;�G/ti��s�[HDa��C�T����P"f%YjT��0����䴬_��xCr
��!K���/�H����J�����6�Utq�$V���������i�iX�pSC�@�z�0kq}��a�Ê��
��t�\� =X���C1������8�)y�q����6w7 �F� ���K������1y��G\|�H�ù�"�ݏk��s��O���a��v��o,Qc�8Z�.3�	��k���5�:y���%��(��9���AE�ʂ��V��!��N[�A���XStSK$��GV*|���W%��ސ������4ȍUP�xn�&��ң�ԣ?(o��WFF/˹3�e��e�d�bWb����O ��[A�O����)v�.W@�e�A=��� ��n�+dә�3�ې�%���[���0���A�R�V��!�]A�"�qs�[Fb$(	�Y�l�UK�Æ�k��%�)�~��������j�}d(�v�H` "�.k���u�<��F< ��qmX��֭7����5���NgtN��-
f9$
��jj����˗�0P�XP$�~��s��0Zl.v(���!Ο���zK>�я�� "ң��`�u�8d�� �˚arĳ8�m��p�N%�d5]*M$�a3�����ą��p!�qI���ԍy^�h'ގ�J̑�X�D:�&��>�m�x�1�9"����w���qryV-�[o���}zF������fe�@�*F�V�V/�t̂ıf�\�T��d3��Ǥ�ϾuDS�xJ�d�4]
\�,���u˪U�CCo�[۳t(��֒�J���`fk4�
�a#4�4A�Ym8K=���Ujã:���:g�����j����`���йb��X��gE��ڵKe��9sQ�ˎR��%M���p͆�ݑ� ����> a�l�v Q�	b(Cb^�a3����X�, �7�E�Y��mYq��v��A���	nP�m�fc�w�%��~��z~��Ap> ��8�F`I�3�[�BW7�#�,^�~�Z���O��԰�^c\*��%�,��pϜ7߷�'^���Um�{���)}�F���|Ýf�8󅇌P�5�NX�j�B��ǽ�U��~��P�,��[/�}��M�+���┈����Դ=U��jW�^��r�(�TZ>.}�CU�4W�T"ֹ.�@L@�F���\�Y7�J]-K�x�Y��N�PS��Z�V1f�E��9��`F7�dJ&\?��iG��wX^��ŦH7�e[7�yV�ɢ&1�Q"eԜ�p¨_C���9��n�F�ա^P� � DXd �T2�VڔY��B'���3g->����%-YԌǣV�����$�5pA�9;��X�M���d��|0Ƃ۟V0��p})�  �7�� � 7�ZБ�0f��p,�	/��Q���b�T�འ��·K�|�(�üp,� ��b�,a� �qM�ƽ��V�tz�3�Ŋ����z�K �Y]�����&պ�7(�/
J����z�����;%$@�jAff�d��.Y�t��]E*��SɈ�]5d�OM�u�2��Ų����A� T2 �@L@�e���̙3�7��x5\��rU�8aV9�t�	E�1-��率 ��ug]�3sŶ���$�T�c=ڹ"-3�ŵg�OZ��-
H|�ǒ��2��B�$��� Z�֙܅���HԕL�oқ21�L�0�ﱏ�e;{.j2��"�B��v&ޱ-*y�8��3� p�{�����hU�=&��7��:�o��1&N��QX�TzX����!�����(c����p�
���sp_�t����4�?G3���\���ʁp,n��=g>��17kL�J"�0�"��vr0z���亐����KT�k��E]���Ւ��-��/R�7/��.U W�m[7�E��l.-�RM��s@�y�e9�����n�z�jU*��` z �-�/g���tetS�d�R���[VPK%����mgmSW96p�� ���v#[�Y� �Jq�ڎ�zn#1N��z��)��x�3Ê�cl�}O��W~"1�?km˺w]RCF�	q����V7�d�g�QK`�`l�=��I�g��f�!9������~ǹ�r�^&=�pd�
/{�\ ���G�}f��� �X4���)�Y\�Dx=RŒ˝�e�/ۭ���4��qm�� i�㇄289t��x@Z�$B��u��bIjz߈W3D@>u��P�@����x|4�x
�~�f����b֫w��.�ԩaU.�w�݊�ő��Ziʺk;�s~6�1e+����*�1�&1������>�W�~�M)*r���w���e��2W�����+����G�=w�+?����/�O�xʊ�kC�H+ �@L@亥X,ER�T�O-�3�����Us��]�F/Yj�EK̚8�J�zu\���!���`�%y����*��D)�,n$v<<���+_1淙�q�t�*3֣��j4Z�N��t-��v��ؼ����� ׂbB>�|w���� p��e�Cخ���z�� l���I (A��`��2���{ B ��+����x n�nn��`=ΰ���lr·�K���'I�θ.�N��f��i��H�q{(P �*���k���/( ��c0�c1���rd�����7���μ+>܉�SP!p��)k���?xV
�eY�t�)��0i��-��&�W��;��j��'�Mo�_��_�W^���Z��ͽ�,��{�ҫ5d�8#7o�lI����<�l�֭����s��/�O��[1� �=�� ��n�����C!���+����e���f�z��7޼I��Y���g�����W_W�*Z��R�V�~�ӿ(?��Oe��jo�e
d�=���s�}G�5+�5���P���;V6�f�r�V��rAP�;6;�5f�')�y��ě�t��ʾ}���u��H�;o`�>W�b�l�t��i+/���! �!��X��'u,�������J���� jK�	 ����1�:��б�8K��v��gxc( �q=~���^8s4?/	k��r8Ix���S{�1�=�����{B9����k�ho:,�E�҅�����{��{���JM\�%����j�3`�[���c'U����qU̦�
O�<�29�$���y��`Ǯ��k��3�0y��q�o��Mij4aɗ������uڳo�l��Vy����#�dj|Bn�i�}��JQ�]	]��Ѓ;��3iߝ�@Y 	 =��d2Wi5�eP��*���ˊ��t3]-�LZAzE�ɉ��k�����c��o�����+[�_�.�jv��9y��~Av���3XT 0��hd5���XԬpl�O��GeŢ^9q|X~�w�oa/?5�<��s=c��$����LciΧeɱ�4-r ��`�� �8�bp/�غ�]��� �c�N[ ���*
��c�Q',s����p���>�_����c�s1uf�3V�1�;3��:������gd�cf>��4�9`ݙ��>�s� Y�2��<P�`i����K�<��t�������"U��\�=Kg�^T ��ҥ�e�h`�dHׯ�p�fl̰Kĵ�z��җ�$�/]U��s����'+���ŪX�����T�|/��$��o1V\��0nH5�Y�����[oEB�pL	d�$ �@�[6o^_z����sgOo���;���H���8��
�u�6��c�N�Z��N?%W���˳f���[2W(ɺ�N�=#���f�<�v��L���|�R����e���e߁��{��y�c�d)W��r�6��wm6��0�u��cΈk �\9�W�̚m��K�kرN)q	j̜F�z�r��-�^"[��o���s�#�@�Чk�����Z:\X� if��}�����z�{t�t�3[>�ՅC���Ħ,C��叐 �
P! �����A�2���Rgm|�����kal�&h���7�+w5��R��F�$��d^��?��P�^���?��*UѺ��vmr��Y9��Ay��7�g~$]����_��#W��g��w�yۈ�Ο9��MFVߴ�y �1����a�V>%��yX�'�,K��tue�:ל�I �\�tw�j,Z6u��C2>6�I�\�i�袑���~��t3����N6�\WFƧƍ;�Jv�@Ak
�`�X+�����P�cA�S;�r��x@֬^&c�#2v��Z��L^l�5� ���5-8)���5Ҙ��0f�ڷ��ڴ��=Ƒ�p |Yo�D9r��5�Ef=�ǵ��ǲ3�Ł�l��q��Y�նz�T�o���k��O��oMJ7<=M�Z��`,̃.��G��$��K���X�[�n�����
gy�sp?h$���]�䈂'c�䋷�i�\�l@X�Fk��[��H�?��6<���T)��� ���GZ�N�/xA���$4<�����/�?����o�������쏟U@�#�Z�ƭ�j&����{q���v/��Y�|H"H����rrj��g�=�츮3�]7�{;7�F	�"	0��)*��$K�xl�=~���qX�Z~kٖ���g��ئdi$R��D��)f� H� rn4�������>�oZ�������Ս{�N�:U<ߎߞ^L�xr��tO޳���;;2� Wv�Ҥ��>t����z���j�&�	��x4F��,��E���KƄ8Fˡf�9ڵ�-*�X�����&;�a���>'n�-��ժ� @�7��p��kf��5��,��[��+���غ��5�]�n]#�V�&S��F-w�8���!�Na8O���A|�st^R>�x`�i)�
����Ph�M٪��~��l��]!�d��k�1�th闞��1w!�a�Ԅ5\��y��/O= VX���h�^��F�5��Њ�_�@�A%�G�?��XV�4b��Xh��Y;�UuZ�B)�V��ޭX�����]TA�!�'�ꪫ��믧����I�Γ	jT����(��q,�)���mx�1(��ȱ��E]���ӳ�2�<��<�螼wA��l�59�cp��d��Ό
�$3tz�-[��������ر�6m�(�Y�^�T:ƖS��������MW���f#��z�$e�z����k�5����~_@�t$dcF����kif:'@�ۇ�S���T sӭ�-C�lD]�ڍL�M��n���vkC	���5��s��,�Q Q*U�i�jǾUI��y0��q����j�.-�R �)�q Xmo���>t�B��X���#[�����$:@�#_�.���0 =� ��ڹ��|��&XGx*�4��ֺ��£
�oB!�v�d<j���RIV���?WXټ�A+,�[�>�rQr>���K��'��z�z����r�f���L�N=Fo��:m����|/Y�J@�2��H"dn���0�y!�ȱ�۟|�I��s�'�Y<@��=K�5�D����ѩ[㱔�d4�$�1z��+��zg���ٙ�+�QWo��GOS���NjT7�'p���޷hF�.Z�����e����[ǥSm�I��t�ƍ�qf��:i͸a��X�����pw���u���n@�� U7�r�kM7,=��q�:{��v\�
��$�l���d�MO��E�x-'S�VU�c�ծ��ʃ���[�qf�B�� SF�T%[Qw�\&yK�T�?P� �x��
�%8� x���Pv�P�����<�E��"���j�� u�����ܺ���y�dZ�<B�}��s~���������K����QZ�fmy�%���G��W_I�V�.�H8�VRR�$�LM��i+�O W��b�Y�X<,��
����8LKV���l���42)=@�伋�,D�W����i��	?,�]���ͽC������a�F��蠴�P���o�Ca˔�'$IQ:;��]��x�����}�Du��mtv�t<����"KHL�3��fز{c����IQ�Wo���4mc����a�]��Uk���[mF4�q�P���PD�:Pjr���od5yc�gJ�b�^jg��+]��&V_m+[V�ܝ��K0w�mc���(]�ޏ��+Q��� ��)��! �€{("��Aܿ��	�-_. �,~��q.J�&�)�-,p(�k�����u���1.>�:+e�&���/Q���
`�A�>���k�40�^z�+E�D�b���a�S��٩i�^N��9@�|�)Z�|%�[��~��Z��"~{Bt���T<N��<e:;�����/�h���E>44H�:�9[����I���w$�p��O�B��'D<@�d!Ҋ%c9�g7+(�1qXbl�����[4;��x+ܬ�#g�M�P0�MN C<H�J�^|���������geC~��?���'h,����^�Ϲ��	 j��{�9�@��o�[tf�-6�V�l��Z�l�g䓤�&Z�������f�e]
2�"�����pS���䬹�5Z���n��/Y+D�R����r�2�i
 ��ĈkN	��-��ӆT��j�k.����a9�k7�,X #\���t��i|[�S/�z ��z@vІh�@�>��Hr�o�I[�n��"Ԯ33Yڽ��v��6�z($I�JA������4��C ��de�Z�����h��7���ҽ�vҎg_�Q~�P�����9~��i�+qGIMHHj^x�9*�<~��������4Y�SB�]�G�N��s��;����:z��؂������/�Y>��o�!Q
E�V�+]�䂈�,Hlˮ7햍R,��R�"�α9��%j�pHX�J����߅]c�Ȥ� (�z�7yX|C�Oѣ?z��A?=��W��I1O����*��
������G᱊�IF�j4:=C�X\2�� o3j�Hn"�4��k�c���Y��vѫ%��[c��Lp��ͯ��w�����q�Wk[����������V�ޏ֨+@]-_X�8O���ư���Ni1�[��^����HT������0��(q(k�J�It��@V:�͆w7o	�s�����~�~�Z�L=]��g�J�)��u���r����o��:����K#?>x��<,�h8&�yA�P�?$���ό����b _��O�Y~M�b3t�,{������K�K46q̪�k[�'D<@�dAbY���Ƃȏ�RF��8o�	ʱ���2o�
GRizjV6LI c���;ʖ|!�5��Ѱ��Z�:k7��8���]�k�� �t���M���S�?��M�>��*z��f�s7hB�S��e>a���!
p����!�!9��^��d���y`^Μ|.�»]�M��[��;�Õ�`�86��-g<\.r���:�^��G�:��c����_`㹼�����V��NXI�c@����O�<)nz-8#6����4�@��Q�B���k��-�/�s����+Vс��Ҟ�T]�A�'r�x�0gi��V�-��L�'�1'Ϣ�xhX��wn�R�N�3�دP�g��A��D_ B�/[*5ff�v`<���螼gA��/~����mi~b�-9��-�I���?�{<������H���2��EbQ
��4�5L]�`��b�,/Kf:\�J�����;�ŋz(7�ы7n�[Kb�ھs@�����{j�����Yz�������3��Z���luek��]ƥ%m�d8���s��Z��r��J�GRO���i�*	���1r *�l������ x���U���QW>��x� ���: NT9���2^���G�xd�����B ��B�%sZ[��z�6u�7`��z�������?��?��ق�,`n_���4xzHH~�s�;�7��L)%y�-}�l<�=BRԒ��܍ [�>��F�+�_����a�!2
	�l��l�=ݓ"�{� ፶:6lX��|�_~ИmT�yJ�['B�).d��`������~�wM,� Xy�Գ3S�J�*._�j'��st����@oZG�?����uwt
��.8��nQ�Sw�[��nP��A}�����D�7|t�oU��k,{�K^�кru��ziݺ��v��w CmO�� ����u���#�.e���z 0��q�ޝ��+^s"�M��pM�Nk�,?~T\��RJ��_\�Q����?<d��q���^
!�-���%p��hzf����@���H( rC!%Bu��	�f]�#]Y�q<�B�W
[�Q��a�kٖ��ū	���-�ϳ�=�0��'�&�ܦ9��Z`l�؜5+���U���ё�p$H�l��XWc�^;sIu�����~�H�*yc�J2[(d�˰�k�@.����ѹejnZ�SAq~�����2?��nV����3-�k�����:�f�k�7Ɋ�����w�����z}����4��@��
����RB��9�1�0��%p��X�;�k\������T��`�P���V���)u��tp �Ѩ͔;��j�Ůk����IƩ�@�q5!�P:-a�<#h{MR�L�/ �O�z�zMMN��1>Gk���8��y�@TC����-�鲓��)����L�=�+x��!+4�1�'�E<@�dA��x�j�Z$ �}��qq7e�E�v<�z��Q��VZj��~q�bS�K����F&2>K8�Ô�E�Ȥ�x� #�/��4�a�9Ǫ~��67Xji����;�>�>Lw�N�s��ݞw�:�Q�cw����Z��DE����2h)��(�d*nf6X� `XŚ������+ ~����������67;��/LD/|?Hr�g8n`�b��>�n��]�L�|�>�9���3�N5D�3a��$��;<�+����b��]�e\�e��Յ�j�,���{B�sߴy��v��)�͉҂k�w�(&�`@�Ϧ�<"I1*9"͆�tH2�C+@�|'�r���'D<@�dAm��l��cy��j6�9rzf3hԪmr�c���GM�n��ʹS2ѕ�L,S>�$&�%{@$|�v�V��*��d�(⿆�~��u�k�����M�+�1��&��=��ֺ��T�r��|ݱw�@�w�\��tl��ݵ��r3 $DK�4�� 8���b$ʽ��K2�V9�&���ذ�U����׬�]o�!�1g 5@<8��;���Lr7o��{�����6TF�:������Np���j�Iwp��Os*�
4���._-�P&�4������(q��N���[��[t�]wR'�KȘ/�����~�|����ZB���V-K�a*����ӆu�������4x�9q���G�(y
M+$�=� ��'��y<�%3؆����Rl��$���I��fK�� `	p$��	�RkH-6��B!GQ��P�c�2�V@S0М:y\6ydc��6��YA2��n��r�[M\�(c�O��p���D(J��kFy\q��mk�MI�d/'v�����9 ;����PK�ݓ\Ig܊��(��x
�����@�1w<'X� k��{d��up,q�1B�Tq=|�s����vxX�������2ڡM.����=39!c�^�R���������؈d�/Z�D�0$�A)@U���k�TE#]s��ŵ���@�z�n�kMK/���>Ip�|f��2��4�D��x>���r��������M�λ��GJ�!��3�Ӗ���K���L�T[88J�|�Wx�(��h���O<� ��'�x<ҪV�v��vG����/���EdږZ���e�	�g���|����3�L�PD����C(�u� �F�"���x��Q{�J�u� {�n  Rt���O���*��3���4��<u�]���0&�Jk�!p-�g�P+\-}=���v����w��ݮx��^7'{�E6�&�q�H�q4Y���`4+])d�Zԭ��mM���,�Q����X��K.�ca��z�߰�q�s��0�C�,s���,���܋6�Ar*5�O��m����)��ߚ����N:68$���/�g],�N:�t�ڴ�`�s�E~��>���mt��J~ ]�)���w�F�_�~�v���9�����������	:|�(����{O<� ��'�V �A�l�[�n�-b�_|�&���h��,�7��E;w�2&�.}�����������䯞�n���s����˷����/��\*�������ϔ�N	�⨠���۵�מ�vS�*�*��Xn��/�tl�j"j��ֵ�������J@�>��J�5�n���#.ۚS8 2g�uN�����-��9α�J��`	67�"���r��v e<C��1Z��↫���_�9IJs����o �_�b�(�j��rP�?)�w��W&:��4)�x"��mO
�i5�BC|��з��99��;ߕ���B�V��lV�PF�g�c���/�?)�	%<P���h�Y��A�S���#�r6U)�/:��a>�t��7�Z�����Z��/��1�ē �{� ��X����I�36c�C��� �%l� ᨻ�G6jl��b��K��n��B����u{�>-IQ?���骫�!X�����(�RQJܔM�:59J~_�V-_��\M�|�ʼQ���$9���Ic��uus+�i���M��jV�Nͺ�Y�r��AQ�h'v���^4�O���G)W�w�<����qw�^�^���(�ntSm�a��9����S�U�]?�KZy�amk�9La�C������5���$9���c�Q�ߩ����e֫�l��0xV�X":<Dp��r���������L����	������kBu�5�=�q� ��tQ��Y�m��&�������r�*
�T�w5��Wl����'r�A�/B�xr�tO$ͦe�b	�R.�E�%�/��2'�da����u9ot}}��>�����}T��2�Z�)� !��-��n�Q�E�ʧw��7�Dbh��I��)I�
��}�#��tvс�G蝽"��R�}AL�9"c���N�s���+k{U��1�]�U��i�� :�WEb~�qxMzS����$3w��\�v?ʥs���;���h��=�#��(pko۶M�e��4�������n�:)/�� /��R�;�'�������hֳ��2.,}m�J��xW�$b-�J���A��R�t�8���(^�`4A��;��f
&���x�9K�K�R�-� �C�a���-^�'J2ܡd��<x^}}'Ba�����ݬ��V���'� #$3!$��;o���o�m�*�Y�\� ݓ	��͛��t�-,�^��a���e&u��A��z�7]l��v~��IL�e����'>NI���zX	8xX����yz�՝�jE�o���:-lt�X������^�����c�l���6���o͹���l2F�u��O 6rX�Ƞךw|p�Cm�v�6ĝ� �n��s%X:77hk�u�˵�V�gp���G=�?��U 0k�U�'�ns(L \�  5~c������3��� ��3�)�T2���o$���E��Z����7@��\�Ƅ ����޴
\����AA�u�9���D�>���l�\)IIٙS�ZX샧OJ5F.g*��PRP��1��q�]�?@,JS㔈�BE�jI����(egr�l�z�?�!����磍ǨQmy�'D<@�dA ݒ>�h���l�+V����O(��.��X:j�cRZ���# 6_�j�h�ǿ7l�DO>�K:p`o�1��C�S���K�J����C��`�U�jՔ�a�6Y�a�r'�0l���]˭������p��dV+@��.+#��.?S0~7:wBZ���e�����q���6?��NxS׽*&�k�RWo����# ��Lq 4X�8 �yxV�w�3r3�c �\?�0W�<{X� JɌwZ�$�Y�#V����0��W����q8�y��F.��9���v�
�s�r笯v��:�_���-]B;_��՚��E������ɽ}���{�����۴%�~����-�z+~��)����Y�H�{��4��;�7B������=Y�0����_HH��dGB�>���E���$e9��>�~���Q�3��Ɇ��w���oڐ����@��<4|F�F� 0*f��lg��+���c��=*;��sx�� A�V(
�JR㶘�-��o~���&�[t��	)���/����C���'�q'ٹ���V��Ν,�Ob���;��Ϸ��U�����{`��!+��c�8��aA+'��7���N@�A�T(_�4�P��o\����@��q�FQ��:'\�Rg���5����j�q2�a���T��wJ -���z՛���AJ���z��<�W_}5����>�)�õ�$u���e�tl�v�x��n��?No��K��T"I3��R*�Q��sKRY1<:&1�tG'=q��oHP�<W�7��*U���'D<@��=����ַ:*�b nXXgEPGG�e������,��3/��-��"�Z.[�Ǐ���s�Y�[o��n��6����/~���j�9���������H���xR�����iJc�a�H0AccTak��V6q+�.wX�)_k�w�`���m���l�ŝ/������Wi��Ẹ�d*����8=���R�T���lɼ���Q,HG�3=�s�7L�O����δ����c��?'�u���f��U�	rj�l�|��`��'$ʊr���k�;���l������Z�6�s�kY�]�6���z���=59�&��b��z��s�d�c��3]�2晑�4�ϵ=��*N�ĖB;h����,���N�]k
c�(<�k������f��낎����f�S��ﯽ�F��?�S��x�f�F'&���G���?I��_��������3;��8_��K��\�c[�"���y,��^_�B<gԫ�2Ѓ'��s�W���ݓ"�{��f���>l�ب<"�;�������UKG�C���ܹS\����e��� C9�2�"Xr`��x-8Ņ=�/�b���N	(tvfd\d8���BI����]��t���B��*Ę�3�l6+��HrxnP,�޻W,vMDS�h�;�)��͚�zu���Ǹ��̍!���N��n:��R����Ķ��6�:�r���C�\��C����s�=�V� �>�G�߰v5�ڈ��Zh���%#��W����R
����;��d�>�t[k�����D9Ͳ��&@�\������������ ��$v�g����o�SgF�+�?@�~�v��Ř��]o�G}�.ٺ�&�'�P� D�b��<�Wӓ��||�G��7e� �A�`Gg�(��H�\A}��_�R���gG1GϏ��޽�'��G� ݓ�e�P(b�"
�l�a��U��&��ϻ�{��ɢ�����J`�g�D��[o�I������*>s�֭]#���7wQ0`��9����Ա�ϖ���7CG���I�U������~w_���&a�EpF��ƤZꎗ�o����BW�v��g�S W��5�Z�q'����1�S��h�ݝ��m�����
� ��ƪ����	�)�@p�����T2���	<mc���&��<m���h8�F��.z�'�h���'�	<W�����p��s�q�6+n���r�oL��1�����￁�%�Ʀf@u$�?����K�xTB'?{���l�*�� ����?i��-�;A��鬸��	�dg��g�;T�6)M���+�c�N$)��*6���������V@���o�"G�xr�tO"v0i��M�X��P���J�{��x;q���o�#��H(��
8�׾}t-o����K�=�B!�o���ǎP"�R���F�$�g�B���Q�Zb��$[�l�U˒��r�� ��N*Ζe,M��֮kJn�=Å7�����2 �`�%S�x�����-[]�u���u�縭}�g�پ�{\�[]��c�Z��r�Zu�+�� ��p�� \�P ��|6���9�=~�x�BV;�m޲E��:��0���u�:B��kz��0����dh}9�7�X�x�|-$�5�)1����_�?���%�/KW����1���:�U���������\�x�&90F��s]q�V��?�"�o�%t��7S�X��_w=����_�Eb)�6ge1��Uc˽L�`���j�:��⧞z�^}�5!�i�[t��W���:���k����'��G� ݓ
[���w�ɜ6]��?����;l� ?l�)���^@�7d���L��2iz��')�����7H�,7l��4\��o��=�3�<C�b�.�h@���<�L�K,8 �Of� ��)�&c��z( ���Ԓ(��0���/�;vP�A��c�,��>�-_�����_"7�N�v��K���%�?i'ƹ��t7������n�����:��������L�|���<q�>t��9��Kd=�}��π��w�b�gi��J���?�u �"ܢ�t�K���H��+h�[u*B��ׅo9O�O����>Mo��� z�����ޖ��Ԭ����-_�\2�7�_/�ƽ����ᓧ�c��7$����~O޻P8�xl��41:I/����h�R.�p��#�u�կ~E�7mB\�s�{r��tO$V˶��(~�٨; ���� [ݰ��Qc���62�Tҭ�R�$3$�Nl��S�[��gw�n���-i����$:9nrX����Xt������tl���^�~bÎ7�,ӄD����X?���~��d���z��;����?}�c�R�}��]�Jc��vw:D�q��ݖ�|�w��A4���L�`�Tu'�Iy��.��Ѷܱ M�����o<?� �(A^+ܫz/����7b舍cU���c,e����rWo�"�GV<�,t��5����{(!���h�H2#+l�~�M��;S�LW�d���Ft�� �yZ�d@�_�z]w�5������Oҥ�7�~��;���w�}�������M��>6[�u$��R
oD_w������1`M���Aj���.�'/�~94,/�ݓ�.�{�a#�e�A����l��jW5�����l�(�1IP���C������*�+Eʠ�4��ykՊ$$������F�#�
%����Z�b	e�����j�R�z�!��\�o2i ��/nx���PwV�%6�v�3�䭿����|P,�0�Vڧ?�i|(%���ص�<L[[�*�i\!�.��� ?��:�Lg��۞�ߖ-k)����f��ۖ�Rq��XWԃ�r&̀�{��d�#+����4��F��C�#I�({`�[�IF��P��>��Z����YMr#�d8|v��W���~IT��嶲��FQ�T�v���>G�2�� ���K���ҫ��q�ѐ�5�9���
}��	��S�I.ބ��x���3�Ҙ����(��,�Z�D	���-j��
��{��U���B��O�ɯZ�<ݓ �{� �D����S�K]�C�����.�o� |&�)�ۖl�l� Dl���5c�a�Hl.�2�=�|����S?�A`\ʫ*ee�Uo N����F�v�/u�Ţ)��,�KΔ����4q;�,��n:��nw��OUw:������t���w���Z��&��z�@�TM��Ys�ו}͝,��r�%����7ԝ\��! }�v��$�����2G���� ���t 2��Ф��]�ַP�R����#�9p�c^X��}`�}��E1)ԫ���ڤ:~W~Vh��7lZ��V��0�Cq��{�r퇎��bb��w�d�c,$���1��g>C�R��}�Yz�?��G�����VX���5^*5$�29���\lr-�����V�.z$y��y�=Y�؍�r@�Pwz<a���@��mAqC�ŝ��	J���w����Ӽ�"��zP�j[s�������~�tU2�W6�v'1�,�f�Wʕ�;�1�6�: �2�^�������Lk�Q6��lY��\����6;��jw���q�c\w���V��x���t�%w��1n>?����owM�����8E�Bwz�O��ɘ(_�k�~�u�ёC�h|dT���*W��x��wg:C'k��%��(?��-����`�Ń ���1� ��l��I����v�x*I$�2��I�3~o�H&'@��}����
��PpM_�F��޷����R�T�c��l��{�K�Yr(�x�����w�BRoD��� K��>���d�C��ɞ'�\ � ݓIö�z�f�B1�q��ٲ7+�έ6Ũ6:P`��'�)c��'��xv�7C�F��z�ħ�}A�Y
���P�a,v���0�6aY~c֚��nKh��EC�ܥ�$������h|^u�c���/w��ɚ�,l��|��Pv4���v����ݠ���d4=G�Y��k�_���7֫ƭ+_�g�����q�����1��{N���`��$�L��n��fn$"�Dr#�ݠ�������Q���`A@�Z,��^!�`��À[.�bRo:�n�1@:�a�xwR��ķ��XI���L7�Q��4=5f%�ԑI�.oՒ��kl�wuw�8p��=����Xq w{�\�$�|u�L��
A^r=0O<9���'���R���!7����}���)IkG:��T.P8�8�f�Z`Ǣ�.�Kq��5���y,��r״�%�cQܨ�G{�E��SY)MC\ܝX& 8��sk�۱m$X1h[Ow[S�����?pNL���ow-9D�j�B�s}~�2=F]��v'չ3��u�:�^s�<4y�+�%Y�<'D*�vނ����{�@�|�*��G�]��hkV -�"x��u����g����g�wDC+��&�i�U�P��Mm{��+x��)��w�F##�hyR� 
�W�_^�-e�C6:�N')_�:V|YB2�J�R�.fK;�'i!��h�����u$S��%,��oR~�D�8����C��[�x(��ݓ�.�{� A��0���,blܚHnll������]�VG�26�D2&�1�_o�+�����mh8I�Z���[�%�4�
yJ�z��^�����g�_Jq��Ξ��s#l�UP��v{��eMP""�X�}��:o�w���[જ &�2���݀�]zq'��q�ou��O�S�WEi~���bא�(.�D-m�<~k�=�c��Ki�w�u ��xR��-־�ϋ���r��qܕ�\C���Nvp�#����qڔ�����]8q�(���AS������0�ې��jh����u�˚
�R�I�����u�n��,Z�]U,jX�#M���Lͻ�ՠ5�.���Yi�����$��g�彃�������@�n���.�(�Yow+�&����^���+T��( *�:�������=Y���j7�u�L:�l�Lŏ0�9�݈m�h6d >�ovufL�3\؍:�QK8���M�>��\V � q\��?�E�z9{��|�gRs�ƅ��m�T66h�)%F��FX@�m>��l��p��~��,��:��M��]�� ���&�q'ɹ����Njj�+ kL��%N��j����YTA�,y��U+~c�5�A�m�Jp���P� ʰ�q���Ic.Hz����n 6��0&���y��a�לX�x���@֬]+�¿Q�ny��I��¬��	~��љ�'��L�m��I���+p��I�v�����h9b 1��L��/��/i�����=gF'�<HO>����}VK�v>��ϋE��O����~��Lx棿q7�Z�����������E/����=Y�X��]��_�he�R��5҄1Ul����X&�]�H��X(�� �e����0[Y-z�G?7l|��N�_q������	���G����a�x��ys���U��*V""U�[��ni��¬,ԃ���Y�M-^\O�˾_�&�n��0�e� =��|>K�f»]����It���	wj}k�\����
�x�3j��ŭ� ���M�W@�0�SY ɋ�R�M��od��,kX���f+XG�ˡ�ֿ���e�u�ȫ�q�\��� �7=�k�:&���X��r�\?��^���[��饗^��)�R��J�$ʀ��Q�����5�;{��1�S��]^���>��O���I:�o?+�Q���nv(*��C�v������^���d�o�d3��g�3}�o��Yy��J�<� ��'��ZMq�wuu�ҥ�9�28����O�GP��n�ի/�x�׿�u'��  %ݑa+g5jѥ�]N�_�Ԁ/_eڥ*�Z��f?[k1�R�$�P(G��x��m�$�����
kS�61�)�Rb���Z��AèH���%��rܼ�87�B����qwaS�\c��:7n/J�Ŗ�o�)���*�ZNC��q� W�� 8(Q�O�igػ�mt>�q�wƅ��5X� rĎq<,n ,�vHhp�*J�_ K^�-o�lz�
��"�e�[s\��`Wap��;��6�cĥ�Ư���ސ� x�Bb�X��h�ʕ��?o�?����?J�����{ĭ~�ݿA��즙�I�ꪫ(NPWw'���� M��Pb�.�zzx�B|��p==���;	��O<9���'��
�K�6nX] ���96cp[')��'>A���/�bG�2� �����K���M��J����J&���k�	�U�R&\���͛����=;��?��MP�aʻ*�9�32���[��ycGs<l,�p4�ve��F0�o��	L�Un;Ip�RQkZ��N-mu㪥�q�|��o�r�-�%>�g��R��)��
���s}`���0����n;JK�햇=k8 �R������R�Rn�:S$�� c�Q���$1�2��ʆ&Ժ	nP�Qg��B \-��IRc<�9��:�g�2nh���i�@�l��2<�D��[ͺ�c�R� ߑi�g�[�Z�d3� ޢl�H��v]y�մd��z������wR*�A=]�T���d���k��B�n����o�L�TLhi���)��^)V��(5ZU�VJ�5�>�9Q� )��}�֒�O,u��!�p�̰59=�Wh���'�U<@�d!b7m�lJ$���VTOO�l��6]�H(L��چ���su�!�Ѭ
{\�Ae�[o�U��O}�S�@��UT�M��瞕����V����F�����3����	 ��9�hN�~�`�R�ʀp���E?u%�y_�bԢ>� GK<�  ��IDAT=��qmP�F�l�RS<�S,�$9�$uHJ�ڞ�l���0����ĸ���>H���A(Xw��İG�8���2�^sb�e�Ȏ �-�jK�ꍒā}� ^�@3�Z] �r2��ՠ!��{�"�oD�&e}k�x�r�+�_:�Sp��W���M�X�~�~�l�Y����}vv��;@�|V�E���Z��A'�?����}�u̕�%�� G�p��Z��`L����9��B���CM��*+_>>���n���xԄ �x}��s7��9���UkR��
�w�������_A��=��WT�������1~���M��]���gE5b4���NӞ���K6Q�.)��sA�"(dA�l͓"�{��;�t*��W�6�U������a�
�L�/ܬ�ûڐ���7����=���{����젩�1� �R	��ݜ� ��kW��y��!���W,���P�"� ���Q���u&�,(�����~��1'�q�[�p�la�"˹R-�\� A\^Cڒ�=���9�����UMZ���9��4$`!9�_�SW���v�d��$R�K��"�����
�6*$��b�5kR'-�5����5����+�A�B��Ut�����}o��e�&$�BX�B&�ܬ�R���xOغ.UK��ĲG�"��%Ȓ*���*�k��2��uv�H"%�~�gg��093+��Cg%N[�H��;	�OZ�"�.��3�~nEz�'?�G�x�*��*�Mf�?��(d����~@�it�����*�����$�y�(e2ݴn�E4xj��ŢT:!����x��M�w�<�����,H�ʵ$93I�O�hP_�Lw����;�r�jZ�~��l�Y�o@n�P�_̠T��G��c�8~`�2�TK�|��8��� [�*�Xr=����٪l:|�!4�i��\
�vOO7%���Ǹ�m۶� n��7�`�~�t$%�Yb��S��u��p��w� E�a��L�����9�<�v���9�da����`$((M��ϭ�El]�~[��xHx��I.(���c+�I:�Yl��9�Eċ ��xxÀ/I�x؀5�J�k3虘|C,eH�Aߕj�O ��L+?�eu$�՜�@�Ȁ]��M��o��Cҡ�(o��IB	q�}N" bߨV0��d:#އw�?��c�o��ü�P��X�9���4���
+OexP���C�Z�y-]��:{R4:|�zR��G?B#�G��@�F����τ}��{������%:x���_�c���Z5
x�y�c'�K�?�` d� O<9���'�?dtәEm�nl�(K�bcE���kN�2꒑�5���5�V��J�ҩ����V��>����Ӳ��ࡇH��'��?��;^k��}��w__�x���tR.?� �-V�C?|���#t��a�o�<��G�1iǪ�+���!�p��b�E���$e��0�X���>�E �@[��)9+�ȴӴA�R��� ��O�Ib�;�qM*�y���* ��%#;(�{0�\�&�P�xL�G��4,��gD�
�p��B�놵О���.b�l�SJV���(Y�����A�
��Ʉ�7��nHKS�������2?o�+��C�}hfrBX٠�4$ҐrDQ�n~�Y(�ihx�����I�<*"P��OIr�����b���Ӱ"V�	@A���������+E-�&�|N8ar,��+��Y^s��;��5�5�]Օ7�fV@����d���J�^y�5�F���(�	^�'D<@�dA�MK��X�;)�h%2A�9���.δ ywO�d����nk�?σ��g� ��������/e�D����:,4dH��;z�.�h-��2�\�H�S�vE��?��?����H�WwO�l� �:�Кe��{���2�#Ng6�ڵ� �|�AS:x�3�W�-Na2�5_.V[Ў2p%ө�u����Ը0��c�Í/���MX$���b����(�k��
�d��{�x|��_��&י�^�ZE�%��
K�������a��x�I��1`a>� ,�BY,f 2~GCAq�7��E�8�Qϖ�l���Y��QP�*�nQQ��(.�PX��|�,?�'�������2"���`m��(�����@q�� ��{��G�y��"�k-MT�)���$�X�8q��a��I�P�n��6ck?ϊ[,��w���*��xm���-���*+;}�������ӿ?�4=����QX��-z���nk��� ݓ���l�M��!�`*%�E������JĿ�= �}_�:tċa9��ba�ݷ�m�����/�"���K��.���S�pj�k���G�!��0`L��ҙ���A���*��)s��7���q��7�.c�F�k�lP��<��	�v��-_7ܶRBf��/�����8,��5�P�p�K/�v�Ԁ�s�L���6>��U���dѷ,�&G�Y[��2T��J�ɢ�
p#d�j�%���+<��o���@K̀��X�-#�)����ߠX�p��u�6*��Kh4[Rڅ<dv�
 ^�BMc�W���M���d,.��OGKѺ��\Wa0���OA���s��̦=BH«�����ˠY!�@P��vc�)�;q�f��@�@[�5�!���7��Ò�8�~���9ާ�T7�����/��l�w���S�*�"rEI�C�_��1���6�4�	���[�#�߷D�(�����N���5���X�N�'��� ݓ���o$��b����]W6XÎ��͠=}fHb���S�nW���1��}��ߧ���tzp�z�A��<����s8�1&��d:DA9}F�P�[E]�Xuh��RWWMLOI��d@�V�����+�7k�u-��ף�.��Rⱶ��Cn�fk�&u�dW��X�H ֶ֬�5�9 #����:j�9&�f ���^Ӛ̥��t'�qh!Fl<�U�$Ð h�֭]N�|^,aű�I����|>Z����,[�߇�8�-�φ.�89(u�蒷z�
Q ��J�V���c�T�NH���U�i�����0e	I��H\��N;NO�x�,^��o��V�x �0 V�п��?!����w�y���A6����ij6Oo��G��Y�D�4��]�D!��5r�x|&��xX'������饗�W^��nZ�%�w���}+!VLg���o}��������0� �CJ� ��4�5�x�%�8��%K$qtl�N1�OL���c��OӒ�U�۳�ϯ���T$:�u\�����,D�[��T����HxJ"��V����X�϶K�P�������$�	a�N� Ha�D���AGeQ�"�D���6ܯ�XR��~
 �a6�wl�dhLSņ4��`���-0Ŏ����g���{�b���7�-7_�N΂�^è�f�lߡ#��C?�d�+V��̧idd����L-wgG7��w�~�Q*�%{�7�e�o���6�QlS��y>��������]�{��R�=������N:p��d��d�����~��l�'��X*�w�B|��]����|�v�m45��l!Oݝ��]2�A��/�Bg��h��e����1w�	�����~��z�@=[�o`�t���%�ɢEKx]2��_���x�q�)�|�et�%[�][�V��s�O�)U�MZy���'����.
�T��T���������z����+[��R&/���
�m�7%��4��M����/
D�P�(ItH������h2B1�������]R7/��HlTyν�cS�{�a)ml�ZR��X�5�m��XN#g�����y1tOοx���BD�Q�d�ޗMd ��q��NX���%�$�	Ԭ��E^��H�\K6�m:���J��o�V��E�M��X�am#�J&EQHD#�M`�=�a?���띛���6��T�7)��I����Ufe�%G��MMy��2P�tvI����>i����D���ʒ�'s�{D,���E��:;��l���'����mI�~5�@H����.�Ơ]�y�x8�mX/�6|v�v�B���<��������u[.Ƴ�t���s�Je[��*U��k�;��o�*Y3����� �����7⽛6m�~�p+'i��ި\ ��
�5��:���{�_V�QQ�&tf������GB���7wʽ���(4�z�-��L����h���W(W��~��Q��l�PQ �	�@#	��5���D(B>o5�	}�x��
ڰa�x�6�o����_��dJ��9 �F˰�S���ߑJK������JE���n�5Y/S����s�����K�"������oyIq�\ � ݓI��-�am!m�i ���A��On�m��4o���2ꏑM&2����}�h4�@��Z�Ir�naQ!3:������t���il�,=���t��i�z�վn��4з����ĂW�Y)�e�>���a�6UbЍ
[�h�a��7v�v{�-<+|]�	�|ߥ�腗_�Lk�S''s�n�f޸g���Sgi`�R,��Hi\���(g�8#Ih�P�V��d�5$���H�ҩ+=���9� ���._��g3�h��u�b�~��/I���-��7����X� �����ٻTz���b��`���Q�Ҡ��%t�M7Pg�b�_�L�)-X�"4:q�v��K�}�q�����Q �`�KQ�a�B�4�;xB�������M���| 3(|S�;�y����J�x�:�h�"Z�j����"�Q̗��^��IRgG�^����t�C�9��t������+.���I���� r(s(M�W ���V�0���n�X�G������v�C��͐�P�C~~���NG�p���Q� �`���+|r<@0�t�� �唒��x Ȫô螜� ݓ�4�j��ʆ�������ĔNUHUZs-D�Q
,\��*IWp���X`��r ^r�܋�[�s�Q`�(R�(�Y�Z��W,C���$^?:>&1r�b�$YIY�.�������3b�(1Ďa�J�)>�932� �mۯ���)��9�������GJ3�2:<�c��d�pI�:���Y&�O��L�Ū���c6K��6b�]�X�P��q.Z���G��Y���]D��S��|�I��|+m�t�(E�b-����AɮwP���^B7�q��<f\ұXT���&fi�P�m۶�o���Q��� @!�V(AC�9I:�x�t�o~J���a,⎾Juw��	]{���{?-�hQ� ��*���xv�b3��˷���={�h��RZ��W��ý���hl|�b���*+=C��;�g��7���x��{���zy��\��M�>Bq�;��=|-tM#?�fg����/ì���f��=_�R�#e�<%���v��(�UC�d[u�vG"$\�i�6n~[і��2�vx5��Oηx���BDʩ�������}׶P�":ݒ��vS�BMwS\�`��;��b�lZb��
A���?3�"nZ���
՛����* ���q�W�m @�4q<�8&�,�����5[b�5��&e�@���|f8���#l���;�u�}�EZ�b-��{@�}��	ڲe�Wud�,[q��l.O-u�i�ԉ��,���R�-R��c�gF��Xe��A9[�Ӂ��r��C���&�&h���⎶�0�s�(Y�M����^�����*e*7��R��h���.�s����jVxjG��3�K�P��{�շ��]��$-_���}��5J<��?8<E���k499.�y���4t�5^���6m��m?:v\�+3S��� ��L6G����LO?���C�����*%>n�	ڻ�8�H<+��Kv�B��.	q��!��"pP�9�=j:�����W�����m��D��M�-p�Zo�I"%�:�@AM��0����	�
S�\�$Z�N�Q<ȊYW��;+�@� �f�&<QB��D0�NZ���'��o� ݓ��g��Δ�n����:,r����o$}و�Z��Q��>Ir��!96r�p�"!���b�(7�����,�T`++� Q>'�B�a�Ih��oI$�ʀ �+��P{��]��v;�jސQC���&}�[ߧo~��R�� p SY�&[�/�~���F{o��CE���I�<�����[c+k���aV ����M* ؎��dgs|�M�d-��=��E\8P��w�ƍ45��&"�&�RZ��赝oK���̔t��fe=���M˓�������$�	 9��`��c��� ��/��=��<߂d�/XD����?"��X	�Ύ�_�՗Yiu�(cKf:��@���V��s�Q��.J�%��X_(���3�TG���ɱ$��P@�c�N�:.JO�&�汖�7������G�֏�r9 Xk���^�΂�/B�8�;�4�U�9)}û��H8 ��+H���ˬd��=6x�0��~	Ws��G<N|���n_����,tOοx���{ް����?�B~ِK� �r��q@m��n	%(���GW.Բ��j&;k��1��K�M_�٬ś;���9J ��IM�Q��C|����m��_Z~�$�:��Ki���g�Rt\�A�W�Y���o�C���a�ǣf�n��ub��)[�9Ðǿ�d0� ��)a���m]�P�5*�*_.2�aE�������<F��TKb�I[XP�JO񀔕��	}��DCq�r�3X�ed$�	���M�V�������oG/om�j� �¶�Jf�P�>����cJ�Y!㼯�O�p;zB����4+E�V�����h4Ӵx� e�]tj�c�j�-�[�/�[C��"�e.��&�{���X���(n~��-�0x�a�<�O/�m:Xxe���>?Ŗs�-� ���P��� [ՠ�Y���GP�`2;A�**�]Р���F�m�T"Tx����9r��7�J[M�� ���y���=Y�����e#V]��*b��>@ +4�.�.Pd��	9��d%��A �q!$95�í�,p��[�$���rڜ����04� |K���E�u��v81	�8;���e%V���f�bC	Iwt�Uh�ƀ
614A�	_�[ZH����q�g��cB��x;��Z�����f�:"E,6Kñ��'�4 �������=B��kBꂸ|�^��fx�P�7>>%J�]/P,hQ�3-JN�R�{I�|C��w�-�nV��T�{$ �d�4幦I��;���k�/:�<��% ^����Л�� 7tzX��e�Iq/�k��xԴ�55�
fB43��ǎSO_/�-�b���6k@yj͂�e��P��Kaq�L����c4f7e]/꣭[�ʸR����w���X��R��� 㽒,}V�p�a�+S[�P
5����˚uk�ڛn��E�t��!�?�]��|M���O���		�ds���4�3�~�n���҇�=�߷�y�FώЩ�hz���v�Z��xr��tO$��ecsGb�:�2��c�Yp?k����l����'ܲ���!i'z�-��%�]N�>���曒T�:k0|�s۾�(�����=�w	� P�[ ��+��:�u6)
\�����S!��c����â`���B 1��N�ak�?�!������͖(@����&w:�I:�q�Mt�e��q�uJ��70���7hY�Zg4֦�d9��-	[�=E�*��p=�i�=�3$�	9N,-n�D,$D=�Y�Ig��T"��ǖe�ǃ�˿T4�x�^��lљkQ�/ ���$e=�`����#^C�1�����Icl5�T�g�So��$���u��2�t����g�}V����NnE��J�k	Ӟӊ9�rA����'����k�<C�$������ eY���[d>��iZ��'L{������Ŭxy������_#��fJ�P
���#s����ipp�~�� �ށ��tO.�x��ɂ6w��$���]+\�(W�����A���+�ӏB,�Z�.1(k��&���mt�w��eK�o���t��
D��[��=��|k�~i��@Y��ua}C�ݏ����(;���  ��/��V�	�ڭWI�b��_�fǣNU���E�fM���F]2���k���,��w8�Bְ��LM��@B�I���gB�Z�6�R�\(�6����.|�!���4�A��>�O�� H�H��ff�R�NFTD6`��S�dZ���a~���ʸu^d�Ǔ&�)`�$���5זi�L9"r�����fg(�Vw��)K�qAUx����e���Nw�4���@��M9W��F�(�I��4��H�zbt���;�g�jt�{����R3��`�RM��6�ox�pj͡���g��N�:a\󁠄�χ�<������zϿ�,�~���gO=M��w��\4�h�Ӣ��V�uW]I��<�,���~��.ɵ�A�kECԝ��y;}��oS��Eq�<����螼ga��|�A��?���������f�Iw�����/���/����/�Y��K�A��;b����D�:{���+�o�r�^�p�r9q�6���Y@|���j�[׀��Wu]>W�O�L�o�#�*=�� W��!Ӎ�n+��$�_��S�־�`��ҟ�ghf�	��� $�"�|�9�8`]k������0�|�
AI�d3�s /@�j���(,>IPl:�{�X樕����kbj�]5���us�c�l�2Y;X�Rg�{�g `�����J�ibr��#L��E2Z�J�Vt����.��l��&-�5Se
 �/I�ȑ�2���ER^���u����yxo��!� ��+n�싵	QFFƄ(k����!���r�B�H7�r;���������]�����A!�e��L��ヴa�
�9OA����K��י��Bގy���=yς����߸Q٪�w@@nw���o���_��-^F۷o�{ｗ���-V$ -������k��C?|�>񛟢���ߦ�L���ڵK@ɸӧ����Xx� ƄW�l�#�x�b��Jk�tZ H�\�#���k'���i��.h��ڊ�[�*���N�U!и�f�kl߰�ڮy <�	ֳV �&��7� zb=�
.��S+pZ��x0S�0�ឧf�t���3z}�
A�259.k�~|��C�����N���4}�Z 8*,ħ�-[�o:ΓX�H!׵��F�(�P�O��));V�ʕ+����xA�M0��N���������������G��s�o�xh����ҾE����>����˶m�C��Ν;�}E�/�k�v4�)I�˖,�5@�}2��	4��Aa-��7��}��ݓ �{��C���V6����a#�k4���X��+<ѭ��J��կ��Ĵ��ٳg;5(�/���/�w�A}=������.�x*���: 5��t�M��#����5�3����eLP4P�t��	z��]���j���Q�&�X��}�ڏ9�:�7�]�:F��8��5Oc����
�5�e�X�o��gpC�yX��N���R�  �g�tq/��(��k�R %��Đ�L;�UxFXWxF$��
@k��c� ����7:��k�-gg=��M���J�wY)sD�A4�����hy*�#G���W��k�,���IRc�6��?;�ա��3�s�h }�}�Q:��2A+hюgw���9+����q�g�ht�,m~�v��L�00��ė/a�P{i�eЛ=��Y�\� ݓ�,�п��6�� $|a��\� �K���.
��ђqOԉ?���Էh� 	2����[�}��t�B�����{�ivUg��|9�W��CuUwW�V��d���A����g�xl<`{�ƾw��0�x�����aB"��$�Z�
չ�+���|���O}�g����;�Q=]��s���h�+��]R��b���z�Fk��9`.(m��>H���c�y��	�6e�mن��2��@n���S�!h�3�!e �	a�5��&����aޘ�%��|1es�������vC�z}�d@�+�<^F���r�K�`����35R)�p.Ȁ1n�lg��NiK�d�T&˝���w�H�z� ��N�����:j�1xہUc�h;�_��╷����������Ӳ����d�k�����g���υ][��	���ɤ)|�0?�P�ݪ�^⽈�����߰a=o4g����%;=#���}2?�(�V��@��sIF�+�����{����::�et�vt|��%���eZ��Wn���5����3��X���p��>08�1@=��0�8!3
E������{�Z�܅�c�N���?�0=���}����#��!�sutu!�l��!P�Ϲ�\[k̜8d]m�R_����+X��c���y]� $�P'd�c�=ݖ~��vX��Ƅ}s��3�l
s�������;�0��E�Qd�8&T�}��m�b�0n��;��^�{�DR�mi�k�W1���G�.y���3���zB�&�o�?�0x���"�Z]P�=����aj#�
R�xsoz +b#�� -rq��
�q֭�x	��X<�xa���0jTa�]gg�g$��"�N�<!}}x�y����l\�ޤ+IP�`���ɟ<dJ��g�׶��?^*G.�M(��Я��j���r��.�Q�?v�8'
;���?~�t���	�5��%��|�+�xq�����f9t�|��?����}�a`�{��ˮ��
p�micNql��G����l�>,��ηRdz�l	=6�J�� ����mw3 ���-	?H	 ��}�х�3�,���?5�0�+�������jߵ��\pM�M�I�0�Ӝ~���'Z��$�">��Qv���y'��</�4��<���`XT� �׍V�����ǽ� �ix�s3���z��'�FMؼQ� �f������<@��F8d��T4^���M�ٲ6��x.\p�4x�h�{��E#X3|]�rz~*�5@ ,�x��G$�c�=�o(�e��#$��ڱ��@����*��!yp��p|te[\\����r��)��Жa����y�W�����u���(4�;{q������9������߬�fʦ� ���n����	�۽m����5�e�/6�/~���i�"�:� v��Q��-�$�~���o|��:��|�ӟ�������$���E6b/uI�%�9bs�!cJ���h�g87�k�殓�6��>6�%W��W��nگ�{���}ZAk���\`� x��7>g۬�
t��9-�����6��|{���V��FL,٭��a
�==}�t�1�u ��Jh�Ӝ�=�MO`�@8! [����(pA��À�����Z)	�k��8��{��[R�]/�;ɖa�����rǵY���À�����} y\�];�4���ݻ�u�S[]�	�)&|W�Y9��)�4r��0����(�HXz�����^#N���	���%5lv��'��_���iӠ���g"u�3��K/ȗ��^S�TV��t�>����������/�+蚃�t^7A F�T��L2�Qo0ɲ3l����w�#��{��06G�\�HＫ!��n��>�����g�zZFGG	L�b���`hГts������f�]Xs�z� 8z�(�� �0l���uR7��X̓�\;��ܻl%��<���[eJIs����es���|0b0OC��������kU�Tf� ���Bu��R��x� x#`�׍@�j���V�M\p���1��C׸y����>iZ��L޼R,N���iң�E��$	".�r)��F 캶�ز@�C��z���1��߃glט|�� �S,���<��јǎrm����Ǜ���p�x���#�BE�Q�6��ܴ��Zu^KM��ر��x2��3�����|��ߦ�8h�/�|0���e���5�	7L���At-�w� �|E&&��3'�� joh���b�g�Q6���:�!ǆ�p��܂LOM�ۇ�9�VG] C�2�������tx���<�-ke��:��>�|ȓzD8iɁ������쿭 o��\����zs��{k9�@ �3��}����i>�q�YG?xi1FZH}����P2��m^����6�����QA��C�Z� =v���n߹CN�8A�#"%D�50�E��y�X�0�.f*\�W� p<�"����n>�2�b?s�1$�5�r�:cȔ�mܰ�9���E�a�mw�����E%=���>�y��R�4_Q�(����_:z\�(�wttR)�H0�9@�#�m߹�]����S|���?����k�I5�R2���]"_]f^wllB^|������P4���
.;;ȿ�����*�G�IR��W�ZB�r�����!O%Mr���l��Jb#��m� ����7�R��9ZP�h�� �?U��Z_ޚ;�<$�
�֋��1�\�<o��wO���sm��[ ��Pxw��5<��WFH$��)��a}�����Ĕ��&vfχ(�A>���W6��مE�o�r˭o�?��)��Xo4���T?�VhZ�=@!�@0��놐<E]rYz֔qEY��M��Ƴa�+�l5�6E`(�����~�tQ�\({5�5Gn�|
{ �!; ybc~xs�v>��ǮSt'F�F�(���S�z�_��:�BI�l��p(�ү��y���Ɓ��ö�͆�u�Ú� OKr�zD �:���拍5�R8^�8r�)��q�&u�-�Hm]��F�gpp�:��S,��9 �5�iyJ���8������& �	�r�[s��m��
q����t6��V������� ��+�c��Y{Ŝ�b�	b�1s0�qХ�������n]�^�nT��L�z�p�NQN�>%�
�{��ǎH�jJ���6�5�|��JL4���������1xp/m�����8��]��;v�/��<�4��Wܦ#0�\��+Ȁo���)����@���oH�-7�D9Ԣ3�є��
� o���[B�~2�LQ��V����wn��sj���@�{WO/#�B����?����k!'�0�� s�dY�W��h6�.�/��ޘ�U���\��+��tK���18$9	vj8@j�J �8�$�D"*���-oy��f ���m�6��qL+ b���:}V���P��g]e�=v��َs%�]뫱�_�	�j�3�����|��[V�5k|���h%��i��"���w|�z���6�fЄ��=@�8���� �h�
�7>���)�֯���Wy����������iI�Z^u�����%N��i>h�kk82��{?�W�,Z�_�!Sv@x�~Ȫ��%���/��U	�׆띛ZKn����U�3Vp��iOp�G�����]��Vi��mV��!��n�,���@��n�^`×x*��D6_��06�����������Woe��J6S/<�S@2�%Xh�j��:7W��ꮧ4^Y4��K�� ��Lp1yjS�ddP�(�߿� m;o�5l�8� /�5���Ы�Q��;K�_-�����o�{�1l��z��k�߷[`�u��}���w�!�f+�{s[tx��l� =�%Z!`��M�=�<�{�� ��������]�D����3�r���y�69��1����<y�J�x�0L=��7�:�����չ�_Y)��j��Xl�2��
%�ݻw�z��5pıQ�������f�ƨyHנ��,|]K���:s�1� h�V1q(�z��x�L5�*���0\+jk<����m,�l�z�g�ډ���>��cMC7gݭ�£D9@�u��3�Q���Cx����dK���C� =��2���ʫͲ�uu� �`�W�0��?�yp��L�>�.����f���JM�א��̓Qo����/���][��6
a�gA܂j븜�g�G/��Uw޶<�R�_����u�w��t��G�&5�!�b�l` a��7ld�uY�ԕ쒜�x�Z �������D���IG@��Ȉ��,�T)@2V��t2�&�AKT0�	kzOY�\�~�6��½Fh��V �ad��?7`�g� ��#S*�=��#* �:��q��,�Q `1p[��k�0ܚ-y��d���xbX��qVv�\c�wt�K��KO_�	��S�C�����t�i�h�٨6M[O�#6�8��	B�W��]IR+���l,�`]o��0V,M����L̇�z�Qg��I=�ɕڍ`i�U/�j7mK��@ F1}�����l[[���0E�R5,h�G���^8F+��z���j��-�֠�����A͋(X�=�����A턬Gj<CޓP�A
��Q�hHtpTx�t:�y�K�=P���vD)���X�K��dh`�l��KR耇y���L�X�ujAO0�Q��[�'����Л����ܚ�<K� :oysH�bݠ�?48`*�\�i���U.Ŀ����b^网�̡gB����������1xL�]�|�n����V�9�ZC��
<;���A��B~^�=�k��>�lA��xȏ����1|@�ǚF �4�ɄQ�S)�ь�b!���b#��GISڰڳy�o�ES3B[Q��H4.����yE�˦[�-v��Q#���	�k��~�.=2�{��{��
���?��8���;����jq�~�VUaf��~mKU*��0�5� ���[�q^.�	z^�G~s^#z�����j�����D�Zq˿ԃt빥`t�f" 5��@����͕�C�RH����\՟w\�:!�eOB>1ak]ܛ�z�}�zyO� W�mfc\�]���-�s�Q���ԉ?<b����`}�j�\��5���B�q526����̜�-,Ɇ�Q�9kz�"�jl�a{�:�R���%Ϋ����Z�+:�tR����D�R ǳ�g�?}�T+�܌aA�dIH5x*%}�t�Q��.���ݿS�_�K6oޤ������3���_8)S#g$V#�Ts��Z ����s>��cM#��y0h���y���(��p������;�M���F7�����4D���_�u�����W��U��׿n�����������O�g�y�D,[�mۋ�C�Q�����o ;@�^l����f�0����䲰�;^7�R,����^QO�aIq���a�p�;���g�W�Wx���[���|ù�=["�Ӥ�!۽5�/-��@YԫC(�
�~�.1ԨL�ƚ"%1�i���*9z�;��V��^DUCI�4�W����+����E��C�K�(���֩
�0h��k������A1H����z��(W�sn�,]S���Y��H�d�8����C�F���TP
��L%ش��0�pm�@C6�둷���nC��_����i���~���}���H��?�+�5^w0�rR��r��>��cM#��	5v�d�!͛o�Y2�mfSv�}b�7x��y��g�ȑcܘ.M+���	���������n���У37��׾�� 
]��G� �06�����9�R��gIT���Qǎ�;�+�-�aZ|�q�z�y��y�A 7Xj��xy�&r�n����elm7�l^k�^|�-Ys\�<~��ф�i���[
�0�u£{\�0�Wn�1�v7���Z�����G�{��mrס�ð3�g`�z������@�.;��`�u��o �ϭyv;_��x��������$H+!d�;�u��/c����)׈p���V`�9lr�7n O�P*�ё���LMLJEA������L�kt4� ��q�M�9!E��2�gG����&���zi��ezfN��l�]ۮ���v�A�+�w�-�r]�z�yY��v���?~�t�i�B �����፾������6n�$�d�\��������>�zw�c�8C�P�;~����~@���:��c�tS�d&��������?N-�M�9",<5=aj˗W��i�x�9|o��-��mA�P��ح�������|��J#�vyk��Jt6��J�kU#�{�[�|���i�h�?q�ٮ����}�،7MϠA�Y0"��C��:�A27�[���˖-ò���r��Y�:C�`���P�s`�m�'J��.���nkV����`���6u�˙�V�"hz�AY��)5y��@�Q�L����RA��#b���z{Q;T���U#k��B��k�uިFNJ�����h�����^��ލ�g���Y��I{w��~�����2��FB�-��9�?�q���XӨ�kRU��-�bY��ݢ������m�2�A��B����t�b77�?������%�zs���	����Q������W
� �'�x�" a�{ʪ��j�PR��6��4*a��~����K�����5�L.N�<L�"73=I0@�S,���^���P�*��Pu�-J]vÐ��ϴ`;AeOػM=�)hx?�����������7j�W�7]�Ԧ4\�3��n:��n� ����3/�m-����e��	i]�#��W;>!A=č7� �>KP���֭[e�SgϞ�rY��|�5��F��l�A���|,Siz�n74��ѿ<$��ݿ����x���nx�(���=����W���СC$G6�$��'@�=��hRv��*��.9v�%�d��yۡ����)i��������28�U��y�#�n��m�d|bYzz@�t��a�:�MΜEd���,�{�?���*�i�YZZ�k�����u���76X4��|��%W�����[o�E�/O>��ttu�{���?���4ù�f���~&��47_��` �v��0(OPT�Æ�o�>���[��36�q��͍�B�8�?��?�0���)�3^#��@�͛Ӌl^V6vY}:�e�l[�e�f���*��Ps�d���r&��i�_��1,n5��HC��Q�4�d����!!�c[[�s�[�~��q���kj�D���/���{�����c4�Ф�(�x��s'��19����G	�b�6*�9�o��=���a�<��u����?ał�G��Q��s�ѐ������f��O����L�1l��F�͸>����vٹc�������7dvz\����ר��K>�G�B�!CD����v�^��u���������XR	Rc�V��m�*z��?�qŇ��X��<�фzT��é7O�	��m�)��P���
�䱟=idV�Q�Q/�����Z��M��}�ѻϴ���\N�]B�W-W��3#o����K��l���m[=��Wu˓l.�O��T���H� ����I��`��h��J�Z����D�4���nU?�^3�I�a�2��y�4�m��j�5����i���+U� ���e.h�a@H�Gd�9q���V�ݜ�R,Q�ϰ�������F����ر#Kܣ��vr(��.I,l���&_�	���ȱ7A'��8��ޖdffNv��ӝ'�[O$LDP���E�[(`��T�&Ԧ�N
p���Wըsy�cM�+G����|����Ї>${wl�'��̙3��kT�C�~��i�O�T�����s�d��k����z��e�����%ԈH![FEA3oT#��+E��+0|@�ǚ�eq7ݖ�`�:u�`�\66��۷��8�4v��Լf#�l���U�|�m���N���۽[������mn� l��cQSS�? >�����\<�v�qwYAɖC�Z�2�Ǧ�6�PC�w�kY�_2��՚'�r9�[��V��)Y�-k�ܽ�W�L`w��cY��\.��lNٜ��*��W��nj�];��!��
�Ș ���f��A6�]ط��^+��_|���ad��7���.z� �h��h/�ʔ[EC�9֤TA�yUBј�f���z�Z�/j���| !l���ٹs'C� ��8}}��F��&����g==���ɋ��X�Q�(��u��۽{��+E��C������NF�%]���y�'���C���^�,�[����r%/�Z�O��d2-�@��,^�}�?�����?�4���(���2�6-����	��D591-�z���w�U��G� �4\�`C^sÍ�u�������%~��������^��o=��fmw2x���m�/-,�[��}i$G@�.-3o�a�8o z{{� ]��Mb%쎕JJ�\"�"��d�bg�l�6��k ���uh��fϚlg�u˔� b �{8��F�5�V|�|�=����eu�	�SBTA�ꖙ����/5(��M��K6�g̞��XHz�*���0�^g�<�&5���뱣w:J����G~bjR��h�����hY�4�P��t0`*�X�X^Z��~*e5j���:�+2>>���߿��b0̬qo{A�- ��O>��fg�=C	�ǵ�^-�Ϟ��+�}Aԃ�	��J��{�����>" f��c��@U����YC���%��Y�����ַ�%i��%��:������y�z�U�4˲}ې�בpD�U�)Sc�r��qpN(�V*���:���?c���5تn��Ŧ51����/���'HX#�;veD����􅍶��\,���9i�2`�:�B>'���7��e����bk�0���'+~G� �f ���>� �s/^"�b��RO0�{4���<���q�QR��g/��Q.;�z�Lڀ=��^����[�4 c$�`�Cݭ�̴6di���a=�ְ�%��0~���0���|<kݝ�[Oo�������_z�`��ॻ5�
�T�����W�i"��Aq�Z]�X$J�iE��p���>����4,t����[���5��&��6���^��H�E�d��FX҈9A��;�6���3��Q��x�0��F,�|Au^�1��hg��;?}�a�Q�:	HBAǕ�I	�ejrF��ѹ�lz���}{�Q�Mm2�Ve�sU�����^�ׁ��
>��W|���5�f3�膉�8�^��Jy�$��t��;︋-9��x� �?���N3�y���|�m���m�߆G�[\��y����҂�)B�O��S�oW�KGw+�P�T��f�)�T�b!1���n����nV�4A��tIC䉋���aj�Zo7�Z[m���j����5Ք8%O�����g[��Ȑ��mLm|Е���$��rͭe�w*��]mTV��� ��b��D��-,����NO����Q�,+s� c�ܨ�,B���S�-`t�BbY�UH0�p�q5��~A�!� wWW���N0�uvu2T��	��!.�HH{g�YI�c}�Wx?a H�h�-C�������{CC�^t����/�Vs���D�=��ޣ?9��s���_j�1�E����>��Fd���n��ߏ����3r�u��dzvJ.����Ã���6s������>����������?���?�4�ߐh8ބwo{~~Q^z�l�&/�|Z������������x@^>u�~iR4�����g�������u�6��|�	��*r�7�FO�Q4���Z $�1S���=wA���0o�>�cs��q��V,�x0�OY>��z�+�᭛s �1�o��G)H}x=d��(�A:���0*�M�S6��a�ݩ#�J�yP���V_j[ƅ�wȕg5LzSgA;R� .s��1�7�=_w�ǫ�0����QO�p� 8��W�O����.�W��*��Y�g:�y�{ט��C4em:��Z�D]x�������4�:4�����=������-2�e:��KGx�\�ɜ>W�r�Ү�x��z��½2�@
c�뮣�����3�=�J��h���:�����j��Ǳ�:����"��a-��ߦ��3��]ݡ�ۙӣ�˖dpk�l�H ?r�y�_�#�5��=��lX�E�iR&g&�S�=�����k���u�o h�	�g:ɬ>y��I�p~T7�i�h��^^ʚf0��I�݅�~�(�?+�>L��h˨Wm�� ��vd�l������Q��ق|���'�m
�������Axmذ�ǄW_(�G����e1=^�^<�B�@�,p��ԃ�!�����6<�&<s��m)
�n�æD-�^(s�M�öyy��r�g��I�O���:��,���o�w$cd@��%ṃ���m���0=�Æ�1 �Ss[�6ٳ\�?�� <�'�=t�ۉ!̭d��Z*r�;�h�[Tp���}�i+�ݻ��gfv���ɗOH�����Ay�-�@����Q�6���I{DȡɟlKJ�z� �Af^=�EgDe�۵g?�?�{ ���s��2�Sn��mN��> +���`�ےQ���k/�L'7��ժ56�!���Iy�N����%i?}RbI��'�ʲ�}@6nآ����25��J��T����?����k�H�V�V ���7e�4�Q���Ar��	��B��+�B$/�8
 ��0�I�8�*ä�2O	d<|ozӛ�����f:��z�h�^��Rf�D؁9���@��V�6dfnV7�(ôd�Cs�bZ��s��xn��>@ǲ�추̦�n�u�6�nAyi���0��$2�P��W���@�|B����.<o�q�6o;�!2`Z�<� �iy���Ca��r��]��&��{i�	b>�J!���}�5L���65A�$���7��55��248�X;��6�z_��h������EN�>+�7�~��\�(%]�;�Cv��%����(�204�u���&�g�ѨŔ>�Q��s4� �8��A�\+��>�N(�C��FF�"%�۰�k5#��`ra}¼w5�*��
��-�|���{�4�D����%Y��Q�!ېD<%�|I��e��I��$[\���E?��+>|@�ǚ�n�
�&6��zO����+����I�� �rC��;'ы�%���	`Bn�eL
d�j�9g�<!�[��� ��52��������p�zR/��^w���h�ɼy�j��MI���<?�<�9e���a#XLE<�ƿ	�֗����K>�#+�
8+�
�5�h�c�{-P]�a�۴M_���껣�1="^�@������_�9ã��gaLDlq=�e�h��LM;^�@��Ԯ~��g�%[�aqK�(K��D�U_��u���� �d<f�T�}�(�r��E��a�᜷�y� ,���=�Q ���^�����E�٣�>*�Ϝ��}����,�4�A��1^������+�ë��Few���xݬtp��&2�;Gξ���Q��쐅��������Uc�rÅ��W�@_BN�HG�����d��������FS��P5D�[^
:�]�{�PY���:����r��>��cMC����n�u	Q �1X��FMA�D�V6dL7C.�K�)�~66Qq�w�b�|'ʶ�j^z��zd�����?�b�摡��O>�6(A��.�yF�ۄ�Q�D)PP���*����֬q��EbQz���V+,�2�j���^��@x^����~|�q�.�° �?�k�4Iu��\P��`�	����i|�R�!S:�V&+�ea!G\*�z�!o*.x�u;�]���C!��0��L��Fʼ�o��]��������4U�@���q�=�5�u�����z��>+��U�0�əI�bB��@�%r���|�vf���l������O��=������g%,h!k�:�!���F�L�&�4X���0�kBA7҄�EU���K�Pgi�4 �8�魞HDP
,�~��W|���5�$��(�{c�ݪ bRwI[
&�D��;p9��ۄ�����֧c#N�gX+�<���n��|��� ��|�Ŭ~G=l΀0�u�B�Jd.���YP�;�y�P.	��-��$�������²�/x�M��o���qYZ���6|�g�H�P5 �H~T�Â�6y�eUM��n�ۂA/� �+�(��L1�\�2�v@�4O�6���������"��p�נ��s2�D)W�v��������^��B.pc����S	ӏ|zfJ�%AC$m�(���S�zQ�%
~A���k�=N���s�@ܛ]�To�&ۆ����	��}�w�C�^dU���r���n���H�jD�pȤ��r���F6u����OkL����FZ>O��{,��%�? �`\�����`�F$��xlouMU��q���2�{iy^��9��I�hV)C[,Ȧ#?��K`AD�����t�i�&٬Tk�tZAP7E���� �V�C����5� P��3mo�.9`B�,!�b#	L�j��
9��Mk��$��<����:���)}%k�Y�lg,�W�y@�T�~zbV=�	�t!��+����S+��Iӫ��'6�3р�фQ������饋�^'74������$.<>(�a�ߵ}�z�������C��Q����'��rY9~�C�����wk�U�wh��tu��>��	���m͍^ ��$�����#R~��@$�9�φ�r��K����o�󇟣�Q��쬦�_��M+نa��-1�)� �l`�.pI$�TP�WKq�gz�ۥ��]N�,�^�	@��_f��uF�.�6�	����c!�Za#���w5���F�@ӕ��y��Z���ť�٠�I�>GjW�hj��}�� x�nG�!�H��"�XX��y�����~>��~T2m=��-������_J������qŇ��X�P�ht��*��KC/�\n��^ �T�I������M�d7x�ꉖ�C��j�F�g�H.��s���3,�4�j<��1��!�;'� d+ �[��V���?$�sFV�:�A��G��Q6����S�AH!蠔�j�4�w�K>����Y�Ruu��W��y��#���}���#��=��#���*k��^s����~�<���tD8�M�T�f	]�tB�6\�ŵ��`�
C�6z�l �v� )x���[���R���`yi^����y4�5+Ive��@�������b��z��0��.��gH����w�y��A�!�
��:�0�q�A�Ȣ'�ta��Bc����0�<Po4��m̰Z��|�3�D'��13��k�W|�k)��:xn�+y�5�y¬$�[\�Z�b��\����#1MF$���w��,[�o�s��?vF�.N�����3R.d��y�$��D�����>��c��̰-r���.,��ع���zol��J��[6@Q��w^��=��ϡ�	r�d��X2�\r�\MC�B^�%���ͼf�9MO'��F�V���}��������0��8B� ���{<�&S�m�vu󭢆H'�:(/�:*�3�d9G�	F)F'-��w��C�do�����/��x��S#类e��낡���`=�͛[�y�����@iҚ�<�aU���q,|Ɗ�@�J}�*�q~�����|�����ٵ}�!���`4F� QJ�Θ�ó���	�4�X�.]�����aF<0�H% �9S��j�Ģ�2�՟�U�z�(�]�������V�{�d�����&nK]Dq6o�*]ݝ��Ϟbi���_�2RDG=��T���ַ�Cn��ZIgT��h��5��K�O����,�g�G��B2������>��cͣQ�9��J�y�ݻ�V0�C�W�͐�������[\���,7�d2BV2 
�* 0�ᑣGe)��M����!��g�s] �
1�t�ؿ�Q�b��A�Y�z�;�)5>�?M���f�B0�Z.��+ez��.sK3�O}������o�>��?a���'C�Z.g$m��cO(����G	��؟�ѣ��G��s�����^�7\Cђ4�,�f2 r�x��`G"�'-����W�8E<@%�i�z!W���'��t���d,�5�-�{MI�9F�F/�5��xX�[����������駟���%��w>�~��~�9FRz�yxǕkֳa0�i��F��`�8zI�7�����0;�_;;���3�7��u��,4���Yo��W��xD^!����w��(��+�K�z���c�|�4���+���QCi
%Ӳ��5r�w��]~�]�?�C9t� ס�/�tO��Pj�Er�{�*{��A
Q�n�N�@�	y��o���я�B�CV��p���^\��?T�XӠ�c 	��[���@�*C�[	�h&�����ʃ>(ǎ'�ՋɤۙK~�-7˯��oɳ�������JF��dS�|�#�ǎ˗��պPn�o�	F�ǹ�X@ ^9:�m��y,����^�����u�����������l	�P�sW��A�B]4��G�`�7��w����FдE�X��C�=9wa�����C�<L��-�~�_Tb�*jL������e`[їŅ9z���?��gE]C�%�
(
���Bj(u�8�=�tMC��&U0���L� t&�Ȕ_a������յ޾}��3?*���mD����
%8����;��v���Q���*�K:ʨ�5;;O��B�mɗ����T4(|F0Z��[�8��nۜ�����:^)!����r^% z uO?av��'�z`-�I�馛Y��>�|X~�C��~H��>'gϞ�p��,7��ZA�
啛7m�L�S�&*��Q����!��?��W��?��_g��_��+?|@�ǚF5�C
���$�l��P$�7^����h�w�L�|���x�[�y@y�Q�NwЛA.��F�1�Q��ߗ���ߙc������}���,�y.�f.n�}7��
�
" �q�׫��w�Ni�J��N'B��W�E���<-[\��dQ�htbC�򣅼l�Mzxh��ղ��B^&����]"��ʳ@.����
�ǔ����qΨ��p���:���wnf��@��I��0�57G^3�gXw��k�f!~�R+��S	�>�29�Tb�� �jE^��e��C񦇼έ�`ڤ\�J0&���^��M�F�ɗ`]�!jD�at�PF�Ȉ�q({[��!�e���O,"���� t�<F�4�g��ӯ�5����0��Cl4-ܛ��d¹��_o:F�'5� J|~$H"������c/!�mo}yP���'�OY��Q~H�:;efzN6o�#���,/��5�*� ��B���|�����/ȷ��	��D*>����������)M�|f�	V Q�۷����g���, 
!����]
zq9{��,N�yݲ <_���S��3��������-s�=}���s�*1��5����4��Q�de=��GH5�6�m�,�596&��u���?:��m���Ș6Wq �3H~ �b~YN�|\A��^v�:��j(H_o�[�m�V�8w�0�K�z�;Y=r�i�	�k[�]A-��蔅�Y�o��N���u� �.��tU
9�Pȳ�dm������߬�/�=պ���py�1�}BD'nr;��i�K�|l* QF�n[V7�`���#2`��j���r�t/t�
ޔ��B?W�A����.u��ra���z��5�x�F&�D)���՛�w�Z"H��}'H��v/ n��(��ϝ����>����c�ʁ����	\$S0���C�%dzrN�}���]�7��&炁��P�988�H����M/p�\���?�4b�Z�Tk�Me�"B���W�9ܼ�(�˞���1K�@�Z�Y�fj{�C����C|�a��[���{L��կ�.�N �nIV��!����D' ؤgg�)���8+[6�JL7߶d̐��3����*b`e�T	� ���%��^8wV��M�a+X����q�dȘv5�u�G�p�.�fX� �z�������>5b(��h*�6����iv�jWC�7~�ר���=�k.�)t���z^�P�jJ��J��%�:���̚�q$�f*���� �(��$Q���Y��:�ޫT��wo� On�X��^wc�-l:�������g� �e�с.�P�P6�G'9����B:7�Z��9�a�(�=jK�IN��D��J�F�h��	p�HTpՇ��K>���p��"�2#�����g+K�j ��E��qGf���dWJ��}]�v�87Gc���G��v��H�d�\.�f�O��Ǖ>��c�����-`X`��GfeH6�1���h��|��?���M�3�����4Jb��������27;#�(7c9P�4�MX7Y�|	X��	�<��&=ƺ�+2>rNA�(��+��T�Nk�� >���)�---�-l]�Y+d~nZ7�H�ʇV�Y��rY����M�7̋m_�ˬ�ZQ��z�󞷜Vp�$iBA�9��[� ���8�jJ�:�u+X�1�Tg=r�;�e�g�n�Oۗ ��zq��R�|��v=z\�]w�E�8��Bd�х`v�z` X��%�Mc���h)���B��� ����[x_ׯ_�[7"P�T�Z���{��7�eF����G=;����A����o?�MF�z����M�:�)P*$�HBд��<�U�OU.���� KK�r�vIb;�����]bJ��^x�9�ȲGI��4�32b����W~���5�����W������U�Kg�R��٧���m;to7�)ȑV�B��zT �)+'�̵�u��jb|\��mRW�|졇xl��$K�T�F�|Eo����e]q����ղ,.�JD

���b$wU��u�գ��4�F�@���AxBkMGj�<?#�BD�ɼi�45�Ã-m�m����/��{I=u�I������xT&�'$��T�dhd���<KW$ƂY�1��֟dh�z�)��J�P���J��l"��,�������[<`;���y�)�}��} 9���Gt)��Q�0]q�,wH���������:��%���u�_/��v��;{Vv��Ő6�~%#�J�Q&�0�b5�"��`H��^q5�md{Z�BFx������/�'�5O��P�F{�*CC�d���|F��eٱm����;���#������aUc��1����H70�Q���j�ƑZ�,���^d�������k�i7t�l ��f'�т�]*V�ĉ�����������o&X �N�:ɐ9@*iw��fy�;}D������(�f���w���<����L����:IQ���Gp�Ў;�˭��9t��g%*K[<(����R��3��lF�6���1�!,�]��ݸca�N
Z]�e(����
�mD��-� ��ԄMsA���\��#���5�rhd�u!�aj�a �c	�*@���]ު��6������V��l � �W]u��>��[n!9�閜�gV10�k0 ����<��K4f>���< x�]��9J���p	h��+r��5�H�����fm7�;�SuE� �4x�ֽc>�|��kt�q��G�:;���V���D��ܫq��%9h�5Fkt.[��G>�����yV�0hy4�����y���^FN2�i#��S�fi9+�{evnZ:{���BC���2���j�]8��<��Is8���D|�8\���?�4t#ut3��=�ϟ��'H^V3ܶ��P.�ȨkF�^#  Lq���=�y����wȗ��W��KGHx�aU�<[lбxd��u�b��0jv��k��k$�A� 뜓:�D$H���"�d��Q E��[�����ʖ.�O�m��J9� 4���T ήh�0,��S5����o�z�祷����uB��Z��!x!�P>L>����w�n}���_8K���x.���+܉�1y��ë�5�����3���2���ؤ��؈�����k%e���M���=�1���>�nc~������M��\<���ʼέ��O��LMN�����s���x�M�Y���hg�?^�"�>7;e��z]/^"Y�\�$/���P�һ8/�$��)�k`y<�V6�~�NP�@�z �.��}��RC�&�TM�yW�gd����;dxx����mˤeQ��~���)D����?�q����X��� 6D��'�ƌ�Y���d��A�]�9�`�%��͸=�EA�H,,�N�����O���y�ͷȯ��W���wI��>��4�<�����hl8��0u�M�v[3�n��*K�����J�Vd[�t��
�(�p4�8%��$ �As��Q�Ԣ�=��Ky���%J�
)�	��=�Րn��8���cc�= �Q��k�;>�P5�Z.�����Ly	�@���_'t�����ko���R܇^��7 Q���I:��W��s(dڮ���Ju�2��)+ ��-�)�;�|�z�{9?#�[f���Q�&P�3�~[6��=w��q6_��P9����fe4�b:��"D�D2�vRC�#LO�\J��['o�ݲm�V���ޞ<yJ��'?)+�շ�wP�5� n�*z����x��0��H4�D���K�R���_�*�\��Yu�k�n���{;�drbZ�uͶl�ȶ�'O��tm�	9u������G�R �T��Ҭ�ү����t�i4��F�Z�c�d]�z6'O�bh���+w$�-$ �z��Y�s���|�BO'�J�8��;����;��vپ}��7c�G~�f<a�t뵚+⊎8׫ss��9R�
e!(�U�:G��y/��W0Y^����V�H!`G-8�u`�c��}���G�ǅ�]c^��p���Z�9�ߵs��O������t�����:�D������K]����+�N�� =�Hؑٙ)J�"b��ɩq2��m#4��
`�]�X�U5�r �
�H�W��5������ ���7�5�;;۽f/5�,�Q���lgu�!:Mz�8�q��;(9="4�KY��-�d��-�Hld���|V����&@ ƎH��s�ۆuM�4��ظn����M���?�jԔC3�z%t���b��#A�e����t�{��AӠ�^?��Q Vm��Ke}����� ڵg�Ԛy���O�a0-#�r�ܸ���mvhd$R�ME��\���?�4B�jM7�jQ=�T2E{U7��G	f��F'�%X��ErU"#���fB҆U�T/�4�h��˩��R�B�
B��U��[���NZaT8	���J` *�r�z�ѰD�;uСR��?����;}�W*��`^<2��I��?��8������0q<s�����i6��U�>x�흒i���A����\��5��nV7W�&u�a�[� өU��s��#��e�fF?.�^4�YP��*p<�t��Y�Ww�P�)"�qY�h<�na����|�l�
p���Q���ѰC5=���H��Ԅ	������6X��tgR-��f�(��J7��!Du������"�kK� Η�<�GF��c t1`��p��֢����RL����?��qIt��E[�-r5�QVW#�[�:�8�*ӳr��9�iF$�4R���t��C�P����pߛN��s�����t�i4��&��lU���zW�*��e��"��ըkV���b�$+%�IÓwL�<�&��պd�&Ϲ4;iJ�j&�l�=�wǭ5���%fa�&Z���ї�pP��f�f8����ˎ�W.������z���^-��.y�Ǐ�7���v�!1-/����D�0��lRwtO�����<?)[�l�TG� ��O�����}B	�,Ǫ�<�����j����Fo�i�#�n�N��W�u�ᔔ�
: o;v�ӧO3V�v������y��S�`���J�H���;w���ٴ~#K�PB�֞1yjq��r����:�x"4Eɥ�za	���,� �0k���/-/�+;��*�DX�o�Dc,�߁�W�TɾG� ���bY.���Y�V�(O0	�{]�UH��229�޻@=�?�������b6+=@���7��0)�l�w�x6ݲ@�F��t,B�LF*��|!�ƕz�ͤ�䭒�AFo��ˬ��ձ[bm!ܧ@U
~�W|���5�H�� ������ag�A0���7O0��E! t[���qB�:�ꜣ��<�*�Q��-����5�Mh��^¼�xD;��X'm�w9��G�n]ꥢ�WФ��1���M"���iCz'����S&�9���J� �K�g�g���X��Nm�~Zj��C�������6��Wox�>���Fl�¦�5�Hm ���"F6@�ꫯV��J����Ȩ���2�~�5��Kޱc�s���qZ����E󛠓��������\���# ��^;�[T��� �
!���Ȥ��wW��:#$乙c+��5  ������$P����T,�.{�\,X�����%�6՘Hv���#r�M���g/�� hC� ������O�<"cS�rn䒫�J�S��+D�cP��G�w����%�< !$&#��Y���UP��ep2b�I��6��tvwɥK#�z��{�����t�i`����GA)
����1����Y�i�U��$CA*C�5�ްYb�E*4H�T*��r�h��+����)S5�&w�r 5��p�zu������|��>�M�z�[*�td:hl��Fn w��A
�X(A[(醭��ut�����':��^+�gQ=V4�V� �\%�I��w���F����u��-Dqۻ6]�q�Z�k�
`� � Y�|�@�%��J�����MCU��s�=�p4@9x��QB�k�5���#
�(jS����F��2��<뮤+�*�x:�L{(�Zq+�cewm�[�m���=oaaY�zz�q�	y<�~|>m�z�l	 �~��ep`�t�AӖLH~eI�;f�b�ոskҋ�[����	U�g{̰�+f>�s�x���z͓�]V�Xt��«p.�lh��'����>�������ҷn���-��|���^H:�p"����Wx���+0�&A�Qb��Qjs7HV�i���6妘͛���s���C �B�S=A���`
��гf�<A�rɭq��f��#<� ���e<`=�Ԇ�p]�_��CE�2��j�l�(��^�{{��H�4�[7�Ύ=W�ٙEI�z<�F	�����D����/2"�����'Xg��Qo�ZB:������E�Y��|�-[1*��N2���a����?��"1F�oPs��
���%b���K�ZZ�9�����VkޜZ��و�a�7��z��V����[>�����_��Ӱ����aG#ʒ4��!�������/:,���;�-�Fq�<>���q�&���Q�'{h�t}@l�46.��;�Ƀϫ!�Q���r��g�۷b�P�Z�����hB�`tp�s����EYX��X�j�Me��Ek��gG::2�4���U�/[�Ǖ>��c�CA�ـ���/�F�G���Je�QsHÎY��遡|���ێ2�is���!8S�DkM7R�]�+=FD�Qz�����	�E��u7���y6FYkldLNC���T�]\�ÄI�2� �ĨS�j�PΥK�$ԡw:j���JN��G\�6��+պ���V�a���K�^��-�4���bv��5�aU\]ץ�z�f������3JxV��j[�^w�u\G���Y�LO��5� B�����G��O���WS��g8YV��Y�>~�!�^�4\ϼ�}������g)#��� �J<%�|��	>�> ���}^1B�US+��I�S�|tL.\���4=s\���3S�$�E�<���{�9
�U��r-�Ȫ��֬�`zJx0�@z���`�W\wE���H�1}fhH���5�@`T�X��J��tv����˒J��R/�ՖK�\���?�<���+XBp���P&r�|݄Y���yt,q
��   `����� �h�V�ȯ:�XG�8A/��� �p�R�*��8۔* cSooK�U��ܼ$�	ܺE6o��/?@R�$>�<tȈ���Y�~�,Qݤ�If� PO=�.C[w�%�XJ�9������J!��f���$��6�B�"��s#���	Y[0g��Y���e���OJ��@m?�nD ֶ[B� S�C�B��>s��돂�`�M���0��M�$���;^��J�ڹZ�����o��L�\�~׉�x_��繆ۇ�Q%�2��w���|{@����g)�+j'"!J�ί���_��du�hX4k�� l�����/�ᾰ"A=tk(�l蘴�s<s�^�-����D,N]x��M%��yY��!�w��۷s���)y��ef��5[�|N�DH��+����t�y4�=�:HF�F9P"i�LQ�l���¢,-�P��b֫C��P<��':o��sG��? �!?�+�B ���!�f�5�ho���*�Y��_ݽ%�^%�bڻ�S�dp�f�g�����\������zva=Ζ�����m$�ojfR�ф�u��i�y�=���Ϊ�0��I��}���BW40����]���a��''�[���58&&�x���?�
�Ü����m u�M7��j "�mɂ o��<�Մ�qX����%�����Y��bH��T[�hq=������|k�`�w\�_��<�&`^����q�u�(�C�8  |wj�]�pA����F�%�鑕|I�(��pj�u]	ئ�[�l�����v�f�H�M��y&K����yí7˥���}N&���{�<s9ٱ}��z�r��z�	��x�����y�����{5�����IN�������?����kIݠ��Ն#���G�8 ����:sV�=��.���b<�-[��3:�@X���mf���$a�E��;�����F1��)��V�����[��f0,>�S��L�f�cW2u��.�NJD7���.zWTwS����Y?�3��` ����p����z�g�^�&<z^��\���n]����;Fu��X�MC�C4� C��j�~P���37nd�^�a`~֣��Ȇ����>����a5W|ǒ��:�`�8�P	i�+o����l�%<o{����Y�Co�����o# 6��,�0��S�#�x����%6��f�eQ5�`�A�R3lw��g�=H&�2~q�M]�MS�\�l<k��-�ɺ�xl���mI�Ӡ�~����P,�e��l�ݿ_>��2��o�n���O����܌tw$�#���x��/<���ڳS��}Cy�?�Ͽ��?���/'?y�Q*�e�#��Y�����t�i���$N�!C���k�b��SA"��2l���c��?~�sR��f�.1ݐ������ o��w�'��������=��Gn~�M�я~T�yɐ�Љ�a����-/(��Ԡ���_��~���_���u��Sϱ�ȴ�9�%?���g@ъ�P�ʱ�'d����ꖗ�gX�^�~R��!*�^�z��<�>|�ൾ�W�� ��wu���#/����$S���:{�< ��L+ЊG�<� �AOT���ȁq�g���)� ߃�~��E�Fc'�r�x����,�Ö�^���Ld3�=&G^w�:�RF�*v�z}�-�cbq�n,�� W�]� ������>�@�i�Z��9�~� ���ٕ�qd�޽29�,�?��z�!2��w$J�8֜C�:�
�xf����ױ����}�g�;���9x�9�������]�?�W�J�z�1�ʗ�����dqvE.���o}���}���p̾XSx��e�Ҽ;qZ�$}�>���������\	��2��#;vl�M�6�溏^�m�NeR)��;\������l�2�(���� 7���	}��W��x:!��v������p�;��`����{v;�5�s}��!�45#���_�׾�f�� T��g��JY�($293-��{/�Ȇ�cy¿�ύ7�ք��+��j�����6*_��W���z\k�]@�=s����S'���۶�~z}�:�r��r�������42���ϛ^�\� �u�B8^����� @p��[P�� /��X�]�x*u0�,Cݖ����՜z�#陜�+E},�φ��ZY���0��"��ɴ��A�@(���,t@F˲jCRi��(�C��-x�:$m]�no��SPc45�t}]aK]7*ck�5A����/�2���|G�G��GDׅ�6mɌ\�7�q�������d߁�dyi�kybD16m�,��^:��Rsr�jP��+<|@�ǚF6;ӯtJ� T��=�j��<2rQ�h^�y����v�ǎ��������<�M�$����}C���������~�dey�� Vaݐ��&<�/h{����^�Zv�ؚ��� ��c?���2=�@��w!W��[�z3A����譣dm@�iH�B�^�@��W���xV�ׯ��	FL���;v� Α_��m	Ҷq���]h*� P�EQ�ؿ�*���5�GGFd9�c{�-%����!qD P2��Q���<�� �����c=~8?B��dg=t�c/UM��j��b_�%��l9���:��U��.5[RՊ!�<�=���A	����z�ջ�Y-�zz��+�l���a!:�v�!�Zض}�[[��D P��H	�6�UAi#:�Y	ڢ)}�|�����������w������Q��յ�:9�ʹCuW��Z���P( �����{���3�べ	�@		ԭ�J�V�:�s�]U]9�:9�����>j�O�޿�1��:a�o{�+�5�|D=�uk�Ȇ+��W^~Q6o�Lo����������I9?xQ/6,�����*���{�t�
	c:��8��НqYcll*����ֶF�%<ԡ��ښ+��;9u�,��0�?��wl��� � 8`a�T���<+�vl7�@���(��D0XGE1���)�+��XT�
Ţ�9�&��O�@��n<�ܦ����n��4�"r���u����c}��_�mjX��ߜ��sTEsY,�b�� <@�9|������e�f�v� vzb\��� ^�p�t�w�;=j(\��_�0��X7x�F#�41���V_�7�|�s��v����3���3R�5�zC�#�����X�����K�p6 �:���)�Ҩ�^�:7���^�����I��ҘA$!p(��ܵ����脇�p_ax �a�#S*W�p��<�/�a,�r�&�����;,�_��]��{��ӀPC ����~��r��)���7Q;?��_HZ׷�i���OMZ=�k�J����U��S2��ܞn�T��IZ�+XwW�RuB�Θ�� �3.k�xV@xִ�ds���WvYŰ�#�����P�s�H����D��O*Un��-07mڤ�[c�6}�g��9۝'M�M��B�<r0�8!Z�h�bJ�nz�9zt �PR3I	�&;9>.c���.�u=��D+���3�5_L�=z��u�]�?��e6=� ��ad�?0�q����O?��y��2GS�NyT ����)������֮�H(�{�V�`5CܺF�`@.��$����MӖ��Ӽ�Nf#E��m�Ҳ3����hY�e76����\*�qi)ץu�e˓f�|�e�{�����|Xa{�;�j��H�"u����?b�׈H��7��U�H��z����p�xdbZA_�s��*!�&z���s�^�n�A::�L���K�Xa>�TO>��454Ȓ�Er�]w�����]���c|zTrE��A��PX��X��	:�e���
�A���8�2Θ�� �3.k���z�5�mz�ؼ�����IY��JpdAB�{�a)�eE��ÓKdR���-���祹�U�X�F~���dth�a�t�sySӮ7B��F��T�w<C�5���R�ݻwʖW_fi�q���ej|��%���b�*>OozӁ=������ܟ�w��ߙ�g�v������}�>Q�_
���ޱ�Y7�!���A��}�*�p��jx�(��u	q���a �`�|�����G�Ҫ�Cyd�M�38�~�f��Vێ^�%f�������ڶ��2y���=rۥb2����VJ��m�-�8�|��l[�j#���{���,K� .T4��(G�b�ӓ�j�i�����yr\�` B�9b�e�u��N�A?��]�.��r�g�ZH�X����i����Y��Z�� �u�Z�B*�<���� ����ݿ_"��4(V������z����gǩS'��e��^O4w ��>@w�e�?�G�L�M�����Jfe�����F�]8�*l�ȡ#L���'Z��.XgΞ�{�����<������7��/eK�
�F�kxRؐ�� ���ߵ�9�l6-˗,�?y��2��K�ϝ��۫/�(gO����s�9iQ����M��c��G,�JQ��V��<�����l߾���/�	\ ���+�6��+V��z\ ��dԻ}&���k���*�ͤ�좆^�F��4�@_�r%{��9}V�F��񇂨U��yp|D�y���6�@E#��9���^�SS�8P�}�-/�.=��ؠn<k&��#H[�x�����X� �K��MD��p�hXS����|&��a}�X����W�pC���-��7���E6�]'>oP��I>�ཎF�l����O�;Z���I���j���I��c.v����} 7����(#%=���6Bt���?r�dΛc��s���f������h��U��챣�w�^R�P����-wg��p ��5
���r��1�K�`��B�Bp�禨����;;�
>=�a幹�ر�D7�ǧ^�z{��p��Ҩ��}�2��g�'����N�#��=�<�Ub#%i�=��d/���1x�`7C'��Y=^���tn�����9�E�2���1�PW�l���i��uk֒$0D7r�P��ȇ�'�u�-��~�sy�/P�{�{d�;;d�+d��w�k4��Z\0�E���'��/+-�2����x} ��������z'ዝ��ġ
�����9x��C@C 9a�_G�(�ŭ>�`����TX����޷����P�~ ��ʥ_�G
�x����4^7�0w���5�A6�Y���Mgj�*�6�z��uk���|��x����M\���z�<zi)dg��9ǝw�)�]{���]������ؿO�ۺ��A�^>��o��sʥSr��1��#?�!# 3�i��;䆍��pE%RA���Q��(�[y�Y4�[��頑V�<7���~�3��?�}t*%q�3fy8���W���]���O�F%iROnB7��,�l�egk{��+yٶe���G?f/�x�ɐ�h��f��y�-Ң@t��7�Lk�sϲƺ���!X�����,b����Y&&�� pS4�`|X���;�HcS������;��ϔ�216IFu1S�B����\���dSY6F�E[,|2�?,[^MƧF��{n!�
a�B�Dm��x�Mb�:�TÔz���6پg����9q��/��<
>.	��;�o�Q\9�����D��U�^ü�9�C�D.�+��i�Vfw6S�]���9|�%�b�j��-����\�������P��:��@Oy]�2��2�׋v�Xs�o�7�� ��^�!��I҈bo�J�t�ӋDm?�=�� [����e�o�M�rQ �W�(�굫e��>��G?�4K1�џ�Q�λoD���1��������hD�#~�h�=�I���THJ,쑞��j�P!��b6%����٭�y��h�c�à�>�L�s�<+o��l��6W^���ݹ��p�)5\��O�u�m�D��{���/C1�?e�_������_G?�����Z{s����Y�;�C�
3�P��/�RMΜ>/�M���fj�SS�C�8uJ^��f��Y�[)��⛂ʾ~���F��_|i3ۀ��o�Ma��z�Vn����:Z�(���5 H0=�b4`���2=:"K�6*!w[��&�wO6��6<4��[�0��_��[_��]�5=="3�	��,�/驊�u~-�M��q |8c������%�ַ�Ź�MN��Y�X���X�IZ�i�C��A��!�kEJ���m&9�PLǹ�Q�	��04��;�8�MrkV#i���r��	��.��Q��F�q����}���(���9jz�%5�J�f��"4�6Kߝ���N5��Va�_w�q�<��R�y�L(���C`�K�b J��P���V�G^Zں�����j��)�J-�p�^���ѭ�n�ͩ�Q���;��<N��?VN˩矕9�]l�z��Y����l��!	�B�o�]Ϙ,��M�]��QkLFǓ29���'@	��ߤ�r��ϩCwƬНqYC�I�M�ԫ`�k�"GƸ��J99v�a +���@��F�
�1���f���c/n�,�v풡���,؜yX������^{���Y��r�8� ��w�̙��w�1�IN��]��^}EΝ:i�=�����ٓrap@�� S�iK65��Ç���U�#G�Gй��+��ڀ�-�\ ��.�0��|�JI�OJC�I�3�~�ٚ�
���|��:|V�z�t��@X��~��)b�y�!j�A�CFQ$c��	!ax�X+��1�پ�y0�qoи��1�Z~eOku1�c�rSs��R�C��"�A�AG	!S	b����N!��=�g���	ߠ�O�]���Ք�ԁ� a�������`�OLIGW�t��U��D:��x�ص�<���.j�g�Iz����:;�$�:()K������|6cڴ�T�ei(�r�����p@�ا��d� ��$s���u�񬍎����D�hK��G����@�|��U2��/V���b�g��p ��5j5O����*LZ��E�;�^eB���+�Ƹ���d!'�S�H���������jx����zex��=��#���oYܐ��,y���?8d�Lj.n��Ĕ~��@,�\Ȳ}�ӧ�5�0(+8�����'��\(IG���c��'?�II��d�O������YE���42|������V����y��Q��\�TM_v�r�$4p���m�Q�ӗ?k���b�3G�m��]D�^z�N>����ф�6IfPB<�c]���=G�+\��+<j����YW�ϫ5��E����cP��T6Z����C�%���
�Q,�:��e0��:�ވL��\B�B�!qz&�:}h@`�_�aD^���Xy}��d&ůbE� ��ћZ;$m�g/��B�J�G����
!-�g�|��(��NA����4Xc��YJyx~kV����LS��Eio�g�\���\�������Exs�ϕx*-�3����Θ��<Tθ�ᮺ�!�m?0�pB��R�>�J����.���mP@-���z(��K�gx���Vj���6eEy�g�C�fdD���� \!�
���C�m�jHLz\tR�&g���7�BZ�S����K���N�2_���z�Jy�������"z���0�|���k�r�� ����?{��� ��P��J�f���������{�Vm@a,!�mj.z���M+S#/�28?*>�߱6��QP���AH�|���9�s�iߚ��z�~����'h�F�t����UTjYS�&k�%r�v;R��i�B�9tIC2����V��hب�r4Dp/��g�$���8Ӊ$���J$��s�xP*��J�>��у����||bFZZ3$G˺�#�J���ΆpI����m�55�������8��"44 hP����T^�ѸLM�p^���Ѩ ��A�m�R@�a&�����g��p ��5���ڞ�-P/ �d�{:�e@�0�y _�z���T���?ۊf�l/ g�4S�@5�ӼUO��y�W�\Z��-���[�����d߅7mlb8��z�J�E;�z�7�ɫ[����
y�������$����麼r��1����Y�a���eV	Y�bt�1pM�9C^ZǺ-�t��+�z/q�cX||��ҵj�3�Y�:A$��(�-�
�������wWM�x /�z�1��\�m]i��'M�R)U���I"j� ]�8����_Q��#;�����^��Co��!2��bN N"�12R���h�À��h�� ?����EA����*qK����{&{F6����Z�B?����ʾ����ǳc���Ĕ^O��-�cײ�
{x��sc^�D��#��s�Z���8��7_=��nV��Z]�(/Ԋ��8��=@w�e��ˋ�$���f#tk�a^2o6P}��<5������P��eB솽��lR=/�ϼ���@���	F���Yb�x�-�':<���o�����-<� ����W^�w��utʃ~�y�ޅ}ra`T^{�m����������W�#.+���ٙ��c�!��a�*C�0���+�j$�O|G[��^��Y��E�<�~��a+��J%��u����k���=���t}$ǎ�0�Ǭ�1r� ��� %mCÃT�[�r����q{������C� W̩�����^�~�ZA@��.���tnj��t2Ź�x�A~Q�����G���AF���H�s�(��/����? �O�����Fr۞w�Ikk;�56g�����t!����U�>��8x萬_���I�c�������*ql�����Fԥ���n�i1��B�ҽ����O�Ղ�]�P#D��g�tJ��\�7�Τ��F�I$��Q�Egf���
��#��Y�;��%&�R!��݆BȺb��Z;'�2��PU%� CO0�fHPs�;6�A�JZ��b�O/
L�h��r[���Vq\��R�`���O�00h��rE2�AV:~��O��:���yw�N�{�B$ �b)Os~�z��}�^���8�%=���,/�?#˗/�?��g$�����u���.�~�z]V�:��)�MY^}�U6��F;$�@��I&Mj� �	qv�3����������z�Q���e	X�h���3g��c�=&����}�s��ŀי�Mz��#��d�T|�8K ���ǖ�h�SP���t�,�PeCi��|�75r��1�|���� ��5:rX��A�� ۋu
�x؏�b�S8c��VԐ;�^=Z�"J3��CS���op*֮�B�9��> ͭ-�>��z�X�˻=�Hͥҵ6���HsS��� �[���=_�P��̈�lѨ%���(�w�3fy8�������"���<)6\ts����z�PR� ���s��T/�����{x���PSl@�l��G���)�d,Ƽb�����FY�`�l~�wK;�<CQ7 s n��m3���u��h8���_�~v�Q4`c����c�v�b=z�^[����^OKs�tv�K.�d�Y�/�e.6idnD�ɩq�ó�I&f�y��a���nz�<��0y�򞸌���<���C�Xc��7���Y���'��������J��ax̙;�k�χ��4�W*��VȨ�65�������?7=]�̤�d��\�qN8am=<w\_D019%?�����½�dSF����I���l���O��܂��4Z��nnl�y�L�N�-��"�T�����Iޫ�I]��ٳK�y��k����ha�L[����x+W%������yz+�z
��O����Ӹ|���d��>��N����\83$'��1��djbL�݀+��3�1��tg\�p�Vjހ��I8�W�H�¾$�asY!wxX3�=�@�O7�h�B&M	���O�я�sU�r�W^y�l߶� �Ps �{ݾ0lmv �ݤ@���l__	g� �A�aB�ؠ�z�)�) 7�t�}|�}�3���˦�Ix��\��nqy�y��P��:u���ŗ_V�4]�i|�_�x1%I���N���(��5aH>���ay[(Ŀ�Τ,���p�|��wf����j�y���[����G�w}^�F��?s��&&��7[���W^�����N�߸�s��b�2��-��� �L���V�c�؆�6"*z2�����G�;�k fCe%c�A�����TD�����ͳ�6? �!���C���z�)�a�w��>19&6\-Ξ�4pS�A�ZL���v��L�����S#���=����0�	׈u,dff��-����4��C�Ի�zd��+dٲ��s�.�pJ�VTTj�C�sƬНqY��������b���Ke��^n��희Î�ǌ�����uG�0�7����h�2���;r�7�|�<�����A��׿�Z�������X����l/^5�8������6�<�zG�Ǥ
�r0��3 ��ƙ�-U\?�ؔM>:_'H�}�����Fz�6����jJ�u�M������a���XБI����Ҩ@���f���"˗-����Ĥ]�@�5�z��eͪ��m�v�g�D�� p#��G��O�9a�Ǜ��Rqk���Xߓ�����˰)�	����KMX_�[��_�ͣ+1�W	�j�)��øh��k��V���zc8�M:)6xa��<K�P���~�S5_�[BM� Ϋ��W��R���%���}9�RQZ�%�����!)B�U�������!����QJ�b�Xa`Eh�.��
�R�\�ׅ���O<����F�n�:IL�3��=�WZ��ok�KwG'9P̧�WO>��[Q�U+���g��p ��=��ZW�o,� k֮�W��=W��E,Q��������g��_��I	�ƌ�Y B�h`�S���X�Ȇ�U��ޕ#��u��i�b�U��bsF}5<���i���?�@���" ���F��y��[.&�T�G��[2�׹/����bȭ���R�a�o!�[�ȥ$��0������祩��Q�4H����k�1��L��QH46�d`pH���]�Z�z,r��Y�!>��1@�o�.pm �h1\�����A���]	��5����Qo?�B!�u��n�ugn��7�w\�y���A��)��>?�C�4Zۚ���
v @��f�����
~��`����4���6��.[İ�a�=.��LN&H�ǔ���?�3�=$������[Z���MNN�: B<c�VN=�{;>9�{A	��#��n+�M�9��g�� �hX׼���$�p�A�M��"PO!��("����}���}���Je��>@w�e��[�-@�</^A�r�Ku����6�� "�
,k�.^Ȑ��mS��x�Q��FV�gZ����+$�����ɓW|T\cx����EӮ4�75�.0t|�n�SgN�=��fY�h����+����i�([�X.�)�X�A��;��zz����!��!{Օ��1�=����;v`:���Eϱ��p`z#� w������tx�1>��ѣ��p�T��#�n���r2 >�<6;�QXŴ�@����T� }塺��& 34@Q�A�@=p��!}����bۣ���nT���=�A��Ax��l���m�4^j�t�Lb�������o�-�S��X� �
�Hp<_��:r��A� ���c�� ����G��D�P����Ul�g����HVDy�)5����: ��&,z-A=/�	�Wt�1����-YL����C4��o~�r��!�5D��I8r�,\��u�'Ύ��%�d�|?�b.�ӯJHL��v��g�Ru ��>@w�eݜ��pDA݈� �A�6���V�Y!ﾻ���m��N��<Tض����;r �a�DX��/��6ѫı�Ի��I4$�#�^��%S��wSc �/*�u���?OC���M>�˕�V��]�V7 q:��k��F6n�J=�݈�V��׾�m@�rɆcq	��A�F8 �ӗ*F�n*�Uc��G����-�ǰ`���nv%��
�)�HF����q�hz��cE��D$\U��o�,0@0_C��a<�4�K�c7J�`< c
`
�������jx��Mc�
z�p�霑{i�l��B�$3�ƒE�h�����w�ex�i����l�5�5�7Q��4�0$v�e8Px����w�X�]��cg��a���Bc�o-�x�HU ��*�BIz���|�K�z�j��?��<��/䪫��_��_���ݗe|t����II�
��Ц��?|\�z����h�o��t�z�xY�Nٚ3f}8��� t��k�4����D "xq+W�R��j��#��N�ܪ�I�Q=#��'Ƨ��}���M���J'���qCf4���Q���¥ 'x�^��fL��
K�Իs{�?�:��+lk���w���ݗ���.C��.�o�\}��*A���	�Za����ѣǥ��C����$�.R�ή���Ъ�8�k�8B��<�bހ4ś���'��;-�t��(P��hmc�z&�p~R��!BcZ���i �!����T���sF��Ng x��&8g[.�ܹRRO������$�麝<y\�8ɰ���Ar���a  ߝ��Xߤ�a���S�%�f2��c�#�FA$d�\�_��6�~�g�
�yMN��#��,s��{܌d ׍�?"3�z�(��1�c�E�� u�tV��GY?��;���QZY"I��J�͐���E���q�,���R*�׾�5ӗ>2�m�5}��9[����7�J�V��N2�������8��������8��<@w�e���S�l&$J�\�^C�����9󥣳EQC<���,
�#C���ƍ������#^����>�Yٶm+�Λ+��x��h[��O�v�2B�G�!pa`c�j ���pCj(x|a�g�y/Y����� ���d篹j���g��FQ<���r���w�PTV�^+��P4����"�\?���1�<�q y�d�U��8F�-۶���� �� �u��yF�� =��ّ�\����z~УG�4:��\�����$������\7�K���|o:����c�� ���:�5��0��ZR�@��`�p9��B����N�Y��WW�#	B9�����>�f:��W�(�~��"8�ĭO��k�
�R�~l��Vm�K�1�I���;֮Wj���"����!��7�E��'>x��ş��Ϲ3��w���FR���j��L����|Q��w�j<554sݪE	�erb��Q���*����Y�C���j�]�V]�\���M���QC]t�ԥ��>�
�Q�
���<==��R��kЯ�5ҡ^zR�h��������뮕��?�e\����.6g��dF���M2���l:�Z%���M��w���9))p�J5	E��sK���I�"���D�U�0� �t�2i�鐪�n�S/_N��6�bq��e�V)@>/���ꥡugH�=��ib�������z�:O��\�: u�w�!
�cht��bnoP���%�w�d�].��`I����	J�S%���:o�����^(KC�`���\�Meh �cX��Wl~�;*J���'����3B�%*�!ڂyn��WB�|��=z��/W�:k��P�C�����W�:z��]�
�^�\�ϥ�Qq�%�����
�>��$�k�&zm>o��P�I%f�U��$�t��5�Y#7��J�Z��t=������|�������� 2`�]�&dIo�L���gd:]��3%��-����	�����4�\O�{��>�wP7t�.g�uƬ�r�e����&]45��8
KҮ)2��Pegws�h�q��9�3��0K�ʬ����?/7�t����.ϰgË7*byؼa,����O���Nom
J������x�T{뭷$����+����GY'�����E��w�/-�m2>5�s�0���><�	ݘ��n�	��JE�j��˟�#�O˻���t��ԩ��ͦ�l�Y`H7�^sE�y�@�lw���� �I����
G���(�F9T�`���`�S��{��:P�C(dE��ff:������X����� ��$�)2��9��]'��C�(�7o3�a�� �z�р�Ü���#�.��5���*����(��e�2��d��ˆ��T��*#�z�{<�<:�s{~�$�Jyv�Ct����@%QB}:� ���'������[}a�D>�	Eb�[���ko�"}KW�ј�u����ys��!ʒE��&Ϟ��[������+��3�1��tg\��U��]C^����X�d1�~e.��{ɒ������1��7�i¶��� Ȫg<|qP����ˇ>�a�����{�Uo�,�����i��Ƹ䭾�v��T����  ���ǎq�G�Њջ�[Ǐ�Q����ѻ#�d믾J:�c���%�<�$�b��4Q���$��ꁖ*e��3w�;~����/X���\�rH�f��`��
���p,h��E����c� F��N��2r�YS	��EA�EI�F�Tҧ^�b���4�IΤI"��� ��� �5�~`�27� Xd����]���װ���.mv��Я�|,��4�m��
Yۚ�l��M�)W�/~����kl���ԥW�0�ۊd�g�M_s�9�s����;R��"~L;W��-�y#����a����0�mT�00ix�QB���:z}g�Lʊ����&5���[7�ƍW�!�2��ӢF]Z���{���Q����1��tg\����%��P�#?	� Z��5�Pr����N>zw�>����O�{�~��������ٴy���{�����m!�%\�3Gn����h��kW���3�:���/������-}�����d����<���{�r#O�\)We��

��M�����#�׮��n�M�~�m�5� �X�A��V�����>���K%�]�v�"���[dx�";o�����	��3���2?�%��5�����<]��?Dxة.�c�d�ɩ��* �	 ~��En�r8��X'�z���܆z�^��U+�����'k\�(���H2x�L �:�B�`��!���Σ^��ظ	��B��j�?�!���f!��j�j1���v��j���k0�pm���w;�O��%�m8��.I����ހ}n�k�����i�n�+r��7��U���O�a�G���i���5���[280.�-���2w�G���>@w�e��[��C�Uÿ�|QF�'�#I�3M(�T` �p��Q���b�A7K°9�ܹ����0�`����V X�7T�%�fL	�D�!O<�HF>�xIo@=s�S���g�����!Vȳ��f)i��l�P'S�06�������3�.��}˂�>�8�>���6�w�X��㨿���wv(0o ���F��z�'^(f��s�.+̍kR��9O��_�����8�U7�1�$�)m�d�2�1r�,زek�)�DbjX-�Aq��'�i��6b48~l#4 P�=X?��Y�N1W	#z�b�r�dHd�M[Ey�HoV#�_���g�F�ǘ��1aT��7��F��Vo�4Tnk��J5��m�� <�[����o{ܶ�o�6"D�\�r�M��U����zw;t	��������V�����_�������TcpP�zk�^_B&Ʋz�sd���F�O���S'�:O�8��<@w�e�j��Η�UR��6Y�/�"�1�3��t�p�_xu N��St�B�0X�]m��Wc��K뱃l1Z��� j4q�����p�q ������ϙ���e5��1&���a��m�t��e�8�	���~���6[��0J(b��B���ak�毠����O<�24�@<f)��x$Jp�d����:v��jh���e�>�}��-v5�b���d>�w�^��� ׎c@�^;�dP���B�_��Zy\������cتr8�i��#��{+
��;�]��ikm�@"h܂h�k֒<�셳�p�f�ղg�Nٰa�t�wpN~5�@8�:@�@PY�Oۺϕ�a��!�Ӹ���k�@��+60��z�� �F[]<�U�N����#'�q`��M��}N�E����^Lȡ�G-�9�tu.�p�QΫѵf�:)�^ĳ�
G����Y�C���	ּo���7�j�k�`���t��;��

¨͞�������6@l��4��2�ө�E��ՠ������qk�ѲQ�����E�BH�D;��3��y���y(��@�.�E��	�Z�(�e �B��p8HOӉ��/��.�{�"�����W���9'T[�҉#�:��������5֟�����%#$�ɦ9�ֆ�L��%VŴ�9�.4QN���ĲjU]UI��;��0b*=�R�e`h��Ćf2��^���0Akk��m���y��M{\v��q~z�(��䡇����I!����Foz5rzΓt��<4�+ղ�}��������Ǐ=J��m0�Xyz���w�2��C>��!�C��n����˙α������������A�J�Ҵv(^�����/�� +Z{��F�F��IiR㳩є�-�c���,i��|<.�W"����Ę��:cև�P9㲆��/z��*9Z�b}3�=%�xF�eF�D�L����f�s4"��R"�VY?���wv�R�D������ɏ�7��[���4�]l���/�H���&��(�I�G=|ݵpdH)F�V�Ur��sVϮV%���H��r��iy���h��C��QS������!�d:#7�|�D�����>*{v�2�`:%!5�ȵj~���<�q�_�1K�9������ԣ���1z�K�>F���PBC=:��m�\ ˶����i��7�e�M����H�K���T������#����6�-��wv�!Y�l�s�eR�3w�,[�B~�O�C`�\�"D��!��N��y�5�kG���-/�K�#���0�M��C�&Oo���/@���]�Z��c��ư�8�M3��������Ź��VYлPj^��5S��\���ɡ;cև�θ�Q�T+�`��e��e�6]T�{H,]���5z�~��jV��*�i��E��<�e�,zl�d��o����#��&�����>Bڨ�P!�ja�y�{�lo	�	cr��B)�fL����B��wn���un!�W��m��{�;�3�ʙS�����r��Aӵ�S��s:���S�+ɲ=x�W]�^N?Be8�E/�ڙ7��
������Rބ��U���M{Q�qW�*�r��>��an�C��DbF�� �� ՠ�	���V��s��JpwAaMLA��~�'�K��wY�A�������s��R)�0T�a��9�cr\߃����w�p��^��O�'s���<!sj7�{0 U��`��g"Fji��b��b��mF>�cs�����s���G�1N�8I��ھ�-9]�I��ʢ��e�6�
Uz�e�4>jz���7�LHCK��kB� N#
Fk tX�Θ�� �3.k�Þ�z�U4a���0��Xfki��52���Xm(���P.=3��X,W)���5�GGFXN�M�56nl�)�[��޴B�x�l{m�mϚ6��i��u0�&�}M�Y��z��}=�qr*!}����>)�<��__�=_�5�jL��2tq@̟�y��W^u�T�>��5�����r�y�ͭ�iW,o��j�3���0�67ĥ%e�8��C��R���5M�$�z�h �F-ȹ���Y�F����y��/���L�\'`�#�B"�r�6������έnh����+$�k����X4,������{4G�y�o~�_���}�Ш ^q�����@�z�86�WK�:���(=�߶��c�+�|�[� ��,#�J!�M��K�l�����鹙*����Ƅ�0�c� �Wb��>gtv<l�Jp�$������?��_��5��LG��`JB��Y�;㲆n��b)_�����eX~Wp��������p��7c���%�+>��O�}�c�°��V�y��ʮ];M����k�GM^=�Z~V�)����;c}  O���O
�T��K���d\���{�֌��z�P�V��(��6m�$ǎ���(>�A8����t�����E� �h��|���1G��m��>*�ny]V�\.�����[��6F
��*�6z�{Exa_[����Sr��YY�j���_���ܱ]^z�%���e��>��߽{���_�9Y�[��̒�/~�"x�<p��q�m�ax=��Gu�?#��.�/}�o����?�������&�Biki%B�'�MS���>�!�3<������Oפ!����0�>$�x��F�t��Y1i)��q;��W��.�iG77<x �����{"2R���9�>���}�����r�R�ÇL.�(ĳSRC4�b1�צϻ�"-m~�W�)�̵LO�HM={�'@�hmm��3�1��tg\�Ѝ����k�LIR��|.���y"��W���wx\%��%B��x�O���{eמ}d��ܸq���_A��{F~��sRIE�4y�p�['j������m�������x=~�˖��0$��nɌ�Λ���o�믿Nֺݛ�z0����~*3��`w�v���rZ�/�e����b�\��!���p��iiX�TV)��)@���wG���jS�c=:�4˧>�)Y��m���򋛙{�xݵ
��Ɂ��exlTV�XF��/�KXo����P2���<p���|�Jg,\��=�m���z�0�Э����Z�[��j������ � w��9xh��]}���j��0�^<�v::ۨ>7�w���G%A(������zo�jƸ��6H{�G����3U�3iЊ~`\Z�v���燞�Ǌ�gHA���M�{����̥�
�3�Ȼ��䆛6Ȝ�m�S����d߾29�������.*�TN����;㲆n���n�C�<���|�ᐴ�w�KC.`��Kl���a}3��[�IO��(,�ƿ|��<<����o��%�����_�Zrټ���YU 24�AL�����Gk&��2�U ,� ěP��n9��X��" rl���sH���I�,Q_��������^xAF�%����1��̨/(���ˆ�{<�2��=��_ɉS��z�U�~/�N*~2!�Bt�C�B�v�.)J� �?~�19r𐴨{���~*o��]���,[�\�y�Yٳ�]���
�y��4eh�����~�3�(+����}^��47�����S`Nw��u�+����nr֍$�<r��o+��5��aL��_yg2)��ڍ���?�w����{���M�|�R�Qo�o�4رіz��H��/=�v4;�D��Sϓ���1���d8��n�j�����<��J����/B�_�z�H} ���y�5�Γ�߲Q"!F*�Z��OP��W�����d�oȡç�]S��T��i����;�F*Uf���y��x�sϽw @.�$/��ի)^�<���
<��c�Y��ںuW�=���\�Z�����KOwER*d5� �1��H�^� x��������O����3)c��Ӎ%f��F�yao���d*9i��f)��)��������:Ϥ\8wJ���v6��X�� ������L���G��Em�{�
�\&C� ��fG�!�W�K�у�u�#F�U�����9TCc��oIT����E��*��k���a����Y5�^���x�0�ʛ� ^=�~C��h��O ���lJ㬼3�$�M�z�Ly�p����u�"�䔰�y�ݻ��^ܷP��d��^r�,�3�ِ��k�;�>M �q]�sf{����V�n�cwC���y��Y����-�������,t.Q�����Ck?��Q��K$�u�WȠ�e�\A���F�/}4�pKE�Ʌ�;o�{5"S1
���I�9��4@w�e�_�z@�&	�խ��*7�t#7`�����G�SU���/�;'O������}���y�����W%o�7�|S��:-��q��K�7<-���"��V�f����e{f��H
{a�f*��n�d��1,
F}(@�w_�b(��,�Պ��aX����/?��Od��iY0�KƖ,���]�l�P�D*+C�3����r��=�Ikx��-P+s�q��9��@�V�v���C^W/���^�[_G'�� �p�@��G�4��w�gr�h�S��'L8��B^�PG�oQ
 �K
F/�7;��ܱ�TxSo�̀ȿ�;˜6^�Q1��=�@<��W�{n�����@���[�&]���k,-u;��zצD��{��6��w�(h�a\��\��`M���X�xS��.\�F�J��}{��=`Ń>C�<2_���5��'+֮�e�7�=�Kjʆ�	4��@"�Fٰ~�<��k�͋K���Y�;㲆_w�x,��ʮ����޻��ȑ��S��\������&����n�W_�b��k���#k��@�ح
s�tˁ�����������v6�v��&���D����ٟ�M7�O~��'B�_��$� ����QA���}������BA��Rc9�|�V����v�����r��~��4 GELj!�`��$s%5z����HC� ��Ks<F �)xN+�������m�s\Kj��k�$@��U�`A�e^�L��k�Yy=V;�
��C$b� p�{��I��ŏ<��g�QCo�U�Y�gSs�t(�
"죞ҹ!��Ⱦ/87�-0n�f��0�(w��M�2x���������{�T�!�����O�(��.{��*T��\��۞4�v�C��Z�ҹ�zVc�,B���V�U��@�#	�J���,���'eѢ^9y�ϵ�ͭr�m���7_����'�Ҹ�6�$W��Z�~�$�)��C�����>��"��� �m�H�Rg8c���θ���֯Y��xV::��ƛ6�&�I21-�(�.���m�0���.6 9w�<ʯeيE�}Db���P�mX�<1:y}�_�%�>���<�Fy��ڼ��u��b���,�\.�� �|�f2���V�x#���Ш"W�Y!?��I�cA����s�9�f�Ź��Fjڹ9��._�ܘ���gN��b�h��Q�n�O>�aI�����o%��P궢��w�N����s�S��������ab�C� ��ym�� ���I��xh�y����Ĩ��J�b�+�,Uc!F �p�<P��ܠV�~�b"�(+0����9o|�����y?��!�{��A�<zo=�ˤ�����X�r�dR3�7�#�2��h��׀05����u�a@��aɦ����ȧ��0Mc"�Ͱd�
����#�߇dp�T0޲����f�����4���6��q#��<�^������R�{�h����$���l$s�ܠ����ge��9�W��|�e�+/�H�H����I|�ؖϱnjj��Ũ���(�z�b�2~�=��&�?��8��=@w�e�����������^��t��IbfJ�ᘑ����	o�Q�e$��4O��"�0�W���/Js{��\�Z��>2��ы\AmA�؆�v�Bĳ����t��m2��@��C��)�R
�n�[E�,o�<5�Q��l�a xtn ǡ�L&W � 4���ʊU�e�w��[��'�T�K1�����>�~�[��L�wv�Թ������N�W�k�N�X�z&\��W�k5!g��b�z� �a� �⑃l�&(+�W���&�����#۷�u�֑�p��Q�����`H)���5V ص��9�������g� �g���O��C��Ģq�������A�� Z�*#�p׽d:&ށ�ё�_��g�����7��*Sj��TC	�����=PC'�1�����G)m��g�R���q�`�Xf���:�1�a��1\ ,T)������ b�[ ���8.����u������oB�B�X2�%�`�/o
����[n��'ϐG�l��L�X�sjX�K�W��)<g8c�������=on�Mw:��cS�T��4��xز�v[Kx����
fy���%�V��w�-�ջ<z���w�_9w���d��FF�5�v�n�Pݵ:� ������3Tߨ�����u%��0y۠����@�`s����ǈ�$SP�cI�#�<"��1Y0�[���Z���eNW+��ăz=SE</7^'7^�����k�ʲ�YK��ȡ=�$=5� �gLo�*�	�lR)2�M��Z=dl���M�H�g�x� ����X}ק���C��6�e�t������ �-�]�X�f�c����Ő<���\��{��["�����)������	�s�.9p@�ٹ��AG�'�C�<��I�5�XN�05���{�C��T����ǚ�؀PPY�n�/@�D �eS���#��#��J⭺� ��Q.,�|��Ft5�RΔ�!o_(����C34�����}�3ʴ�ٿo����ԼR*�dF�Ά������=�T� ���i��|�@����Θ�� �3.k�s96[l�`\C�-GM�*7��d޼yl��:�r�"n���t�iǈ�l|���7�%����K���?�q)��֛o�K�~+i�[2�5j^h�R���y����Q�<22"�#��9���s�yZv����Jz�K���5�0��G�"%���4<����*�4��d��H�gY�C��OJ�+���ѧ3yʯ��;���+8�ڿ�e��259�P9J�pL�����Any���o~��R1��($��a����R��F�M\����=���1D<�%g��y���kX������Yϸ����C}�!qpVyױ'�n����\-#��U*�t�����Ŵ���w��E�L3}��w��_H�ټ�L- ��^��JI$g��N��`H�iF:������`7���n����G �_Z����^���^S(��x�} �ُ'�\��}D�wӍ�r�
�eSlV362D=����=������z���ǖ7���i�W_-mme\���^��{�� U�kf&g8c�������n������|��J~࢜:}L:$��t����L� �ʎ���[���?s�]� �N�>-�?���ww1	ŭp�4� �&;\�!�����
�+�R��!^�O|��-o��ߒH0 s��]ާ�)O�+s�/�����h���0�}�����!�\�|�3˖�7IWO7��Ȑf0�$���̤�6=�������;��Y�&�(po yW�5/ds�˟�B��ͼ6���m�~�ht���p��{ǎ�A����W��3N��11>���s���w�
+�v�U=�Tvܰ��������>����dǎw� {��)������Y�=,{��}�XQ���%�^9T ��e�P�;:i���1�l�Z�Y���g��|��7�{X�4i��&�`������/�� SO����j_�H�V�$�h��4���|xI� ��n��&��׿��6 �|	Z�Ui�k:���8y\�u�X��`�A<'�׃�Ap	p߻�:؏Ǉ�_ϜN�����Q��y=��d��ݲg�.rR��+5�v�֜1��tg\�ЍХ��ʠ��n�F��O�_���Uoo5�2 �0:�)h@�t`p��Ml�� q	�P �����Y�U��)z���2Z�rSL�p$fB�"�%��u��w�QcC�p�45Fd��U�J���6���X=�B�K/����!�b��m����n�������
����%u>)�T 1^)�;������o2��S��"aK���w�)�c+��{۶m��c�T��z&�� p��=�JXq- nD$�<�6miޏ��կ��8G� ��K���в[��0��x�<�-��50
 �E_t|���ԎG���`��ut\{��g���S�6��u��7�,+W.gy�w�&/��U��|��E�ʡ�G(:d7T�yC��������%�M�s��l"�y�:w�������ܸ��D����Jkg���_��\�f��ՠ7��#8L��y��F��ׯ�F���8� i`Sx��dD�A̵�o��9{Zn��6����YP�U����Z��g���F���d�����g��p ���M޳�k��yA�9���%}��X-5��g���lS���	z����k�0�O|�S�G.udl�x�
�k��G�������R�W��J�!*T#�{���!�=��S��sϨ�:.{׫�TU�uX���;�9oeۙS'�?�����.�7J���<�� L������Бc
,
~!�	�Jd�����H��Eɪg_ �/ ���R��eٚu��k[���%ndsA^����уE�n���@�OܖsE����ҧv����Z�Z�ה�.}(�G��l5�
>0����G��� .v��Č��'>)���y��W�駟2�
p�hL:;�����$�L$/�u�]�HK�0qm��VAGwk�C��lg�mOQmp��QiWP}��-FI�X�����=8���̛�D�+��f���+�9�
L*�S ���q9!W��F��5B
��z�\�B�B�`���T�X�*�"P�tRc�!q"܎��M��ٯVae�jAr���R��c����C|�Ϟ?����T�Xɻ�����:cև�P9�2�Dx��wn�ݏ�#<�b�B��g�k]�t��u�]r��A�;q�@����=s�'t ����`�o��d��(������)����R���8'<�r�L�yaS�l��(�
U�̋��zޭ-MrH����=(��88u��^D��,�h��� ���!�� �J�۠_�=CO�����D�j���Y5��iw�\
輽}'��J�4�)"iK��{�[n����O�d��>�;���p(���k�;�Z!m��h5�l�u�v��Y����(�\�]	�0(�b.��H�5����:�5�'z��P��_�<��+���&��IvE�cG��7���/�~�̙3��3�ú��\,��� �x��u��m-2��[����q�d�5���|��߰�J!'F�h,�,.��2���޹�c�����/�� ���O�q�~�����rT,mF� ���&I����ѮUǽƺ�9���_�����F<Ͽ�I�ီ�\2���:�F"�gq_�듸^���&&��g��p ��>9�������W 
�t�Z!uy��y��7į�,<�Qݼ1���/���瘫���kY.�M|NOK��~k�{�1l 8����b���u��r�i �z����=��fHb�� W�X7��~���կ���՛��6ƃ��� :��D�!&]��r�1��Qҩ ����/��sd��j���@y����/��oB�`����?�R3���=�̽��P/� (D D��6���-a�;u�aDẰN��Gc�iDJp,|��ۃ� O�̔ J��\g��5�&C���G�S�%�$z�.�/�Kj�m��������:��PB�uY�;_�X�JΝ>Ŋ�^������3
.EB����d��"���q�s0���u���޾^����$��[m��]5I}�y��	�:��'��M͊���+�TϫTK�w�z�(�@*���ıc\+�� �	^$��{b�iv��5�:��OI�ܪ��>��\��7*�p�,Н��D�����"F��jaZ���gw��t����5`�zM	6���O�k
B~��r��w���0ˆFG��ȡCd�{����v��U$LX���7CѮ��'vKA7gl�02�/곛c��,_>� �2%�zy�lδNU�Ĭ�xc�='��b�������Zs����?v���ٽ[bQ�e��}�A��'>I��_<��Və)����g˥�a��P`�����na6���g�l��;<o���>�W̍����q+ꁿ�/Z�"k׮eH �(
r�۷o����T�E�+ZZ�EFp�s��rM�F`������Rմ#u���񐆩+���<>�u���+�-��O�8�m��-:�$�l~����>b�)��2��=��IY?;2ԯ���czF�&�$�7�sE�{.��j�r�暫��ֲ_�_�L�p$���b����L����µ㳈�@����5�$�������[��lI�nD��eB���#a�֕��8��<@w�<���m������ۅ>�U�k\�y?EI\�n�eZ�����L�8�U@`B��������{��uUYûr��I�n�eɒe�9`l���`Hü�`0����<�,g[�eY��d+�V�s������k�{K�������u��#��ֽ��{}�k�}�]w�S��k�Z�'g�yw?��%y=�@4�O���ܠE
�2Ӝ%R��n�Q�c�A�L��2:�G}T�%�޷�>�f5���B�.�gf��'���6�0�m'����eL�THI��$�}ۖM�{(4��{�	z)	��n"a��i��o�s��S����2j1�0��Q�x�~�/�6���ODJ��tʮ�;�ְ;XǴ6љ$�!ώdv�T\ V��O|���~B����S�`v�g�2E�<ET
А�/�,��<�><���Voˠ{_!�nvM���y=$��Q���pe����*"5z?�O����^3������ �JU�-nOI�[t��!���T���ԲP�t���Z��-"&� b��ky��GG�u^+�(�gKL�p�����싞/@� �vY�'p�-��8���Eb��5�z��*��]�f6HT�-F�����	�,-�j�����L(6Px�Ua􉞐'{\�l��R�t2��l°����𧪛�l5R����+�"֯�X��je�QO=GO3�HK":������N���Rp�#ǎ����us���)��l�Z�b���q�Lim�l)�S�D�eQ����"A��@�Թ�i�Ȝ!-䬲1c� x� ux�X�@�S��k7uA�>|�A^;��o#_�� �Q�kȚ�a�>r� ~<x�o���epȧ�K�1 �R)�ﰥ�^����w0
�`���O�]М�r�r�n��=�K�`E"a�	sC�F��D'���G��V>�I�	�Ct�+�L{�ۅ�.ϙnm�DG�$�>����j����+7nA:%���ͤ(	�7�ms�p����~p̐��ŏbC�LaP�AZT���˦i�D"!�l�ю�~L6�~�BB(�#�:��8��q.#?{�̑l>�VhpB���1�R�d$>tcv�鈅�ᙣ3��� 
�7���kEh=�`�P���t�6.ʋ��B��i���/\OX,X��0��Eo�+��� ���	|�Rѡ�T����G]���Oʴ�3��e���M����9��T�z�%݌�0B�{ۤ�]�vI���g����m��+�G�c��n�')F�Mp@�޳]���Z��m�����$��8 z�`��| $�y>�n$����  H�O?�s �p ��t�ʕ+	�&�>*_��ef=�}e�+�O��a� R��C"#״Y�XS����F�����M� ������>0���%S��H�9V��'��������KVn��J�٫��(�D|��p�`�$&s�;�F��髧k�LC�(��z���Ri��~�����4�����I[��cj���>A����\އ�A�������>}�NJ��|H?��Wy�Ϭ��$�qA��d�.���8ϣ�q.�s�T�4����b=N��8�%�#��^ج��+7�B� A�V��}�$|� C��"l����[ ���xM�9��_�e]��ZV��[�!����������������Y+�p|k�T�G�)�R/�k�e(�s���Co����M�T(tB���eos����|�?'t���K��T��;�BUR�^֥Zω\=��Cx��=����+���f���g��rH�34T���n�aD@�w��۷G�,Y��8tŃk���rm�-����&�_K�"r�0 X�U(�ۑ�����ҙ��&��!R��b�Zu�`�O&R������i��9*sg_ǢDx��kU�w�p�,]vǞ3ݒ�Ee|dX6oݬ���/�Y�UX��c�>��9Sϳy�f�2:���0fUT ���w}7��[[��3�c�]���WK!����TC�|�Bd�E5*Bj���h�@�ʨ��<*�^oLNV�ٷo�n�N[V�X9����cμdm��h9��(�ۆ���p�d&k�OvEcW0s<�|�E6��4y���EP�3?Fƴ*����AX��XW�^?��m�ن��ͯI:>���
Ѣ)��_M��Bո7 ��v��4�H��P��4�g����'���́�9�7�c]rΡ��Ǥ��2��������k�����&�d��L�P0�Q1��ZBM�^��'Ήc�����ڭMqN�<�9s���0�m�}46�C����%��}�&9t��x������5�MY�;�і)����:TE̚���
�Q�&������-�W|�薭�@԰:��ͦ'h'��N[��r��1MV�]�p��Y�إ���7�@둅��)��V�G<z?�̤��g��iҫy���ǧ�^8�Fޤd�x���XF��^ ����yM��Ӵ��zC <�G�_�X]�9��e���<�d����#r��Iٽ��?tR��\L�8K��TFe��Q��x�c,����j�EmYV��OV9��)�m��DdJK+7�޾n�z�)��F=0ژf���K��<���w��V��@BH�f��dZ�z� C�6�\;dlx�z�5��r��tv�SZ�*(��!�x��1w����ߣk*���,MO��}~xm>�ݩ̐�.�`�$���2ۮ���ק9���wC
�bz{��_������Ќ-Z������ �gI\�<�{~��Zr\è�9�}#���� ���cMlз�v���D	���/�'�=�r���r�r��y׹@�ǫ�E��K/�,�^����~�i5z|�r_r|FDI���	��b�ye\$@����7z�j@��,��%6l�������&�^zY���=uj���\+�r�h�[� ����Koo7ea���
5�� �(�+��@������6<}����ݱfx >Q�xg�e����ZJ�!�5m�lX��鎞<��_-E�G\���^}5�7>��lڲ]<N5r}lؒ�ʨ��<*�^o{D�1.��!q��z.N�{����3d�zY+W����f��R���y`������9(�9��둯���r�k宻�%q��)�ҥK���Y��N9������
y��<������Y@�������$S�?� ^/�p���!	��exBdނ��)G$�DH�Z�EӼ�@�s�e̾���u�8+�-g�6wDМ��(A!Z��%�\¶��z��`�d��;Ը�+��!٢�P@�&�l�����e�Vss���d˒�y������Kz��j,?k�*K�.'@!l�Ndl�r�0�m��a<~�fwo��3�����vz�0 �����lY��a�(�/�(?��${5���U���y@=pT,�C�z�
jN��gr� �@��OA-��ۡk�:��!�U���ɓ���{�G�����z#�F>�C��葃l����)M��;Ŝtu��k[_�|�jȅX��~�E�J1[����@�yu��S�Q�t�!3�,d
c<:�B���4�P�Mǥ��$�f���C���������ך��t�y	���뮕��ny��	��Y���+㼏
�W��!�3�s�����5�6ˌ�3�+��5k�ғnh�/�q�_�N�_DM�|а��\��V�^#+� �;���r�W˲e������Ш���)�;!�
�u¶�i���^k �If%py�����oH=�t�"zsc�e��d`pD[ڍ 
��|^����7��(?���Pl�ʥ�݂5~�U�
 �`�������F�^��[n��\�zТ��2¸ �S��#�����Az�N���6Y�F���&���������p<��烬*�u� $ԝ777Rm�����Ϟ=[�=N@O*ȡ*���,O�s��R��z��g����`U���"�덜�~�н��i�]^�}$DR܎ �Dqzz���-������ȡ7c��3����(�<��AĀ*�j��hH��� ��<I�q?4|L��O�aw�����M�9�f�@�U-5u�j��r������d��޳K��	�;q��(�����g�c����6O�E/Y-�f/U��/u�Z5`��N䤘���X�x����{�!�Ta�W�y@���=���D��X�98�7K���
�  &�(�NƢR_�hHm�ID�g޳g�;v�ʩ��ҳ��G>"۶�&7�t�z�U��|�]6�d=0B�۽¡�eJ���w���j�p�ۧ���M;_��c[���ӹ��V���H�0%U��� cB�t\�پ�52�� ��� ���V����e����u���@G8J�z<�tfy�8-T������{��ʤ4�X�"(G�V�h7�6�VY�������P�MT�g=o۶M�C-�� �Rt�21�EGS�s�x�a2���6��#V��<��R�ϴ�t�D����g �@Dbp0�G���ř� "��F%d�c�!0��5�����*9u��p��n����{#��Dȝ'O��x>��ϧ��1�L���X�`M`0���6��	�R��=q�ǃ0��Cn�ʗ���M:H��)Su{YV�w#���;R'=]Q�U��¥%������֭a�{Z���6i�eK���W)�OH*�(�U�y@��s��%��v>���|6������f���n���V`�p�2I�����?r����L�a��
��ؐ�����!�@յ5$��졳�ʪ{vXyxlش!�2:<"����#�����@��3�Ĥ��C�(��2���r���O�[�[���<��3��y�ׅ������hH�s������f�&@���R ���nK��aI�@��~��d�*��sV�T����t�];��~�����,��	�ܵwL�� 0�ڤ80�O(h�Ο˰=���t��!7[��a����Dk��|��s�N��j8%3,|��!���BT���IN�:y�R^�r z~_�G�Nf�(硐M��
���b��ã���X�h;�̙�Ƞ�O��C�+"aj�]��A4"��ү���T�RF�FA���)�rJ�2��xX�+.�L���\�/�G��AP�(Uᠩ��Bς����	�#�����{<��ǔ�-�ؤ��9�C$�H��FE.���O���>*�^�2���d@��a���2U7g���m�S(\��(C�K��<[Xb�̦?(C���M/"/�O�R�8Aю4������;���qXlx�\w�x�hՊ�(�>�Nm��i���T� |YEک����+ܻ�b����}��Kk�}J��m���������a��<��5��<٩�i�����!�����2/��!\*�ɘ8��15b��5�L.����`B�T"��y��l��F�լ@��a&��Q��!�����îvmSejk3�$�3�j���YMm��G���8�RQ���3Ϙ��
lj5)6�z�`1/��(����1]�<zm��� -m�h���L���Ei ؚ�o��ed�d�.��ƶ�,�����޻h,f��腡�� ��hi����t��?3c>@$E��֭[Ձ��Kj�@`�}�\����5F�j$�5���L��~o�:M"��w�A�\�Q�E��z|FƆiP:Q�Q�q�G奪��=�ɑ�����@7J�1kJΰiN$RM��ߡ�6k���A�2��(��x�]� ϊ��8��R]f;O�dP��(����H���
��d &�����d�9>�;=��N��{���ﯪ�
���ή��K&�!��ss���jڇ�ۏ�;�t�z��<g+�!�˲:�&�Ȁ�!KLz��E���/}�K1��  �!IDAT���׿&0�h�2��a�za`��~��,h��R:����z��"���� �O?��\�a=�� ن�&�{jp�Pps�M����qY�j��}睲q�S�[�Dv:�t�~`G11Q��?X����w��l<7�tSvXt�h��#5��kT�[#F㤲�E��!��󗉋8��%"B�`-}0@�$�"ԙ��N��a�5��lP�Y�x	�h���_���6��ܒv˖M����Y�uu��������sF�/�@H�&	E���'��H>C��W�xtlH%����o�o*�2�� ze��1��Su��������acSD������,<����I0`�b2\��3��pVt�E���������R[WCO�NV]x�\}��r�]wJ_o��¥T΍�r2摗��;�ƹ��Ep ��L�"������K�&��.Zg��I���^��R��fP�s�I.��D	}a������m`��=��rި��@H�Bt�VI�PM(��,h&�#��01R���@$@#�����Ѝ(J� o{��a��k�Ex��`)�D��9|��_0O��yG�5@����F_��������֖&�!q0Αc�5c�-M͍��C����kd���V���u�~
�45�赂4���oji�0����9Ͱ�X녇��-����ݱ��X[��i��ǀ�?�q�:��=t|�0��#1�}����ܧ�ᕗ�R�� �'��qih�ȩ�#�6s����^5����
iiE}���d|Xv��.yɨ���W�����ʨ��4*�^o{L��N��\i�IN��{y����>MF�GY�@���ӭoh����G}��9f��A��Ƿb�r���?)?��e���r����� ����!a��cz��?vX
q�����u�־	0G��۾������~��5���VS�	0�%� ���r7���&�KMD=�(����aF'`$`�_9�à����(A �{}C�����܇n^_��Wy}��'i�wۍB ^6�ap[5�s��n���ƽ����g�k����@�W�FJYg�XR�N�>�����{﹋�������r�dxxHZ�"Yvҩ�ն5+�6m�\ W��0��LLf��뮓�~�+z�P�[�`�x���������Q
,�eb��d��ݖ�7����9'&S7��eD(���z37��р�B[��cɼ�R�H��:�2Lm����~��ҵ�J��p��{�̘�B�/�!SZj�}�f9߾]d��[����S&ғ�ze��Q��x�Ý���b%6@ 
��(j��۔)meB� �����;��9˟����ӳ����?J���3嫷�ƺg�q
/kn[�[���oſm☝K�f�ɔ���G�����z��\42��W {�PԪ�/�=��F��e�����S9�u�M7������7�=KІ�x��Ο�K/l�)�-�O}R6l�� ����xP��Teۻ��O�x�{^����k�M A��$�����j1��`y@*��nw��U�0��)��w,΂��K%3̯S2�(�M[ؑ��mx-^���n5>� �y}2]=S\��ǇM#�зo�*�#� �1?�SG����dhdT�M>p㇥E�,x�����$֯_��eΗ3�O�0u�:��˺u��~ "��s�I_� ����y	�H�`�h�R��$�!�)mS���~70�<;u�a,�A(�9��0���$OHC(,;v�k�y���x�O�_�J��#E���{O�=w�F�g���0�|����W�y@���=�Z&�j�O�823�|0ڡr�L�z�iz��fB^�p��������۾cG���7	ooP�������� �ʶ��cCE���<O�p!�j{�����xF�������>�[7�I���b�� Fv�M�u)>hD�GX�/��NKK��C����HQ���A5b��w\s�<��C4CF��-�KK�U~��_���2k�,���W� �Y�t[�� s�f�s�vT��1R���;{��vZ�{˱4�L!���O~�����3����a	�)ȓN����#�u�$����}����Ƨ�U�z?��z���q���d���g?����5���7������_v٥l|SWW�����R���1ft�w���/�� �m{e;#h��:���u6W ���뮻�x��l�o�y2�@>D����q�w�jL�}Z05c�q��C��W_&3�̤���7��'�]����}R����F�5F��4�ފ�^�uT �2��hj�1��⋶t�>q�����&%7s� B����O08~�$��h#�)�5n¹CnSn��_��@/t>�e>��yݔ�D^�ͦ/�r(��?ȱ�Qr�Ժ��ˇw�4 =V="	ӦM��� Wr����轝�G^���Y{����>ٷ�i�
�k�G�Ǣ���[61 �Gi������Db�^%�b4��A�~yf�$,�+B�&�P*G"�:�H����z�J�$���6�y�T.�h�����4�f��)Z��:�9|���Q��a�ȇ�/�c#d�����?}�������NM���J����n���[���������m�5��:�!j���x�B�.����_��e�X4��{B��ITB��A�^=Ͼ={�]�'N������[ϲ�����7��!.X5��:�C�hu�3��ў�Cg�TZ�EOP
��<����~?6��-��]"�Ɍ^�J�j�20�����x�Q�mT �2�e�͝ohj,��Ƈfx��\���86C��p ��*Pf^���5=��jlݼ�̂
z
����+5��r�9^1mZ��Ur���6�5��A�Mw��/�,��>�Զʜ��e2��]=*�׀��d�^�?�A���b.:�>f��y���>q<�q����_(d�S�A8�����[ ���k�ԱV)�4�D/;�,
l�;0�"3Ɛ(�Uӕ��[A��A�������|r�[����^`h���g��SO�SFI\R���tN�U`N�w]�5�WABG�Μ!�_�^^����t������@�\s������
l[��9	oޜY2>2��p<w@(�5c����u{�5�����e��	骼!J��P��Z�*]{���Z�2�m)��:�0m#ѼV� �3{�L�!���_����R]g�ytM�6��J���p��/T�?�pȕ���ȿV�y@��s���ǎ��j����3wY���D7ׂÄ��_�ݼt�N��V��C��H�=��L=OB�Nʪ�L�����cQ�rC��_X���d�sރV4� w�q`T�����x<����*����z�N�!�P�V�h����(G&3�W�pmM�:���䥻ׄ֡�V�Po��\2c�,�S���n=�g ٩^h�Y�]{n6�H�:o�u��@oe���'n�ߝr6⮟!|�ܰ�a��<E�N������h�R����X7�L$��N������Ω��I�5�C&�Q�:�E<nlNR ��.���͞-;��`�,=}�S0� �%(�=�=��`���f{W�L���/^�0����{˥ihۇ�+�L������������5zKF⯆!��)�a������1}w�$�%,��3M$�����hL��Z]c��y����b��_�T���F�+�m���td۶m�qD�%�O7F�<�2Y�H���G�Mݴm�Q���&�;]K�)a��R�I����`%1:� C[� p�9hĂ�-)�F	b�)ꪱ��	6z�5��m�U��q�x���V���ʰ8���Woq���2�}��68��lx۰p��Ǳ�'��jI�^7���@�u�/�Q7�F�5���gXK�}K}�=�{�r�ˬ�w�=y���ӰA��#�ys�C
�_�P � @�ܒH�:�~Q?�¯��@_��2�l�j�����Q?���ǭ�cBBUKM-j��j�/\-����7�������@���~�I�
���u�XWKAT�1�B<X����,��a��|���e��s6�s�2�0��V~�l�t��W׳��*\�w�.�&4�����u�z_^��UҦ��ht���*���8����G:�q�����6��D��ɿ�V����dr�E+t
F	�O7Wt��3����`������ջ����4>G�4:2,5�uE����w�o:�1c��m��[�n��pHl��d8)��wA�Pr����7�X2h۩��%:�g	E�0|��#�>{�\�����+M�8вn;W��AJ®7�`M����e�Q�<W,��=/{�vn㬗.�(CN���Q,���/@k���z�u�
��C�?�t�s�m�T�[��^�=ֈ��l_�¿����X2+��L��nYtՕRLg�ﺚZr|#i0��V�Cy��)�#^���+����X5���|���I���
�`:Zb@o%�� k#��(�ߡ��2�0s�%�Ǩ�(jpT;$���ѱ��_��+�����1]�[��R�q�G�+�m�X,Wz�Lr�*^6� 찑�i��AY�4<;l�`�c�X	�g�w�I	����tJR�\��>�P���'J�|��0kk�8o7�XI�31�uFq��i�00�Zt<���	r�ɉI�M}�OA��B����7��3]��j�Z��1��B�zA�%:���S���B=��U�u?_=Ť�7F�k��u6MR�QF��Wj�a�7���9W�߶��������ڠN�v8���dK�Z��2�^�z�%��7�ְ��TZ=�0?Og3� q���ed�N�L�s��H�C?��E:k�%��?���/!S�ġ#��8�����B
�z�dR�_�N�z�u4�z��0t�D"/�w�|ɤ�A�nIn�D���fv�>���N0_��^B���a-Dk� 쟷�{�����"t��J���Z��������dE����3n	��R��������>c�VFe��Q��xۣ��:��L&s�"=S�}��5jγ�"�N��l`�{�F6@5�TdC�YQ�E
^Yx���[7�n�Ep�C�#˰��6�8͞�w���K�l��7邩A�(B���\$�p���%�H0R#����
ֱ�|s�����)��<D�����Ƌ�W-��߾ �I����8tN�xKG�|�3���'T�����9�h�«����DG��Uo{�(�@�ո�1�l.k���F��3��e�%��.B%Y���Ψ����X{6_,����j �P<k���>���ԖV���e/z<_c0�P��U���*�)���Ճ�j����T/|
5���R[]/�h\�F�28�w��߭b�����q��dB�eR����H��h�,�炪��4u��]�����a��A���9�"�Z�P)np�_��kR�"( x6W✲E�?���]����z#�����Dl�Qg�!��[|ά�L��5J"L;�u�����{��6I��k��k�O����� �)Y���8O���G[[�dG��O<��Z���F���i�ܠ��U +��Vl��b��S6� H����G�t�k��d2��wU�PK�s#r���&\���^:� �s�����Zt��<KC��M80
nU�5�v��Qz� ���!i���9�f��'��Mv��@X6UG�=�>yc������g�q��)����
����ڵK-\luO�X	�F ����Y��y�7mZ�`�T-@�0B�l��5DB�	?�}c��"4�}����v�+J�0g��'�����i���Q j��S��ĩ��`kkkd������XL:::�����;|�0C�RC# ��ʰ�]G[�E>+�*DW���x�)"
~ |��y}�*�O��涙R
�q=/쥗n�U�Vr.C��2�Ɋ���|q�����}��:�&��K�1-�f��F���������D�(��j���X:E���^�yF߯ںF-j \uŕ��X'�?�(#4����)j|U\�z�"��p�4����z��"a}��"/���?�]�m���`(y\��Jze��Q��8��[�pa�#�<���cn��Q�3����07�z ��v�0�F.�Gт�������7� �-1y�|�R~��+[^�f�JdX�\n�bm�vh�&��$/���aD4˴�3����v�':O��L�˶�[���ȡ��G�u��[&�,�T�@��oY ��w�sց��y����{r"�9��-������p����=d�תQ��?>/�����eyz�?�0=l����׌�n��~����-�?�-]����=��#������_n��6����o ��>�1~�{��.%X����(��~]~������/���!��ԧ�������Y�9��/��"���!�����X��`�*�*��{��n��ɟ��g$�-S䦛>*a[)g������������t�p��j^��%By���^qS���p��r�����~9|�0���>#<�J��5�&5��zlZ�G&��G�:���F����v�P_�����}�V;�;��{�{�$�,A�w��:���p�|��|���b)'�aٰ�Jik�h4+]]�R�V����T#��Oڦwȯ����a���œ��*�oe��Qy�*�\�3�H���eX^��!]�t�!��ysd�u�����x�����D�=���W�X��M2�� ڛ�.du���"�|Z7z�=�2?NF7�ܳٿ�n�M�w�����	v�G���=r��X�����{��r��7ʶ�q�>���=X�CGʝ��-�#�'7>� @j����w��a��}r�t�<��sl�ZRGq^t�$S@@:_�fs��7.tIK�s4ka��AI�e^o�OU9D`x<���<�a�����.���{��1Q㋿ñY?�������΀� �^. ����7�7�Z�zڱ�;�����hl2�B�h�jV��k6g�F``�(��8�Ii׾�.Fl��)ٍF-�	�1m�z�9��b/�6ly�q�ԣ�;26*�%,.+��eE���fٯ���ۤ,�(���3Hm47��154%f��0�\��\q�e|nXCD_6>��=zX����W])���o��Mʔym��� GO��r\�z�S�Ζ�sfJ]}�d�	z���\ �Ϝ�9��ޔ�i(ɬԡW�y@���=t��n޴un|2�vXm*�Oko��s稧x�����*FEΡ�d�Pl��������x,*O<�Q���K,>�R��|����5<��;)fR 2��j���1ӯuZ�<��Tp��RC�Z�F�YW�t	�{�A)HA{�	��
����K 4��_8O�,[���V�cE�u��ռ�k@� �H���NɆ���UoP�e��I��$�$��е)�� �L�wmPE���/��;����G�����������w��g�F�w����������P���{�5��uu|4���V�V����g�[� ���غ�e��/Z��!�.iD`��~6mٹk�d�����
T�C%��������~�I����+�g���xB7���g:	��,���и����G}$F�i������,�c��>���D��2�9r4��w*���R�U�.l6=�KLrN�]w�\p�
������l�b��f�?SD�w�V0/�E�6�eW�����S�����ٔ�����%����I��2*�F�+�m�l'N�t���p��f�t���
��?�Q���wѻ��7B��I��?�����{L3�����q���b�Jy�ŗt�N��9SfϚK��i����Z���.�j��Ҕ%H��f��O��{�>���+e���
�9�Q72_�^�|6�x���r6l�B�8@��z��\{����?����r)S�b?���hu˙��׹�"�r9���?/����<v@�["7��������� �4�)חKv� N��0��� rl*Rc�����px�v<B���h��n��v�^0���(�u�Ñ*�6"�g�`����}��ځ(�ɓ�jmd�����癜���j6a��p�Ե4��������LN��"�4h���^%��� ��;��g�bVoi�|w@Dd���T��7٥��·`�B���M/q����y�K���!��D-^)��f��XTF�b����Ғ�LK0�c��w���0C������؍KeT�y@���=Z[[s�-�z���-M^?ac_8��:qLڦ����L�ou��_��1<ޕ�.��w��Gum��G���vʻ��7��u�� >�����~o�9n��O#Њ�-˯��~/�j��T��w�)?�(A*�V�Z�*zy�O�MK��#�^��jÉ�V�f�4?���H��v�<OH.mr� A�Ćk�y��T)p��Y�r%�g�+&G��y�ү�^X�o��q� 5�F�A���C�H��y�Zem6p��s��ݑ�6@˃����|���g�?̃9rH�	���+�n{�;��r���gh�?����?�I���x<Hv]���=H�<��w��P�J=��x)]�H�Z=�,k�!�LH[�t����HMJ��`��;z 8��hH	�/�c��A~�B�z��kO���g'݂z���Ө�Y�o4|���AQpBP90:��B� �6�[0��iB���ys�3���d"I��O��R���%�3��󝆱��xG�����8���q.��p��~�ח/�^�n�`�c�۾��%O(�����%���OA,˰�nh x�;v�e�W��W\Cp���g$�l~�(��]��jwP��6��ޤ�3K�!��K�)����̙8�	Wɐ%����N�OfҬ��B�8�D,�\lM8"��w��VOMI�Vm��2frU�������b~��組drPԳ �t�������Y4C�s��9�K�ێ����{��ӫΛ�=X�8$T�f`���|��q>����t����w�����o|������\}��4>����(�z뭼����^�W�9�{B9߲eKe떗�6'9-o�|��S��bw�n?A���C�)S0]ѐ�/du�]
�x�rE��^���a}c�z}�ԇ��%�<�ɤY��֓j� z��0���ߝa緋/����ӝ�I�e����]��`��y����)k֮V��t�z�}^�`�����'#�Q�yT �2�e��U��z��x|��46dx4���K����̔�e�e`����k�`d_�N�}��/��Ɠ��w��1
��wv[�|΄I)|��vMu���ظE� ��!_z�|�+���{C��[n�K֯�O}�S�;��q�r��>ʰ�Wn�����H��l�E�6j��
���q���H�x8dT�p���H�^�_�����>���7����b�9�`+���$)�}�o��mذ�-@���I��,C淟�G� x�����=2��=� mם��`�q0�x����	p���?�a�P�4��ڧ��@���׫[_���w�����[G:���hiJ=F<��T'O>�y�Ǥ�O��fr��/�嫗��[%?��L�7K>t�$��뱏+H��s��y�d���� ��g̜ɵ>y��:rX��KMk����73�s��qy����(b�gS�b���ܲe+]�i<�R�P+.^G���ǎq=��8'��H�$R}�[)p��&�,� >z=�ʛ{���+!mZ*�2�� ze�큐�O>�-9�% H�X2����.�|R�@7�h4.C#'eՅk	v㓮�3d�.cI��r���ɷ��=��o���e�{d��r�UW��Ȱl|�19tp?�Q���R���z�^5�̃'�uk�����A��+VPS��w�K��أ,k�>�eRS#/1�Wx�k׮%0UG"jd���g��7�浩
��E��!�c�e�<4�|�۷��4�C���Q~�� g竩�����z���#�s됐��̰9�����_�E��ܹs�@ �,�cl� �ED^x�j<��@�%��]h�)����	�A�?���;�x!�Dn��~��r���a�%�mX�|�t�:&c�잆����d��E4�}ة`������_��+��T}f��|��o��/�R:�������?"����\y����}�ލ��c������N�w���+��52ej��{�]$��]��>��쥗^ʴ
R��#�� ���{��#ᵫBq�O@)��]��v�RC!%S;�$��r�HN�8�sm�r^��^�}T �2�u�NW	^�GA,��Wt��U���a��.M�w;�c��u�F����L�U���w����uy��G$:6.�m�
H,>n���<&L��o�Ac� Bκ���)�b� lb���#�������~��,:�A�ddxX���os��wN����y�/����K����,v�;7���U����{���,%X!ߺc�+��w��f��4��V� p@6��,��X'��W#z?lA� ���]��/�`H�������@x�8�9������Gdyp����.m��n c�l���*Ќe�����.�L�'��a��3�<˹X���"P�����'%�T`��������_��Ng����뮗��u���i�>x�5�����ȣ?"�\��!u�ȇ�/��|����;���7J��w|�A�:uJ�c�<���x?�Fx�=�(����73ʀ\�����ګ��a5D�L��"_�kw��A��`��y��]I��ZԸ��T4��zQ^۾W�	5j"2�H�2*�<�
�W�9�;X���Ka�yII��{	I���Ț�6�Kͨ�54D���� �6qR���M��{%�W��/~�����?�/�:�&��ς�~��[�%l��V3<�O����&�����oHl<�\�S'���,�?�r� �D,�F�G7n��TE�<q�j�,Y�D}B=�	(q�(D� �9"/�d�B�E�x�Ϛ>MZ�UArphPB���.���A�kb�r
��;���߰�y&�*�nx	<`_�^���F���[⚸K��R��{��k�/��r�@�I��1;o��~Д��wX{Դ��G�׵���S��W&��hÿa��cG�\��PȩϿZ���;���d��t&bI��V��.��xB��n�>�+�֬��3g�z\�.}���ky����� �{��d��r��A}W��Ç幧�f�;��u�� 0T�n`����~��7oz��	�F����M��%Ԟ��ǥM��d�		E<r����n�8�^�?�3 ��Sv�ث�_�^���R�q�G�+㜆n���pU)WȲ,�`ש^�B�ٵ{��������߬^�@x� I��M' ��ƍO�c�="�Ǐ2g�m�Ay橍,7C���3)vZ9W� ���=�V@��b# !䋰0���<�Q����A�ē�6�y�U"��9�y�7<6�{D������=���d^�#5$����g%><����H�㓆p��wz�t�˔�����6��!w��+0l��#�`�§M�N�5���z�y���Y<c(��댬_����.]o/$QsF�=]ៈ`�-X���nGxv>��9A�aD���Gc����U����@��5��O��
z��t����c��Le~=�H�G
K���}j@������>�9�Ŀ���Ȼ�q�$&bR�}�kx�D\�CE5���U�*}��ɠ�>��{�K*���}j�>uBЇ�����(�(��
���j �������Ts�!�N�*)|�0ŉ��e�+�_�&�V���QN�R��N��8#��t�ڋ�ʡ����/!�Q�yT �2�i8���nҥH����pʒ�Nw�&y�+�d��X�mk�c�Ǩ�
3���P��+����a|rB~����p\Aʴa�S5�ނE�@B�_7i=��Z�~��Ϝ9-���*���
�����z��˛����ydlx��XlC�k��F�=�y�D+̡��O=K5`-�z#�#�^�hm
o#�^�m��Ǟ��ߔy��5�m�܎8`�)\�n�s!�a�PALs�9O���d����� + 1�7ae�f��� p� ��ڹc�Ug_*���1`4���Юk�<Z�Y�.k�r���)H.o���=����u/^(�N�f	���(������!��׾ʨG@�sh�>z���:��-_�t!'�g� ?���K6��}���{d��9����r��!^���#�/�������S���6J�m�`��=sv���D2ٔU�P���zQȱ�Ȏ'�.5B����cR�����.I�2��%��]��r��K2��ѢTFe��Q��8��(8
U�@��5X��1B���X�R?s����ꭍ���db�3Sl7A}8J�N+���FP�P�'@����^��EP�2�|_��רQ>��Wn�� �I&dHAr��e����Z�������"����Bi#�OŲ@HN��y@`$�W��Q�Zc�\R�\/�PS�^5�ﺰ�ڿG��#T�{�٧M#�Y"��Ҩ��끐��v���nwO������~9����� ���)΃|;����]�Ʀ&��Ǝr����>�bx���o����7��^����:�#�u"hI���	��y���c���Le���)D4��Aܮ"��@h@��ӧ�ʮ]��r)f&����!/>���S	��w�Apt�����d�O�p�)�鏾C��J�?��K�բC��e��I��3�}��!a��h@��H�s������D(�y��F�t�Q��8.oI�./U�R���<6$�J#|�!py�?0�-��OIu]�d����8���qN���no��6�nʦ��9+$nJ�|^S�+�u#�r����!;�͖����	�ֶ�S/�.���M&&��ߡ�K��z��x�4-Zw�W��;�2{�<� �\� ?��_�m����=&������fMѐ�X��mjn6�b
Dcј\���z��;5�Yu�&u��Q���D
����i�n�`{C��u�ֱq
��dє���:s;m`�����Ϲ��������M�X���Ɵ�������
T q��e��x2�,��- kww��T�ӵ�9G��X���q^�Q�'85�hЃTD\����4JvY}��H����b4�2�s�Ёߴ�Eٽk'��{�G�(�Z������3�?CO:�NP2;{w�.�_���;g= ��/�G�����	Av7�����:u��]so�أjat|��@S�H��k�XM�y��#AGX<��#���k#|�q��������	�q5bgϝ-C�c���2����T�qN����
�*����
óF8�^ Ox�B�aq��&P�Vw��
���}A���1l�̱;��e�ӂ����T�\�����Y���=���mV�wu�f�0��0�=^����IP �����MM<�k�3�A� 	Y�ދϫ����pL��ihi�l:���^�ð��$O*�{�^�~�"u�SP�g7>�����~Mz�tXح�h,ǑCG�F)�uURWS��ٺe��1�N�:eB��W+����:u .8 �����a���!�ŁB�]O߀�VA�����Aą����
���!�:�ƁC�:�(�;�n.5�z����`
����pt�hc�_AzP����KC�a��y�}F� `
T��q���(�>�����\S��c�F�z��iG�5��ޏֲV�^tҼ�2<h�F)#�}�x�;��Q�3a�A6����[ �Wr@���C#��n�D�h���g���u�VY~�J�#�S�q�G�+�<䯍��!��0���]^�	�'
IO��T�r:��TK�fyt��wˢ&�`�N�"�mT٠cr��Po�vR7^ 8r�v�4����y�u�v9��.uKe��Ùv=2A2o:G�N+��䩓���1C>x㇌�i�l��\��b�}�ꝁܕ��x\~���ȸ�3��U��T¨�Y�l �݌�n�b{�8[�T�f����		����S�8�����$1��Q�ෛ���������L2MC������ϱS�[��L��&����7]<t-3y�-���j��q@�[�"?�pX�I<�b��-_����~HF�Ǩ��~x�h�:(�ć�M
�v��f
��#��}��w�V���0l�����=h�bB�����GD<��u�>FSH�y��)���cH�(�C�����e:����;���낮�n4*�(I� ��M����*9��8��qNá;g&�*a/E	{�뮏�+ ���P'm뀧Ha7K�!�nt^�F�4��,��S�9�Gۻ�$Py�!bMNNЋB]06^�b��O�DF=��H �
�u�uR���ʇG���u�6��ୣS6yD֬Y�?�y/��靎���7�<��߽s�n�.��}B#�aC�O�V^#��^ѽLs�?úb^�,k�̡T����b���u���ڧ�~�v��`����1���#ɉ8l]7K	��'��U�@μ1DUt��N7+ `��~�(�̜%�(Ӱ.0&�Dr�LΩk����o�1�<u�i��Y=�'�2S����V���_HldL���;�)�hl����%�d�S_����9vڅ�%�"fg�)پ�5��z/(,��\<������a��%+@
u�#xo't��<\�2��H8(Y50����@�٪���Dc#$��pҌӤ��Z&��aoU%�^�}T �2�i�|��n�dj��^��%��ƘZ��� #4� �9�*�ON�x<̑;�� �b�4B-KT�(fV��F��v��y^�7��o����!S�?#�/��BZ�zmPT�wjÐ5�3�xy��z�����%�F����=�
���K�a ��>���%����Az�H #�Ȇ4а�!%�<+<:��]e��mL 쑓�����z������7����*Lcׇc�@C^��a�l�ܘ;�Ɏ�&Y0�蟞R���� ):��v}��.�<��� � ��.p���x|&��R4��o����/�ۿ�npjd�Ͻ�wѓF{Q�s��:%����R��R��F+Hà<np�_��\q�r�5W�e���X��A�|ꩧ�5�t�t���<�?G�[p.�" _^8	��|�d�z}/ۼ"
6Sc�$'�RCI=������U�b�2�>p�W�mWcb�<te����,_vA��2��� ze���M��K)� ��-芻��\��d9K<%��0̉&Qv�2���6��P6T+�^e�c����µ���cV���<�3�� ��R���w^r27n`��t���И<���z�4��ཛ�9A��x�)SZ��7HmuD�͛��k�@A��;vJ_��ׯ��B5�)I�n2I�V4h�����<��C�����5�w�e�\���v�O��\!���#a���Yo�H0�q�|�;ɂ���?,##C$��E��V��P{~��W �n�*�<��Qq:���p.'���Y��ϮI�P��t	�"��n4�ry}+Jzl@:,�j�L�"ߺ���^�������i��{t�y�M<�enJ���(��)���g��CZ�J=�^B 9O���A��xh��|�5�]E���2sTo)��>��)2g�,Y}�
�={&���^�B���?��N5t��	����Z���Z�1s����%�:�]�_�NG�����t�K<���S��JJeT�y@��s��;��1��
��Α��l$N�a̪p5���=N �&�P`+2�ij��7���8eH��H�� 	����S�Г7���>�����l�lPώ�;F6c� 9@%n�q����v;o��z�*��x\�z[�������z�	���Ua���R��x�(���QFV���(=�6P+�Ovr��
t�\����Y�x����[���׍�@��dg��_�9�R���+6�	O�%o����]G���'���X޵�g�i�8��sZ��wpxHR���!=���˴3��5�ՀH��:9��بz��I$��e
Egҹ	i4l��FI��(�z,;�Y�yA��Z���9�Wa��9ϒ�+�G�cr�ĉ��=�p��D`�y��>��>v�sy���Z>��O�qYE�fb2��b�!",�� [(ɂ�sdZ[+K,s9}GC~iW�*61�?q�7w��~������|��W�{z��2*�<�
�W�9IW6�t�����Ml��Y�{Fg��s�)�6��9�َG�}�v���<�65��u��r���\��}��YR�P/�bU0��i�	o���$�
�)�}�\uܬ=�qMim�טͨ�����!e��O/.�𱛜0��zp�_�PAtǹ�PF5�}R��/��^$�-2���ǏQ#F<;�."({`��z"�*{ո;]`x.˻4=�kk���GdӦM�� ��b1��9n��F�^9}��Qf�5�2����`��c,&�>��!���
���Z3�]��ᱳ{X����!֖������a�Ľ��@���t����"C��{T����������=�,ǆ>P��g �`�n���K�y�yH�xg��������}��3��:�IFIJ�3  7�6/u�N�4�k�e��7������tK(�����,����~5��̚�������e���a}W�f���E���q���Rэ�G���D���9*�^�4��#\]Ŝ9�a�E�0��eXx�����W�^)N�S��W˚��h�H�"��ӟ���?�u��,7��nz�(�Bx���Aw�b�{� ��۵�بq.l���Px�ؐ�)�;������gJ��3`���vK��_���(�z��W���/c�}�F}��ԩW��|`�OH��`L�Ũ�=�B���k�j07��@�A�4 y�; �z����T�!���CKK3���s�4:��bq����J
�t5�z��G��24<�P��}��]TO��3�2b��Q0�HQ��a���5�:���,k��i (� �&[�R �K뻁���zy�R��T:cU:LH�J�%g�P6�gmK�ڑ4��c����ߓ�4S)N��T�;������u�XpJ"��-������#��)��l����9�tH��q��T__k�%�r�UWHuM��IFr�	���J��.l��S.��y�Oˑ�G�3�
�W��@��s��ǡ��^*���#�v�*je77����n4a��z,�p�G��;���-<6X���%�d�?����1c�n�Ez��O!ת��*��ɶ7j�\04"7���N0�ˎm>��|���!�"�@/�z��ЎՍ2-�>�o��-�}2w�
)�|�+C��F-K�����a���d<F���t�5h������$���6�3X�g[��-涇B)㡎x�lx�$l�r������u�I3!��[[�ȡ�G��� 2�h��g�NHUu��}�F���/��1���p�H#,_C��[�X�t�M�w��ߚ���:eϞ=�O*�f$��������uAR�n��e��|AFF�e񲥲h�Ry}�>�%�H�$����|�h�w0�p> ?J#C5U�Ԁ_�����AV���(��c�l�#��r&�7�#�]wݥ�Q��^}����ʈL�|�Vq��A�B]}�����i���&]�2m��3�E�9Cv̢ٞ�P�[q�R6��vJeT�y@��s U�'<B�E�[�p^~y��x}/	\��;d��7c���v������m�y��C��=o쓛o�Y��Yq��?�����I����9~�(+{��{�f�]^���6���nɒl�r�lp��n�MK�InnnH!@�IB�(	�H��ĕcw�"[��Q�hz=����w�����?�3����~���9gw~�k��%�;@��T�e��O҈��� C�< �R�QZQ��(���icE�T<�2�dϮ��w갸Q�X�Z>(s,�T2MvC�1��(��]Ft_���"��ֿ|[~������>K���&�W�1m��Q���F3� U)�1�k��^c�1ӌ�Nv��n����}g����0���"�0�˞V�?��  ±�y�ܹ�t����ٲ�*��_���/��;�����fd`pX�� q\���<��ȩc�lIus���EN��!Ȧ�cӡ�@��K�}�(f�;fϒ
f�]��LJ����H${ʵފŋ�����I���k8���p�y��/T�ӄ��[��3��w�&o���X/%u �����o�o��5&�ᄓY��d벥dD)e玽z=B�v���<cA�i�̞�)�y���p���y� ���%�Ѫ.�^�d��	]�P/�	f�W�X�1���!����Hg����P�p�<*���g	LX�1Z��楛�dp`�$1O<��<����ls�tg'b1FQ�F�,�H��tՀ����Op�Xt�Nh�|	�f.�Q�:���#�f#�'�o�
�.u���@fh[K�v̯�XR��j+j''���9���g"� hQ,������/�G���g��@.pQD��;ƺ������a���'>��)��q�=y�)���F��,���;���!�Pmd������w����;��F������}r��o���w��~`��׼�g�(G#�`\�F5J��E-���9�';v�欶�rIL�/�=D?J!x.�͛C��i�|`kCV�\�0�9�a������s�.��sX*$!�S�͍R����䝷�.�#Cr��t�>%+�.������R���'��,N*�$�0�!s�.�#y��af>��I�y��019!Cz��L�&b��λ�،L��Z.U=��]wJT���e�t��MH֡��-,��
��+h �C`��E`�h��'Oq�F�۳:g��3ݜs�xQNh �l,�b�P�c�R�ZE0�<���+�a~��5B"Mmr��q���#�pԤ��9�@c8F��ZJ�����j�d��Μ�%x 
D�5�����/���d�5�vq����-����=�|�r��w�#��k��NN�� K�jS�#x�ǽiTcFP>@������)�h�l�>�<R�h$�8 ��}GHނsQ0��MO��kkk�|�C����wHqrP��~��'6]|�l\���g���G�H��@y[��;fu�r��'�Ͳj���$���`��z�i��Iw�)}^\Υ�Z5�ש��3�R��Mfk�/<���WG �I���������z�<��G�'�ʭ.^�@��I��L�NW��d떫����òb�J�sDc)�& ��R�	(��څ��۵}���9��%�=1���ԂLՠ�y� ���E�9����뢚#���ji���QY�d�Oh�b
:�]]�LS]�yy��(����_}�e�Νr��k�N��V��o�^>�������������
E6�!U���Q-�ϧӣ�M���ӊ� �;����N�^�n�ē)C�}t+��0�d�"�N�Mi`��mDA �FUNd��yT{�p�juT�ə�dc0�����o�Q?_����OH^�)w���r�Iֽtx!��c�ǟ|��e-�-������~�C�y�,Y��Mz�;��x\�/��/���fy�Ձ9"��ڢޏc b��^~Q�>&	u(�u�Q��y�0DB
lW_%o��f)�)U�E�ɏ���ޓ�J'��+.�+��T��:"��qM�<����[n�����t8.ڴI>�7#��x�Q�;Z�|]z�&ߊ%K��_��|��T�;�۽�-��e
�;�T�!��nx������>c��mo��(�앧�~R���HҰM��OL#dF��Β��v�:|�NԜY�����%y_P"@�&�I3ˁ����4�������A�a�,	�_8�~�"5�ŉq��w =�Y(�b��Q�mLCZu��%\'5b蓪FX�7��Ex�4*�  �HfY�r>w9��,����+=���[�[e��9r��I���2�B*�)�֭#���?.���gYƼ��7�\�F��t2�D�1a�b�ۚ��o��Ψ�嗷�O�Sը�l�P>|X�{�oˢ9�����{HFsy�i�ɴ/uZRG�Zٰ�B=�a�;#�(0�E�B����G�f2�!��q�R�@�{8
h��KLuh���Q@����&��zdΜ���
޻������.�T��O?,��ֿȳ�>ˈ{Ӧ��7���O�3��W�{��=﹓]�]IƓ��ϗ舁;=�2t�}��l$��@u�ת��Ǡ��l�H��h6��^�QF�W^y���'���Шދ��eP�wǬv�ù@f���tZ�ڷo��3�k��2ݒ��t��3��}G\u,P�)��G̔����(`�WOc�"*M-�
�	鈵ˢ%�J2��}�ꬡ���B�_2������o{�:	o���1D���u�F��1���-Ȇ̟�rRkK�F���hLv����@���j��;� z`3�����z��XZ�D�����v���@zߩ{���Y�FF9��g�NΖcj\H!$��u�]t���\sYΞ~�iC��������i4s��7����x�a��?���LoZձl6_s�{���5�b꾜'hΟ��)nl�h A}�ca��F&iu|��{�M֮X��\Z�.\L5�R�0��p� h���Fd���0���HԑD2BSS��_0��k�g����`1�$J8ac�H��;jq��})��s�a���b!F̔��e��R�̙��}й��3�ŵ�l��T8����)t��#`\�b>G^}|�\D�C��ǏvɂE�%��܋�	Y�p�:M1�3:��}���:���������gg��ػ{�l�t�<����of����W�ftxX��G���˖������� �Ͼj�G�Ȣ\}�՜?_�z�̞޳h<KH�'���#q���"X��{�Iu�z�<�[��6���H���� ߩ۪˴��C8�0wN��W���H��>y���e��#z`��(�SF�$*�{`��@l�(�Ԛ�ܪ'�g�ʳ�|��2h�C��������m\ ����ܰQ,bc�ٞy�{����4^*˷��H�t���^6(�7=��<�HE�d��5�f��t�֍��y�$/��]�ek���j���)�jtC������/�$�/X+�M��F��w=k�/���/�U"=;2��l�,���G��+�x GM�#u��-���8���
.+)h���=F��3� ;�*�ؔ=:֑) "zň��`V+�lRko��hl2T��,S��&(�<�0t[c���c��P`^����N	u���AW<��\�� �1�1�>uZo��K��n�Ɋ��HGM$�Q�~ %�2��Č����/��N��?E ���^�:�#Qyeۋr��G�v���X/�dT���Y���vKS[+�o�م��F8_���S����C�ɔLf����3�P�����h�x���c,��*m{�En���`�����ohh��:��x�2�ݺ/��ٝmr��O~�l"�����g���@R��x�������+ ��Λ�،�r!�R�R�t]W��t�8���F�'uq��4�� ,��X����m W&����(]Gh�G|�T0���S�r�`TŐ�N�������o���R�������={X���Q,�ѮF�al�5�iO?��̞5W�{õ�~݅윏+p$��F8G^�	��g�S�dǞ}�J߰�"��O��]����ȏ�޳S),�#�>6�MH�����Y�x��UKK�d�\3�gv{��K�T���G�/4�f��u��w��9l̾�Y�4��HA�VG �Qu{kIt���ǥ0����80�U9
�Q?�_�T�nz�IY�'�idȈN�WxL�x�F�)uf&�`�PkBA3�ǎsU@�;{V��eѢ���ϫc�A�8 7�t���9:�w�D�Ȅ"�T�h���2�ɤ����qlom��:|���D����s �t,%���作'�����hw���Ks]�6ކY{��~dǳ
�f� ���A�D=��!���R2=�ْ>�!���J7���䋸�)��-��$�����3�<)�����X`��@lF����!�C��(G�V�hqb�",n����M�A��8�p��2�nbjML���-AI,j�سɇ	���U=_��B�rPu�icX�.�H�N(����r��A�m�V0h��@F�o��;�ˈ-�J�a�7[����G�~vpD����Y���b��͌�!*S��n�����	���)�����PA�����`�42H?�,��J�rd �����T2���Q�f*�\�r���(C�u_d���Ld&К�v1��������x�N≌O}k�=R���!����1Т�,����z�Ca���H��4'�9�4�+���/��o���w�/���D:��N/�ߢ��?����@^���?G>j�(W�,�雜dv�����E��욦8�;��%�#��
(�5)�q��1���f�h�ٔ�3=<�L�0�����J��ƱD������3��>��;."���v<��8�"�-TX��lsk;���2�>}+	,��d�6#S��WJ尥´�� ���X ���ъ�.�0�-=�ioD���f'�.�!�����oh��<F�%/8��@�	Mp�yc��\9�9<8D�EC����B\��Ƽ�^&f�*�J2RΫ��ՅuiS{�2�M* �wt��<���f��6�����'`oٲ�s��
���jt��#c8p4�Ɔ�-�SG5µ:�pF&'rr�W�]p���wP~��g-`0��s$�T��C��c��)�#�����g�=h���,��U���m��W�(wͺ�(��XT]�r�@�F��F�h�{ߝ�+/�,g�X��nb�]8rW��;{�Bɏ��|}P*���{ꩧ�ȱ��ַ�C��[`������]G��x����b(|��ᬠ[-�秊Y��,w�^�&��9р2�>@pH8g_(֚���+�k�i���}�x��O
<w+k��*x�"pL4���>���${��(�Ye��+K2����TM�d:�X��o�(�v�, ��fdCC��
�q�+�P[�LfX�h �I�`���"l(�!�I�vGC-���[q2��J���� ۙ�"����Ξ�ś����t��ڌ�щ�"��S��g"��R7*o���2�C�skG;���5b�(��ϥ�t����avm#���F�C���P��B4�f�J�#�Gz}���,)`� =��������/{õ�ʃ=$�3�^�n<i@���-x���y����=^��-X�Q�$�/��X}���)un
����)�'�7\'M����[���N��z��-$Zٻg�i���qL�ΐ'�S؄�>�N�m&�>3�:�����_�lꨞ7���ٍ��&=����%x�9�� u
Ǥ�.]��ԁ����ۿ�}t���^ukǃ��=l*̚�U�|G�R[ *��GĤ�j���ngt�5���:.��xNI�k<,����v��(�d��<��n�6#IV*n�\�0��t�0�ѴƨiPr��1�����uJ]���M1>|Lf'��I"�t�ˆf��c.ӹX4Ѱd8�#,ܖub�2�h<#;S��jHas�M#�R�8!HU��w��Ȱ�-W�g�Y���m/�Ky�ؿgwM4)al��l�ȃ>�q ��W ��k6g�K��/��'���y�3}��ժ�Y�z4��I{��2��"����a���K+,T+�b@].$�C&B�藠�0��qT�|��Br\J�b���7�ճ� �Q7:����2�S�-#C^]c��]���CC#r�=�2������0Rfo�kt{�0Y��9?�7���c����̀�T��D��e"�i䃳X�j��mæ-�ཋ/�X����L�O�R�9/_f�$ �B�sd�@h�T�!�q$��@�i{/Z�s��4p��I��7D����%��� �;� z`32]��p����d�B��� �KɊ�
ծ.�N��Ya_Y,�Q:@!�Q9��W�Z��cǎ0{��A�@�>�@ي��� Q4l� X{���l��`!��E�Z&��E��j�k�<<2���)z��F�Jc'9꼈��	5]���S'��g?{��ph�CP	B���~���|��G�n�� �����6>c"ư�@*�?��qޘ��3w6�p`PC��Z�[�&�n����v=N��"c_*Uǌ�پ�7���`��`�|V{��Fx̨���U��� I�7v�}��_�'ٽ{�̞3�]���P� '>�讟cm�p0p����@F�8�+��L�9B���˧�kg�f[�S����ŀ�����)X��)���A�)P�gY�l��L��w<a���P��FB�?��ې�&	��*�%�lh��uB���F�#_��FB!=N)`�y� ������"����>v֡���夢�$u���ʦǙ��u贂ʻ��n֣1W<11.+V������ޟ�޽{#F�\�m����<^r�&9}���BHD�8�Ijr��F�ji�*S��.�K�[A#ׁ�>ٸi�W��(v���|�{X��t b����u��O��]	J��3��������[�4� D� Iht�v�yp&p>P2kЈ
h(?��%��hif��sĈ��8��Q��9�s�(�R'L0��:L(`��k06�K���t�4���'?�)�#T����e��E|���ַhT=���{���*]4���D��O|���3OS�i���
��V�<�c�RIa"!F� KL- TAT�h `���=��1a��U����8w��H������F?[ú��F>��,?�q��*���/�k�
���e��&�xt��@��vuD\�~��I7$d��%�~�ξ��q��|�}��<Jj�T�EܭBAZ�=1s�v�, ��ffUÂi�h(�8�"M-���x&B4���Z�X�E7�9b���N�x�F]w��CFTH���> W]��ihHt�s�h��&�}``�@�(z*�77�5noF�јQ�#0�3R��6I���.��-;F�,5*��l�
��z��F��@���wH����ui���{@^x���C��n|��K���u���Lm�� kP�^vŕ��1�#���?�q*�}���y�+��/�h�8���+]]]r�eW0�],�(��	�����E6����@��ɧ���'N�m����/|�w��&L�669��W�D�z�GDv"��ǰg�F�8p��F�?F�j�|��g������|Ե8>�;�<ܲ^ע��1N �3<:h�>�
�I+�cAc$@d4�/t�{b������խ s��J|���]0k��q��Ȝ���ڌq�3��c����|���38IF�7���W^*��. QMZ��&S.�喛�s���<�Գ̮�A+�X���;O z`3�H<�4�5u�pu�z��Y��s��ֆ�ܵ�M_!��yaID#��~��y\���A9t�^�)_|q�\����k�5d��Ms��t�",Dҵ�d�s��E, �V��n,�`" @� R����/VB'���b��n�rG1�E�s��
h�bW�;���L����A�u<�`M���n[�|�H}c�d'r�\�I0@�h8�f�əguVp~ ���p��?�����-[��\iZ#���,�L"q���(�|�*��#Z��l�T:��o�f��]%�e��u���Ѩ:_zݲ�㤾����e�~W��PP��j	u��r�	6:���=8f�Sr��έ��K�ٔ��76�U,�~����	��104�����ѣG����@V�^%��M�����Q���^ɛ}�g�զ�A�J��\N�OJ��(�'>x�� hl|X��8%dA����$_��7�iA��"vʊ�K�h���.�,͍ͬ�GÞ,Y<[>������?�}�K8��E0�[ ��Ț��A�AqԸ=]��Q^�|�������PJ������}���~��jݩ�&lQ�C
��!�h�QbwL���Ozщ�1FW�H��Q j�gVC���8��ś�G�,(X7n���jH]b��8�T�Y�.��9�5�c�l8��!n"b��O%R��ҪQn�������؈%F��4�Utq���?L����o�\�ϛ�����p�c.\(����$��7�����%�6˩���ǲ�+�myWD�W_��b.��d_~�ev�#��3g�����Qx):\h�CC�Ui.��靀�y��|����q�Ӣ�k$����s�������1
o�ZF�dULD�s�1C��{�0��;v�`#�W\�y�\!/���+u�[�x-�3<ds0Rȉ���l�3J�9u�����2'(���Y�t)�W׉�����7^w���'?%�7n`drb���p :;gK&ݠ׭�P'3�)�\��g>��w��/ex��Q< ��j`��@lF���G"��F[��"-͍�b�
��+�P#"qȢ%K�����~��ӟ�������7t���۷k��jX)���aini��{�����Z��멄�hż��ƿEfЉ�� "��e�]&-�h�)����{X�;;��jGY�'���NNL�.�&),����s��~�UH�L,#xW#��$'l�'e��Q��x��$	D�}g%��0�1�q�~�6��8��\V�b�̞5� D�k֬a����i���v�7!��kb�JP�X�d�tΞM�ji됵n�,9�߆�F	��f ҆�=F�|�م��av�Á	�c��#�A�E3�`$X#��2�X�k��o�F�l\��{���Z�����H���stv��~v��C5<8hg��z�8A��~�Y��7^�^.X,s�dlb��hQ�=j6H�6��R�Ѩ�����:�[�v���=æ�y�g�Y:~��/�%h�oVǲN2�zO�;;$��#��>�A�K%}B��\�y��^�V�{�e}�J��a	,��h�6#�帊�ꢹ�!G���s�:�Zo[�,�5�i͸�_>[Tp�S*���G^y���.pFV/��`208L�K��$�	x��Gt���u�XPmDgǘ�Dgk�
g�_q�Ul;��+Ԯ | ,��f�/_*�W���k�ʡ��9�擺��Ă�Uy3%F����bDZ�Xƿ���nے� ��-m��1�~`D�VČ�g��� d\d�q�9�t�M�<�ϔ�^���z3�mJ�Z�o�F�n�J��h�x˛o"�;g�Qvn�#}��uj��^,�!���F�$/�DR�dC�/y8�d547q�+�����0��{
p���6*�cy0�+���8G�F � F7����L���絏����<�C��Oɺ5ȩ�]�6͎�`;6��Ʌ��:ijm��;wȏ������[�T��:*���o�����'x��r�lq!�a�-������R#����u2�s�,�?O�Ι�N�^_=���V�cO<�RR0��y� ���%҉�b1�WT#�ʙ�%���.M(�
)���)�<9|p��\IS"x��}���e��92�8ñ8�,��I*S-K�3jW�FG�����;��)xl���� �u]���9r��p :"�|���x�ʉ�,�94�%��it?,q
��pv�Ԙ��?�t��D'��Ҭ�.�E����:1����J�ᣣ�2��Iƣ
������a�H��8���GĈ�}P�r4���?\GP��z��C�)r?r�#���^��78%���}\+��q�t�[�9�밀O�D�N�瓸@�!�>;S�јߠFAF�ǻNr����(�Ȏ�+�s�O��6u�&}�N�͘��2R=�}��ҷo��R2'N�6Y�f\�\k�D� �=�+�?�{��!����&9����#�dr|�R�84 ��&u��&�������L7���P�(�DF�X��5��H*��?%��Σ�،��º�c�)�ʙ���q��KǏo�:iji��0���L��9g��Ѯ�
zI���7�����[~�ིo�.M؋��5�b�̶#�}��eժU\ı�#�j�1����L�U����h���]{���X�O��0��4 Q1�lk6���Ƚ)�9?en#N�\g�O�aCւ�����|@�Mt� ؔK��O*��s�.���q]+
 l+���[�qb�+W��[�+#w�v 0�u�i{��V�e0U �Җ�V�(ͼ<�gѩn���Q3������!S$e����IȚ��F�k-������q3?ڷs�8vԶ�Y�q���ܑ��M�}�������b���;b�����}}��fs�ф����P���O.��b����:O���̓Oȿ|��2:8$�	Å_��I�������#�Y��T���g�_o��ޯ�+��JH�v>- ��fd�C״� �&��E�� ���]:;:�(��94�/���e��)���?:��)����F���rՖ-� t��m��k���G�%IɄ?g�IQ�J\H�����ݡV!��qp*ȴ��@���ܳ[���J�mG'�b>d9�6vz����=�?�]���V�&�c@��;ߦ��;��F�9���Q0;/�� ]^e��d?�4:D-�b ;�Jc�FZX@V2�xz�rc&��:�""Ih�gsct�%iI#~�]�U ��q�r���c�ۙ��.�B���G�C�[�����x�-p)@×�fY�l�Ť�iiie�:���T��Ą:g���d��z\�a��yWMt��Z��q���Эٲ�uĬC�ϣ Uo��6l� ��=�vJG{�\�~��~��T�{�'�J]Z�����i�l{�9�xQi�5W��3��G�h֬&=�F�:v@Nw�D���!	"��Ϋ�،loqĬ����>i�kT����I�?o��s;e,�;�N�9�߼��|��o��_$����P��x�ER�Jj D~�_+�J�kin��E���`xޱH��cIy�2f?��3��*���T6�G��x�G�UC��.���>�N���lԎ�7#t��Y����������L�S)k���k�7:6̨]��=����T�E�H�'ň���Fi�49R��M�{��Hۤ�I،�^ !��k���3�NK�١~7�Gb����Z��#~$TeD�T�+�XF�:ȣ|���:<^864�Q�G�q�ᘠO��Fr=0�Q�M_p�U��8��x$���ɮ�^�����V*���L�>�{�P�5���7�s��/�����Ô䝫�W��%�|�e���?ȴ��c���L�َg�~B2��|�B}�]
݀6��{�g�����u{M�F�A�{`��@lF�'���LV�h���Wf�u����ua{A�����HF�ޓ�9u�[z{ �bɕ�ƸLd��,^�X.�K�E��wJ�H	��tS35�㺐C�
فx,E��2A�
pD�gN�HǬNu8b$q��H=������qv�[����Q����6	KE#ّ�A֏�~'=���n�vm�L���7p�cp�[Ǡd�:!�
p�1�8�w}j\|����ıcSLx��6#p��s �2���>��O�;؎�7�憎����w���Ԩ2��T#��0�v&�����%�/���@�����T�R%c`��g!_�;م3��vg�nF�@�K�w=Hp�G� ��!`K�p��'�ǃF@8^�zߠ����45��:F�=�H��=��K�#����:���I�+7�)]�A�b� ���W��:ҐNq����I���;���$���)xp�LVdpؕ��Cr���'�b%O:ڱ�Y�r�t���}w�{��~�+�L���"�h�̢v^- ��fdH�c��^4���i���֨k��6čhD��?,'Nuˮ���%�8fa�XcM6s��Qmm-�JӺ���9}RJ���ڕR�F=
gs��P��F.[`g4�ЬG�����N�l��j��>n';9�����q��	)\(~a~�z�D�!'d��9?m��ac�F�F�ly��C����{��� %# �(��(��#_˴f��:Q?�?��ƖX��n�|x�~�h_Ɵ���������k=I�� ��z"�s$�o$j�������y���|}v ;+65�3�v�U�̀��QN��b�����V�lN<�H�E�w�pP�COz)쬿�cwL��>��X�`],��<��:&C��㝷��D(��D���!�T>�-9u|�oX+k/\��϶�6I�d��<����O>��?��9�
Mq��_ =��.�n$�J�)��ɢE�dV{�<������ə�I��O�<-ǺN���S�i���WdY�t�����M�g��L1D@@��H��F#���@n�^���m��#��e����9��0"��:
H'�K�t� X�� T�Lq��5:��4���;D���6�f�9\K�㧕s���tN{�3�w<;�dj�7E[����H��?�����9��Ba�)�ӞN1��LՒ���j�Ŀ�M�-3T	�"�B��T&~���;(=W~MӠ�=���7U�0�X�� õsxw�s�{��|(e45�1"��-�XJ��=ʶ���^u(c<a�q L�#o������[�|�#�D�q�LNN��a���:+!
��!L�vFF���/�ɾ�����M���S]�r�|�u�j�Z���>�	'	 =��j�63�d�.ꈌ��yK'���=���9]���;$㓓Lk#
D� �(�����(X�G4:}ꔼ���f�Ȃ�c����h�6	�U����V�Ԑ�Ge#HD[͍����MG�>S�ȟ�rA�X���:��D�$b�>u�ѻ�)E��F�:\6|�Պ�+�U:�=��khF�"M��o[���*?���@�.�*S5{ېW��ᩦ3oZ����v�Ӂږ<�ٯ�x^�y�{�6������)2,x�=��I,E'w�Z�97ix_ͧFh�#�W�f5�؟�F�8:ɻϜ���3��gL�:>��Y6�g/������'��U`� _A���F�r%9t�0���Q�RH�o0�U+�l~,bJ0_��Õ�l��� ��#~��/!��d��&�ʉ�O%�RSSE�<Z ���R��W�H���ȉ"}	 �!uM�L�W��X4�su�L��k+HN0�v�����[��K����n�F��|�:����ҡ��<e�Bm�f7�P<�������.:���E]�Z)I>���ա�7o��k����˦��]�6]N�r�o~c�6@�ejQ&^ ����(3�N�C����S'O���5���R�w}t���Y�LE�qǭ1�M�اt�Q*`��wl-ނ�݇2�u[�R��?O�7�?t�c��a��Kg�4�a�5�j٨��Ke���pl���D�L��@ �a������`��H�����ζ��GZ;ڥ.��x��tw#y� VJE�#G\���H��O"A'׳PD#�:%�D6 ���p�1�������pF��$�T0�)ܫc�ⶠ��wBz��K]S�\q�r���J�ptx8`��Z ���<߰�S�\�3=g%��4�͆�#��<_��HVFa�}54DO`�����x���w�n�S�N��m/I�dR���"
T�RG��Yn9�}������uȩ�Q�0lk��M���g���|� ����Cۦ祝.��̴nؤ����z���87:fu�t�_{�Vy�;�i��:�Z����G�0�aϝ�"Lۿ����3�^�iۭu�O��M�[s<�������ۧjZ���q���5r��1Ϊ�9e�M�4���ANS� ��.���#b�G��wx k8���8hj�k���P�9�r�؜e1D6Q�pol��{�$9 p~x6@�GұC#���!�rG���$�"�-���̠�M��H�4Sz�9���
�"�t�<Z ���tw!R2��$؀�`�m #�Ʉu�2c/�g!JtB��q��K����{X���ҷ��ݜ#�:~\�_��ɸe��==-l�ld�mcp����9�$�W8� I�5���:$PI��+;�gf�c��\բ[ȃ"3�?���Mrv�
�� ��������9����-�/�@��j�=1#j�pV"����&�ZT���i쐿o���o8�3��ͿW�ا�w���mo�řj���1o6fF�ʮ�\�F��	���7������q�11��a{~6mG,d�~��U���i�33���r ���lDVpM1��h��襨�i���L����l���Ƕ����\�Z����Ï>B
ت�k����J��.��O��r,�]q��M��#�{/�_!eHs �������D,�d�yJ�v, ��fd�h��Q�k�(���w4^b���bf.�\��J�0�Y"�&jߧO��S]�j@�H	Mq�G�2�k#-X,e�Li6r�Q+dDY1]lQ@��S��5�8{D�)I&��W#b�À:xq���$�qw��D��#_̯�4r������7\ô�U�u����~��W� ���Fʵr��1��c�՟�ׂ���{�]���n�~�WA�=WD�ֺ]j��O�z���Q���^]2��l�9��L9�l�
ƒJ�dN���y��r<Cy�<�+��fA�d�s���Y�>�'o�Lc�>K����;��3���CfϞ%�����5��=�W\�U�ʜ{�����t�8.�T�T�H����Y��"X�8���X ���(�yX���Ff�b-��B�E�R�0C��4��,��7j�X��Y|��j��[���X@�X�́,�1��v8�QWQ&$���1@g4s�Lƨ�� �e�R�&{j��g�^�;����S���g�P��v4��+6˭7���qP�{\�E�g�KP�{��6�`���� V�����.z{m,`Ow�����������s'&X�b�Z�<f�m���-��8���M�䑟?��r��W�Ow[]u8E�'�1s��ܔ�ƑAv�GQ`�{�J���>hZD��d�ʆH�ϑz�t�hjó���a�����H>R��q�m6�Z��=��}�k_��~���}�WL��;��/r��B0XR�D�
9��~W�P��o���I�2�܌���0���2���I�?����b��Ϋ���,bF�F̑ޞ�(����D�a�?˺C��F� �I�? ���w�ٍ�TqI S� ���
Ivb��l�s�,]_'!�8W{��TZ����`���G-0C���`q�F�(�"�F��&����q<����˯H�0��������\�����{cS=S�P���'k3�V-cs�����,;��f??ޣ6�^/+�j�Ѧ;�N�ۺ�t>zkv���Lu�ێ}#O�˒:q��h�V6�&U�Ow��Z ����,\(�/��3�j8lz
�ZZ\2�M��|����x��?���x�\��*F��:G�N�v�����q'ҖI�u����]\�={�ș޳���{hތ�#��K��gn�����?)O�,�q��� Im>���W�Z��x��G}�5����.���ff��Q�T��1y�ѧ��--{w�bV(�#�ck��W =���a����MB�MD� ֤.h�M�DQ�����$۪A�C=#G]L#�8շ�
 �@���/�u[�����j��(��?~�s���Mr���JE�r�Lǀis�0��n��c�ݭ�"SɆэ��@x���S�k�%s���j�5]n��8�֣�נaw��y�o����PgF����� �~N�js��D��?�O�eW���HG񖜡x�B#5�T���[S��WSѷ=ƨ�%ՒS)}F���8Ʀ�#>[�<��-���L����^u��޽W�|�tP"�u�*P��LyGj�	>�s�<Q�vdا�MRZ+��%���؆F:��H�Ա��9%���&���Y��"���sD��?��t�=� ��ٸ92&;��l�2t싼��l�J��n+�<'Ƈu_�i˺W���dͪ5�O�t�$%����r�ߜ�; z`32��mt�Mj��>%������)�H8&ǎ���zF���j)��u#*M+����|7�L1��}�$`#&��q����,l��X��1*�ܶ��I}�H�p	 �&��j�X#�aw�F�`%��Lj�/�T�d�!��N��ɩ�6��k���uމɱZ�7�q�h�)\�[�|&��`;$k)k�( e�������9�{��a��[��ULu��Kܧ<�H"Ƴ�~�N�E��$q.�가4�f�ׯ�E��ə���Q�	qR R�u8����r�#� ^8O�D���Ԯ���R�.������@����c�rX�y׮]ܯ�5�j� f�恟>D>!dG��<6�wS����J�B���`�
���&�wKʅ
����}� �����_���|���(A9ޯkX,�X ���4��*(zH��{�\-��.��K3m�y�fC�`��4��R����)T���dG.Z"Wn�*�����7�|��t�M��;rT>���J��DP���Mxp�/X�� T_�H� a2mt�q���,^�t�������Ia�gsҤ�A$>y�|w��]�ݴ��u�-�LT�i�3���F�辆�Aj�>����cA:ijl�Fc� f6�G�X�k�~�]����Uj�����5lR���sR���Lב�5ep�#­SP3��v�OP�h��2��!�t��r�7����Wޗ���E ��N4��:8xA^�����5�c�:�)J麔i�s��w8���~F�`)��>�Fm߾��1��wz�p������k�8O�#� Y��~�3��鹦eٲ�r��q�h�%rɦ�8��I7��R��{�F�Ey�{�+O?����mT�z��z`��@lF��R'+>4�͙�)�W.����ˢE(�(h8���}銥r�7�}�= ��=$�E("�뮿A��%9z⤬Z{�l߹��tц%7�R8�|��4�>��s�=��cm	�낌�-�o����NZ�6B����w�G�?�l�&S�c� Tv��!C� &�rv(h�B��$3��lm���}J��:14��5�`���\>��� �s����ݻ�G%@X.��2���ˍ��Lq�s�?�E]~���3ئ��jHhJ
֤��������ʎ�F�����v֜��v]�t��=���i[j��=����s䐲�H��}ý�h�qμ�����y ?�g�
��$�˂��4Rn��'�1�Z: �o�>���ޜ���ر.�(��oP^|�F�ǎw� � F]|G�Α:1P
#�T_Aڿި�G�Ƞ�_kK�r�f�jY�r���Lʬy��Y��g�����i.\���Me�^Ku]�T*��;� z`3��=�!������d����p�*}�"f�|1¸��tQ��[HOH��3~;L���	��7��eނE��?ʮy,�	t�W+����F,#ŋ�$
49!z�0̚5����C$�hB$��M�Y�B0����,]����!��+��+;�a�O��uf�,PV}B�W�M[bHfnٲE�4���!0�F��f;ǭ z�c��vף��}q"��jyx��~�q�߭|����h��'e���Վ���dHǫ�^8�p��#��3)eֿ=�n{�D���:��m/���H&�Se;;oޭV(�b�ma��?�פ���կ~U������O��x�t����:��dW�·���e���Y,Z,���_�f��؋�xC=QP'W���H5=l�Qn{�;d�%�('�♚��!��I�B3s�Β����F�d�>��U��ĉ�)�j˯X�L2uxvK�v�- ��fd���M����~��h��U��[��3�jo�d�|hdT�.[!��-���)7�p�<��S���П9�+<�����K�N7Ȏ]��n{��y,����KϪ�Ar�L}����9G��MN ��"��h�Fw��DZ(�K.����裿`ǵG��#IDr�)��2�'���g�Q| �I��)����=zT.��i�T:Ip4s�.	KzN tS�'���x�l&aFƹb�ǟ�Gk ���������ݝ2�����`K$�&@����tV8;����9��<����^������7�KˆQ��Ϡv���?��4��Ș:j!̅�Mͽ��b8<.��:�3a�>::&����E�vu
�ώ�4� �����t�Ѧ�Q:v܏#jHS���R��ԣ�7����<fu,"ndm ����+8iL�'�`O,���-0�E��>�=$�ioi5Y	�.��T�Ӏ���V��A`���@lF� P)�.�q��Q?�sd���*��HTi�"�w�za�\8҄���S�^^{�Q���t�Q���/]��3��s�ɀFg�J�E����,�UE�|�h_<r��ޓ���V0��L�c��olf�`iol�X]Cc�`���!�huwf�}�x�jv����ǌ=z��|/��jqgz{��G~.��.�(LT�$�.�|����n�i-}�w�8Vb#�CZ���v�8��^/P���l����V�̰�95���{U���O�b� 5�ˤ?��$-8.4Õ*�.�t�l�ݣC��ܤ�^[���B���u�<��I�җ�ĬK8��:'���� �h�9z,�be�B���a��T��y��
�!��#���O�����4z!:�P��r�ӑ���lt��f��68Q�̀sr���́x��p���~���gz����r�80Ep#8���f��NHG�,��3tx�N)�&x_._)^I��B)���C%T�V��z`��@lF�p�&��3 y��aA]�t�FJ��ؐe�Z)����]��*���M�n5��?������� r��-����QX������9qJ��$]�Փ���j�e4�Mcݏ�T���t8�}V�"�88!�� ¶n�.lvpK�6o�O��ͦ7',-�1d$:a�pL����1:�{� ������AQZ��@�:]4�z^ ѩ�T	�8n��Hd��T��L��̠O��ٚ8J�j��?�p{�n��q���]S�/W-�l�_ތ�!c @p��B�p=���r���G��ڥ�&B��Ma���U��;��3��E`� k�8�l�9.eg̍ӑL�`�l��X\��A�/�9z�	���>{�~��]�0�0`T2�ڸ�օK��u�]'��w�4���^�\n�p�$��_ٶ��T(��K7_��{?�>�Of�n�[�^+.�K�q�N�K&�pزz�y	,��h�6#â�А��4������9�۷o���3���{wm��QFg`QC�q��Er���u��y�oQ���'���|JA��QnXLW2c��� ���P��:@?�pL���"�N�|���T�%��C����( ��a��s����d{ӹ�Q9i��������}�s��ё!���7P/�!S/�z���m:��`�mz;g^��l��q��(@Y�s�֧j���n�pdJ}mz��j�}�����&|����9]���8q9���L���ҋ/+X��]�H�3�az��[ء,*�5������{��H&?�{ȕHL��F��(A�f��AD��9����E��p<b1�'��K�L�d�]�p�1��A}}����;�#;w�$MKc��O�2�����#24xV�]�Q�;�����ʬ�=�^PT�nm�%�C#�2��#Ǐt�+/o�����E��̚5+ ��Ϋ�،,�;������߳�]{��e˖��d߾L�R�CM��Iu��#�������� H��Z�J~��?��|H�;*w�+��}F�O��x]*����ڪ��k�:h��Q�:I (�ʒ�� �E��Ns��)w� �����8������6G�2a�:��(�*|�H�[�T���냅�ۼ�k_����r����0�T�q3D�與sA�.�k�L�Ƽ�����_8G�l�}J�|:�@�2�M'���vְW;��p:�B��P����ϙ˿!��+N	�� U���o?Cd�1�|���k�S�QX���m��S�MXډ�����^�:XdAP+GT�U�J�<&&&�TƓ��M�t���������>�%K�pt.71���sTK&S|�~��{���6Ҩ��u�>�2�s�dꥭ����Ւ+������G���棛6m�Wgz�%��΃�،l͚���u�~y⡮744ևuݵs��PPG����l����f�QA}�K/�7�����K2:Z���v΃#E���]w}�MK'O�d��s�v9r�L���9���hC���љd� z��
Rf�����D$-y���-f��x��H������r�ixx���x"�}`�'�jmX�K��L���	ՀRd�k�W*�\#��a��Jfj��%֫�l8��(\3������Ʒ��uЮ{�Tj-�^�I���;�:�Z�ݝb]�����Q-��	�K��ڲM��I,�โ�ݔ L����#�>� ����FTgHn|�v��@����SR�G�(8��ut���ߐUI���2Ci}�6n�H����>X��T�b~Xr���,B!D�h�;p�����;٣o �e�ʉǍ޻����3��9 ]��2}ԏ�%�\"M-m<7�����+_�����>
�3�f��ٲ��$��γ�،Qƃ>�����;�⪺L�yYS,�K/�����$)`A�o�>y���_>��rJ���������.��'?)�4*Z�b�,_�Bn��z�^x����Iʂ�(���!g15UCˊ�6K��Q��&"L�Q���¡*�h������5kY�Mh䅮�ɬFkn��OS%G-���T����:����� �]2���l.��L�|�S˹�������o��!�A_�Md�2���U�	K\&�*�R��h��t�2�o�Ng��/�Zc^�@n��	���)��F8&jQ�H͉�Ӂf��h�.(S�0}Pq�	2��s�=�Mի���S�j2aF]�j������#�[>�ֶ6"���t��}�[JAcu��A��Li��pM��*	v�eӑ�Ϡ!���<������K1���Nt��~��~� �Q�ס��i�n�7g�<��S�h�"f������!�ՙ�3w�w���2o���;� z`3�[n������?���?�D�P���sh����}򔴷w�R]�A���Ȉ�4�"��76�"�Htp�6ٶ��E�@ #7>�E�f0�\��J*��HYţ�&�C�T��qtbPRuW�g�K9��+ ��)@546QU,���UA�Mc�#R���㧍��_�
�0�aH3*����uQ�sk[�46���
�7v����Ѳ��Z�@3j���㧍*�XƢ�×UJ��,����Kv��;[����&N��H>u�^�Yw�������#��g��D�quB�� �e8MQ����r/���9��`<6�ȯ�GC�ַ���Fz������Ty ϑ���X�>S?��O���g�1��bp#8$���"�N��G��zN�Ž��ȟ|�stB,l�ft�i�����
�MwO��y�O�����#R���Y�m�g��~�������&%���, ��fl��u��.ң?����T��K��a����4�!��ʕH���*
�j�Q�m+W]�����nuu���,��&5�uˬ�"B-�\�˞��)})���)b�����R�3�X�Ou�&�p����(�:�t)R�3��E��[)R�O��K��e�F1�p����k���~�\Ʃ��M� Uv|+xP�w�{ $��O{>�����i�sצ�aI\㹾���;��n����j��m�lg;�JV�Lq	}O�Qv�á��u|4��c�F84�y^I|��i�f3�a�d@F=��c:r��>��8�b΍D���\�~��c�2�u^Y��;�Ig<{&N��=��d>���F�q�6�:NU}��T^�;���v���y�l���x<��E/��wtt���475a���hS>
��Rɑё�lGG{O�.�}饛��~�[_�{?$���d�v^Lޒ.�v��z������?~�]�(h����cq$��
�!��:�������A�~;_`�8YL�1�vn��>��Q�=C�j�H�j��`[�jQ����g�ay���Z[����3�w�́�j���a�T�9�5!-ǧx���[�Ƕ9���Wya���?���<����M��(͋�C����]]]����)p�1c� ǆj�� 4� }����~7�a~
�zn��t��6�ՄT¦l`f�C��z[s�����3�W�� ���ԯ86��ʣn�F4h����U���w/\�hG8� Y��J�JAtB#�I���!��!�*��H��.�{���P��P�sL������̏^�j4�`�>9ǭ��7�V]���\��ש�/��.����B�1�#�w�S �,��;�JU�W��Y��W���¥�>�au��b�\i�F���6����C�|�	�D]}�1�X��x����g��u��*��c�	,��L =��f~��]�?��o|�k����������D�p��l_G.���N$	�C�H#6ԥ���)�;�k]�]lO�h�O@��!1Dzۉ����,	���uĩF$�E4���w4BX����ׅ
U��x�^��1W�
�x*�wl�Ճ��U���rK���w*�P%R�}T*јƈn(��ʕ��g�Rz6����D��.[�d�����*�X�钦 �D�-[A�F#�ʕ�Ys�g�����_��_5#�j�Ws�B��ӿ��.s�B�Ǵa�E�,�*t(��9,���X��{���o~ӟm��g��e��8N@�X`����y7�_5��<�C{�F���ϕJG�F���6V�t;�?6\��*u0hm@�;&ǎ�h(Qc���ӈ��˧�>����7��G��~��U�U�"Nm;�!c|�p��X�0�!�R������J��|�.��L��X`����kf��-͉EB���xn��X%o���Q��}sk��i{F�l||��G]�����'�P�&Qf3�&�ȜLm~ӝ�ȫ�.8�t|q��b0H�C�c]8�x:E�4R������`X`���X`���&'+Ԏ/M3�?������G@�i�CC5��4�f4.�+�j����I�[v������v�R�Nզ��H�X��gz�a��������P*��8$/K ��_b��kk�e�)��L�M�����cP��/�O�dR������CW��bӚ�~]=]���W:�CFqmz�}:#~�1 "��D"��d&!n(�NyL4�r9���5����� ��5��d�T\�V��H�.�!P�9jC�B�hHZ3F��R�Mgεy�r���W7���Qξo#u2�Y�ڪ%�)���`������ݶ�K͗�}�<}��<�t�q�5��{�- ��{����cc׏������;�hLfϝKu/�|A�԰�����z]C��Y�e��E��hH��}�Z�}��	Հؒ���s�U�]�a���	����8�,:�������S0�e�2�^x�#u��O��w�gsX`��f z`��F6�wf˱c�>s������-r��K��N��,��8�����N���X��S�H|���f9+"bA�Ε�q�)��W+�Y�ߦ)�ըk���-�ۨ���'�;`�C�>�dÑp�X��[�������}��7@:$��kb��kd���{�F����6]��K�7B>.�Qw�s����l ��E	�I��n͂m,���4жLu5~w�;yլ���W{u��i�|��m�� �棤y����r��ɑ��^s�X.����,_��^70��kd��kd�憇�\��7�4�Z���������"�����l6[� � ��R��Q�����b`�5������5�1ּiҰ���Ύ�Y	U�U�������ں�;;�_V��K�}��o<�_�m$��{�, ��{����}R��Gbh���8�P�
ʍ����>}z�c��{k*��(x�5:&%����Yـ�U�ZŬ[4�N(�:���z=��7d�u9��\�L?W��Q��/8�Nccc^��1 |^�6��S@�ONN�؎͞={��cE�t����X`����:���	}�U�<��������H(`F����� �|�cBg���g�LU�_#iVm�=��g��~��W�n����`X`�}- ���o`>��Q��X`��_Z �X`��:� �,���u`�X`����@,��,�ׁ�X`�X`� =��,��^ z`�X`��, ��,��{X �X`��:� �,���u`�X`����@,��,�ׁ����W2    �����D 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t :  � B�����`@� 0 t {uUcrC%%    IEND�B`�PK
     mdZ�S��*  �*  /   images/cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.png�PNG

   IHDR   d   d   p�T   	pHYs  �  ��+  *�IDATx��}	���WU}�=��9��HIH ƀ0�`X�������6���x^k��lq��`#N	�����4�h4�}�t�}�]��W��}�"^���Y-I4��]U����/��?�/>�y%*d�ɇ
�g�B�|��y&*d�ɼQȃ��$ɀL6#%�d*%	�"#��@��,�,�K�e2q�B��	��+��l6����@/#dzo4)Ch^ׂ+7l�|�y��'�=	��8�v'���42<�$&����D����fYK�I�0�l�D�?/ɚr:��:W���bP �d����{{���I�B**+�lU3އɰ� �)g4�Y3*)C�x�C�Ȋ$�U����J"e�#+J����YVT�٬��T��h�Y>H���\.�'�7
I�∄��EbגB62�,W�H:0����,Yrpk�Y��)F���s�ZX�`���}�
aV��<�J�0�d�(� �$h�3j
U4[�.���I���2t�Q(���s��T*Kߥ�;�P�v=}��BU�-UMe�'��4����lN$�4l��m44�p��9�N�������Y��l�>�$0��e��L�I�B�n��5�`+�)O���y��Y�pͅk�s�*� %���s��y�����$c>ɼQc}0�I�ɬE��,�"I�Y�!Y���D"!�a4�D���QUF�O������ ���^YI�|�y��_蘒����z��s�_Ba��C���Bd�����>#��j�)R�5Lz����ItWȳ�=�Á��!D�i��SD)�ww!�;J�=&i��0T�'D	ˠc����lk�� �b�T�N���'>�����`JnwN3��W��p;F�Kp�m��K�ǻo�����i�-�*�_���:�<gO�v�����sh�<�[Tկ�֭���x	�AF*�FZ�Y4�xǃ����0%|EP��]�&8Z��T�Y�p��N\RS��^�,f2��Ukq �A�>����Euu��c>}��z��
�XX���M���S���n�\X�~��+�\q�1��`���`����Գ�CI���r�C�����M~�������,�V��X���sp���^q�Շ���G�����wg����w��p<��������|�n�m#�*����	����U���>fYPӀg_x�&+�$ʊ�q����ƃ}�h�o`*�B�Yi��T��T:%>���l��S�
�-�/��ccî�҂��,k05>�5��lQ<>O�3������z��
	G��;ή�兗���=#��2��I���cA��I$�Q5A���V���U��"��!�cF�-ј����"�;�����cIS"4	�D�8|�~�������C���:�K��誐H\��V��w�K�N�'�PѰp	�v',d% ���VL����'q�qAͱ�C��VF.��L$��Xa��&���$�F�VÖ�ν�Ѕ�X����1�")���W��`�ؤ��� ��Ǡ���I�Y�A~�[.Eg� |3A�-H'b���$��.C���pm&���
��'�}DXGV@:��.��Y��gggdVE����LN���%��� 	���ͨ���[�?�J��T"�EW���aLO�`���X��2�W�a��V4-^��gN�Y_UQ�q_R���1l�(�� ^ӈ�b�����s_ɭ��5��ј�R����BJ�+�7<-��<��d�K�6�7�o ���#�矠�誐L� ��\mkkW'=����H�+��P2�F 5��X��9���am(���_���~ψ�fQ������.+b�\Ϳ�g00؇� �v~�SS��{�<�c~P�z��
q�������K���	��
���6��*Q^^��������l�e�K�3���[���N�?�F"��7��511t� �x\X+���Ʊ����Lk+]c�o"���'�xI���Ϡ���C2bq��Љ�n���0�������qb�cP�>���H�g4�B�gV�z�`���m.�+`-��,V�S@0���\�����L {��0�P�a���_G~d��_������-&��7����.]��)r�	r�L��E�4`
J+�16�!v\���LJ4[�X�%�H$���A�����ő��Y���9{EXE2��{a��E~������3��3t-'1S��r���U�%BY�L��
I�Ė����z�\RY����ӭ`4���]	�UX'�Caa����C�EE�!h��lb�/d{�gccc�3�+f�Y��f�2�����B:;;0�ϐ����~�xP?���X�6�.F+�P���ߠ��\T(�1����0g�L��AqY).l�)��t@���ⵑ(sVL�|+�-'���S'XJR�J�{�ɺ8���Ҙ�0��s�s��ش����#�a�?�B��PE���G?��}�LN�E����o�;��C�~,^�
}�=�������J�j��+`�!�_s��QgA��U����Aq;s�m��PyNY��Z��z��rhp�a$�-7l!�~7n����ص{o���փAo�U!6�j�"+F�"9q]�=4�V�-�F�@?�.�1�C0��$v�1Is!��`e��2X�X����s�:��}��4?����5
O��,6L�M ���`�ӹCO�U!�e�p��#�ۤ��;�v�����K����^*�¹D���2+C�eW��VCn�	b���`1�g���gr��{0\Y,��0�Mz&��J��T9t�,׃m/�Wށ͑7�G���������C�s�ݤ�b4ȱhP�(+�YA�f$GK�ee(�(�!AȖ��I��ҙ��Fn�Z�&��l�Ă.ʄ������(RN�,DXJ2!����٬�jl6;
���~�K��/v�PS]�@0�*+p��׿"EW��;�[�r	����㥗_���A�/\���L���؞��CXN$r�9A
���b̕�h�o+O�PWs��c�\F�_lA�VT^���>��7$2�`���8{l�\}.��#8�v˖-#�6�EW�Ȋ�gh��_}~�����-������D�&`��')2b2h%���H[��Ա3�c�"�.�)-����/������Ur�w�g��r�X�r���?^>vR:�֍U�k��誐��H�������3��L�7���wv�UP�a}��*�#/����<����r
%�+�s�Ba��ȅZߴ��ʐ/�.�qJE���;�E		���m��N�d�㍷�b����S'�E��[�e��ѐ��3������&�0�lg"�G�΢�4Fb�F���^���%������+��U^^.����+� .b�<dE����I�y1W��X�T�����3�ԗn�ӦE��
aX����*��O�=^m7>8r��k���%����HZBFղ�i^���`�m������ʂ8T�����H9x+��O��\���`�F�18�O�t3���PWW�k>q,��*�z���?�	�]28Lxm���z㞩��>������q@�����P^�΃j�Z4�d2� � �3�|�bQs�sk ��@���f2��H�S��=������]o�Bxfm��1>�G��h�Ǯ�M���zq'c���ci_�YQ�@
��3�|���%pY
E�GEe�R�\>*W� 2���[��K�dr��?� �8(�e���e6sQv�7al*��a�ۦirRH�g�S��ȣ��k��V�,�1��.�)��t�'��?���@Ii"� F�F�S#�k\*P���N$)2^XdB��D��J��a.dH��bk&��VH0�����bQC��3m��!�E��z�-ho;��k�㲍��܋;����;�Խ[�%\��3�3Jmm�ܲ�k[6�d['�+��CeE
��������w۶aÆ��k.�� �(�f��	YIKHr֖��CZ����D9?�Z�X�b%+yx�Oo L�[e:���i����(v�Swf�o�=������y�Oy���)"���)1serУ�d!��~��,4�=�I-_��!JG��
V����33WI�N�>���Ĵ�Zv�lNli�\����)�B?	�c0(f���O��S��}��o{V��ޢ�B�����d���	'n���y�
Jʱj�:T���	fDI9��}��"e�Yܹ�h9�Y%��ҙ\բ�s��֬���d0jۼ��S�e��wq)Y�g*�Ν{0�ۍ)�!.�Ѡ�|�G�f�^�-�9d#�����k��/߃w�݋��D�%K��� k��ġ��tٕpXͨ�����ag�"�V��WA��G�q6�W!�b��&@�&�F1��t��1���_(�1�_�	=�ڰn�������J�����n�z��
a���A��H8�<b�<�Ņ��񡴢c.?ފw��K3�N�Z�Q�
kQ�(Z���ɞ$KR�l\N�V��'` ��V6����E��'֭���W��m�8|�0.^�H4%5-�(���[tU���D]m�z������-JK���L�<**`t܃���	�W���7�Z���E�n,$��[�V��0k�����:�k?�eK������l�&��jCS�%8q�V�\�}b;��|�\��uu��&�~c'YU
�z���a������v�0�]�L�s��Y�AV�N+)$#�δϋ��Jb��f��7����,����sx)
��h!E�g�A�Zڻ&����C�4�GØ�	axz/)/��=^
���o�lv���[�߂��b"�c���y�Ld滍���c#����#��&���ܰ�@?��������q�\���2�Z��|f�O�1&�����s\^�(��u"��&�s�k�RS��U�c&r���)�2�hi`Hcc��qa���;�^��-��7>��n��V;|��z/���g����ن��
��Rϴ��4EY\�`�dGlu;i���'���h�[�� *f�H!��ϩEc�4K<�Q*}����"�"������ٳV�O��=� J˪���&�Z�ZJ�/�*N�-�.Ϟ>yJ}����A���^y�T�]�إems���s�k��$�!用j�(#��l�|-��w�X���G�SbFQQ!��+�p���*���{�"II��_ǒk�5k[$N��-�FY4C}�I5�mWW�]�ށ�
�
��bT��D,��K� ��v�koΕ_��(f���S�YY�b�<��DB����B�6��R���,�z{PXP�(�F��S,(t������ÁCm��ýRC�E��L�044����R��NDbi��_`Ś58t`���ZP]E��b�X��kڪ,Jzĺ����dr]��Ė�"N�g��O'㈑��-f�"ڟ�U�f �SK�,'h*�����Q\�������j�ͪ��?I����ޢ�B$��5����!����'��,1��' ��;08<B0f��bCm������H��K��}V�u؊�Cz��3�3����ӗ��X(z+*v�h�t�pf����y_	�F�s��3��[n��	z��Q��Ƞ+��e_}����HS��Eό���EQVY�<��(W>��]my��/�n���oa��{�0��V���������JI�.��e"�I�D �px��]"�M>\��!�`d,������n����Y���Xo�ׇ�����%�y�m��g)��:߃�j�=y���(*-C��U(��k�1Q��lq#��v��FSm%�6+<�#G��514�DB�j�����p�c��$.�Pa&�&���k�Dج�ϊ��M���-8s�����z�V����WwHK7@o�U!	��C�j]ݥ��ի�|�|��?��] ��ru����}9�������$X�U�2�]���uxg�[I��>.�&��B�]�E���"��;;��\*��8Q�#�J��{_4�VV�c�@��+ω��>�'y�D��Z�z���;���?&��X������c1�N��o�q����!�>Wp��]m����)Z
��)ֲ��^�#ַ�D˺��U���������"��z� ����0��/�����Z{ǹ3���I��O ��k�����Š��ˢA�s;T�ק�Rh0Y��!�Ոĺ-���х��6[P�e�U��>L�"0���wZ�5�/H$�p:�[n�
�k��sQD|WLT�4-Y��L�ߎ"�I�}|��MAN4�$kQ4�O��r&���4�.�ҫ��Oi��P��.��#��څ�pd�^��3�$*�ax�BX��P�'��������[a2�p��Y<���zյ�tU�oe�@������@Y���f�H,Kpv�ͷ�p���^E�4������Cx�w�<�o�������bH�X�Tc:�2� ��T#�M���H�&� ���եy�&�vY�=A�`�y�sW��*��A���VBza� �B1���N���>+������v��P�oބ��a�,�艏GBŹ�!�Ҭ���uR͂j�-�󐆦z��|?����D9g:#���v F�"2�ĬO=�ȴ��Z��
�za9�f�h0;�sG7���㉨h -/�j�Y�;r�(�sb����N65aղE�A7[�q��8t���z<���ff�������+���6���S�[��!4��ĺC~���� d&"lFQ&�
��<��O�D~!3>���I��\�����a$�x��a�{?fg���I�Ϋ����E,_�\� ݟ�MRt������qW.@�+���&��'�A����^�b�1<�GOO��Z����c�`� .�R��0Y���_�F�]T���TޤQZ�B��������1���P�[\R��#G��n[6,V�ݙ��l��;�"*M81�ʦ�Ŵ="*��� �܎�*%\��z�ƆQSjŵ�n�ٶ���G��y%���Գ�/�W=Sb0���"�`s�5�F3���҅�p:���m���L���0F~�<>��%豹�f�Mљ�"�]XB>AFO�y�aŖcu�(���T�W�(���E
��֣d!�Q�^��J�5��b��-�l���4?{��-��_?%��7�X��pth�c�)�M�"p��c�����@�߇rʳS>
��t?��7���&����gd��,V�l��K%�()-���^'gE���� m�^�*��+]������e��eJ,�.���@e$����y���0C��׏k?~#���S�MzE%�������Ս�q�XPP�鄑�f��K�!��2�nb�I��s�.�u ��@
�6�ESi-m�����{���ʐ �rin��M8z���ct�z��
i^^��������>�F�����_R"v��%Y�ق��2�T�#��)DFg�{av�!����C��s�<�r���eee��skCw� 9�$��JK�yJ��s����ˤ133�[n��:!G�PRԀ�U���;X��	z��]�&�˖�O���_|�E��`�lU3IX�_��S�Lx��xQ1ƆzE����a�K��;�q�>�İe1�M�m6}g%��b��ň���o=��e=Y�⥍��酛,����#��ލ��?+�j�����?�=�R~^��AoѹrQ!Rl|c��{?��H&��c������D-)J>C���clM��v&�2 �@L4��j`�;Ol
�~��������|�X�5MX��������z	�����)��B$'&F���<���&g��WRb�FgїJY�!��|�|�g��$s��u8`!��H���
ь]C��]�Qb�ee��s �>��x���O�[��d%f����Lb�#���s�OV[VE))����E��L$���gPV݈�`������؀����<��-, ��[tUW�3����H�ml!��©��(,-�e���Y�;.���b�S��������0=�\O7�t	�8r_!�"	��,�g�߲9�(�iD$���(��
x�Xl�������v9ɏL!U�%(�d6�IE�@wѽغ�� =�ko�����j�K����ZAs��5S'�AeY���2a��9�Q��*�ML�.*���h�<�@P�%h& 2��He�h^��+���&DW���kP^Q���ދ��>�uww��+)�s�>C���d�׈�
	�m��d%G[O�Z�G䣵�����}H8��b�N�1Idp��UB�e�(�Y��q���!���p5J�L������0���4�r8�P��$��-,)�bAV�"�9fHF�_��������]�qn ��PLV��#�Ȑ�*x���q͍�»o����d2�����ɒ���R4-]�������F����t���L��]z��Ѱx	�.AQq9�ɲ��Ӕ��a��{��q�q�팀Ы�������C~'���'����z��
��#�H'�R�D�Z��f���Ǥ�z��:-c��C�ɡ��;�׃��j,ij@w�X�����ɓ��n]�8^��2�mk,<8;����s�g��Cl��w܁��^d���j��ڍ$L��op#���^�()5iR/��$��J
2�:ڲ�k۳"�$���ϋRN�x�GS�	L�n�C>�OlL3C���!��7R ��1FS�)���TTV�v���X��NؒLf+)�����E�����w���Ь����5������}��ܡ(4��,�儢IѺ�=$-*��`ݪe�����A1Y�a�2�M����4pє�ID�4D��EY���xR�_�w����.]��6]*��"���3�� ��Q
m�zZ,!��7�u��0>r�����3=�u
�E�M0���<���b�k_���b|��G÷�wvR$4 ���z��h�G��K/!�RaLGQ� X#�w��-8��&��1T���p����=�Fi�캵�4�!G=�yY���]m]-��b3BD����P�h9��]&�u�V�����#r}C��ۢ�-F5��}���;&Db�"*�ɽ��MX�t�	��B�o܄�1�)4�?�w���n�/��&�m{_��]h;�&�	��ƆKp��	�����wcjj�y����i
����!@��C�O��8|�R��3?8<�]���]grZ��^��!�T�[����Y<A>��_��|�۳KXΕWl�G?�]���V�o��;^����0���Ά�~�J��a?��������:o*S��]�TU� ����12�CP(��a�pۭ8r�0�,������}x���E3����~�,E`�R}�%2G�-:W�H�g	�����b6�U�MK	�:��F轃|	��(Y��#	���_w�Up�c��}�!���$[T���Ξŕ�ՕU0Hx㭷p�L;zz�(���n��F 3q��,|o}��y(�"e����;����h=u^r��[���x��!�غ�����Y�u�})���I"t!:�L(-viU$̘���:D�j��f���p�R�	�<���OR�v

�=��S�3�"!is$`(7
�i�F�,2YZ�*��r㺏~�v�Oљ	z��Q�B�Vái�����$9v7ʫK�.r����]��6�.��Z-.�`尲�n'zη�F���sD?1��{<��r�=�Jlq�	��&e~�W,P��Ef
��k�k����J�t�"/��MJ]n�L�_������)%�9u��S\�XT����G��GB�bwn7 9�˖���b�f9祤�vV�UN۝�s#����D"���U���ʒrr���W~�h���G���	�lR0� z�8��"���V�F.������a7����b�~8x\_(zC��4���2Q�;a£�
&�_���]	z:�	�|(+)��\x���LL���XpMϣ{`L�{=z���Z��?�5�r��U+��
��e��7�wI�=��\T�ޢoE2�]���6��?}�0Z\��u�31���^:z_����=���w���#2�q
m�;���e���x�����s�k��+�����W^���E����������5�c�uå����P��gX��l�`��&�,�X�b��>�4[/r��6,h��?8|~���~#���$a���e��L�11�%˘��$���J#�D�^y7l�^�i���IB�[�9O�	[l@<���ᳳ�t"������Y=êb0������	�ӥ��,������Yu{fz6�N����Ɔ��[tU�wr�f���"o��?5Ks���:�u;R^A!F'<���1��J5�,��BcZ�����i������_���l��;� r[s{h���/�����nj�l��_�}���P�%��$�ɧ^��u��3j�T�ɬ:x K֛M�����یw�~Gl%��誐{�r���o��{�L�r����h){�d3�Q���C�wj: Be��j���פ���X_/� x�xl��\PQ��}꼟/��V�%��Ǿ;�܋/Sx�x5*Ii�����l�5�b�zIDEwomen���oJ��Cc��W�"}rח�(����޽S'����~��_�O>�\w�w�TY�M&N�KiY��V�*?�S<�-�t������{�݊�Kq�UW�?���]v��#����IJ�u+)C���Z��#�dI�?knc3��ͳ���9��]��(�+���/���.�B�|��y&*d�ɇ
�g�B�|��y&�(��5�N�    IEND�B`�PK
     mdZF�i~�  �  /   images/85e66502-362d-4a26-afcd-97fbc4859675.png�PNG

   IHDR  �  �   �lC   sRGB ���    IDATx^�y�o�U߹�������$��$YÓml����ӡCU�ؖ��bl�iL7Ch��!@H��ҡ����Օ�*����ƃl��,����7�������]l� ���٪�{~g�:{��k�9^�   @ h0���m�i�   @ p^� �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   @�����^@ �  ���  @ � M ����q�   @ ^l �   <TU��tYE����^��}�w!�   @��J�����s�Ҵ�1˒��䞝��_�t)��(���EQ��8veY�eEeU��M��$��yQ����CKK��6�%?�}���v?����|���   �<����}�K���f?�mw����˭V+���]�v��p�i��s��%x%|��4s���E���(��^��q����o<}�ռ����o��+� �W 2@ ��_��[���r��p4��<��N�'q�z�~�eY����n\u���E��(rE��5�k��*��*w.*�8n��[U�$���<�'���Ao����>�W��}K�����K@ �  p@���_�-��o�Uu�sѠ(�YQT�4I�0��W9�+W����]7����v�-�y�$�Ue����$)�$��0.�"^XXpG�������?�.��	 x�|F��   |I��_�g4�LQV��Ey�fi⽲R���\�f��v{.��������q���E��o�����)�Aq�ī������������ر����7��!��K@�b!�   @�/H����O�]W��8]��&ij�Zye�[bZ�\�W1���ή��]9WV�%����%ᬟ��z)���j�+��?�}��C?F5�_Є�s@ �  �	������sQ�3�V۵���b_yA"�G+D
Sp*<�BcUY���=7�\QN��*�g�6x|��g���������������/��g�   <�~�g��ue���v'U%	^��Z)^	� �+W���Gn�?t���%��*��ƉD���UY������i������O,-.��7��۞zN��8!/����! @ x�D�ϟO666������8_�Y��>���O�x>��\��\��-�4���]�WB$�$b%x�vw]�Ԥ�]Y.IcWv�ݨ�q��eY�i��ǎ͏�-��Mo���=g4^�F��;�ۇ   @�Y#���oM��]�g�������J++�[�9�F�ϟW2��t:�{����?�c���'��:�v��z�8��,��r����4sY��7��w��ļ�u�1_���t+��^��Kb7����Ve�����r��v�E�o�c���]�۰�9�   |�Ο?��Z{�E�B�f��|���v#�W�|>���N9���۝͕7r������,͞|������yy��j�ť�:q������ͦ���c��N�m7�繉_��*�-ސ�vX�:M�s�,M��`��xÉ���~�~G�~��@ �@���mok/,LW�i��ҕ���������#��d�L糹sլ��~`^Y[;�@��w�4��iֺt���.J�?�y~c�j�+++i\{x}H��\
e������W�{������!
m�	l���u]�!xzu�.S�n�[�r�/z���G�-�Zs��J.@ �������[�&Y�����;����,�LƓ��S7�F�ao6����Y�n��w���7�tz+��kUU]lg�Ս͍WW.:[�r��vkG����g�4�{+�Z�+��=�ԓ&�����t:���N�c���^>�k�@b�9�����۝��go>��7��/T���}� ��wv�KY�2n�Y̋WN���E�����^\\\*�����gY�&�I����\�����x4�~o�$�t�8�tUV����v��\�ӽ<dۛ�������!��u'p}@ � ��D��ߛ-�^tn<y�x<���h��py\��W]���p4����|��4s�O����;n<�Q�$�����y��Y֊WVV�����ʻ;�͝�f��Ӂ���=��&t�VW��+W���UkPȮޗ�������u4q"�����G��P���O�'O�x���w��k_�ڃ��4���~A^��q{����׍��o~�'��������f����jd|
ש%���-t�uUI��p��I�<����ʭ�rqi!�J�,�r0X�vB��v�p4,v:��u��^w���t��j}���>2��W�vze>ɟ^YY}2I��<o���gS���������@l^�   <	�{�ə���O�:�����[���O�E���4����b����իW-�LUN�V��&әtC)�!�mY�q�jۿWWVܑ��\UQ
AHL���g��w���-,�x<v�V�b|���v:9P$    IDAT� �,�G*[潻����W�D��=s��ͭ�������*yra���ӹZ���v��x�b�WY�<o���'d}<��{�wskkmoo��Ҭ5���Z�&I�U�p8r�N'�9�Y+�]�rcGiQ�&���[\Z,u\_�ݎ�����ڪ���,��,���1#�Q����m�M���T��f��oQ�J������l:�������M/}�ՙ^+++&���tʅ�������Ǐ�g��~���=L[�F����WVv���S��������r��v���ne����Y��?��y>LӢ�nz�����"�����S8o_�`?`n	� �{�ϟ�wv�3���;z�h�e�c�?�x��z$����M�3w��I��[ZZr�/_��]��������q)A<s�<�.q�O��y�&TC��Y�0w�.^t[��nqa�zݎ˲�'��J^e�� �l�
˵+.�Jl�����dmm��G�9��N����s�X���Ӂ^���t �4�İ~oν$.uh�����H�n��EY�Y[}j>�(�>��葅�ړ�Ї�/�����|珟�p��?�r��=�����MA�k;�'�ټ����Ι�i�R�v�]�}�����6�����b)����d:���=7��}��JFVJܪn�l>7a[�2&��d�Y�SQ��N�k���iZ������knuu�mnn�����j����ZeY��.�:u*�Wݓ<�Z�i����c���h����`�O&�X'&��p�ot�`�߳�$z��,�*.}���z d�>�=.{ݞ	q�S�Ntɋܼκv��c݋^�^�T����^Y�f��dF������q��[��tsyiy���+I�&i�'}˹h���o��t#���V+ݟN'�s��R�jR��EQ,�ǎ�>��.T���է?��ꮻ�:��x�y-������'@ �+I���#�N���J����`�8����v'��/ݰ�?t+�+��j��d	��dj�Q�P�C�+W����b)���[_d����|,׬�E+K����{衇,�aia�v��CJ�0��z���Xh��Z����y>��������[��x��)�,��y�/�()#W�
�H�Ԏ;�.�.��\�Ib�9˲T�7L�����uUmggǴױcG.�v�m����~�o��7>o�x^^�����t��zW����p����mi�eY��u�ťXbLVb͋��)�a�H�*�@B�o��ޣՏ��p�9��� ��ܒ�˵u�؛/������$�f���î���rww�l�[n>�cms�b�����>[;��������ŋ�3E��F�$A<�ڶ�|��m����4-�BטO�q�nǭV�&�=h��4I��`�����d<��ՙ�E)�E��_���q^�Y^j=���3l��������ի� ��q�^��N�]����:�{0��u�45�����X���E��w�� b���G���&��/�L�3�3����ask�?v,�\�u_�~�V¹:3�S}?�ά����5�8P�&q,���VҠ"Q����'��L���8��ι�(�v�4fY�RG��h��neq_���v%{eYΒ���&�YUӪ��ը*�$)��h�P��~�·��jg�_--mU�����_�����B�! <D��{o����Ϝ>��˗�������z����z��:�Lb���敥�E��ZN�1�淽=w��	7�L�Q������l�Ξ��u{}?�ƾ�B��n��]�$6��G?j!K��n<�V��U���+��%�� �噕Ksߣ�>�>�яh��G��[�P�2���\�H,�l^��j��+	N�ҿ�$��컍����M���������}����^�����:��ox�w|����ϼ���[�ο�|t�䅤��^�ۍ^2�L���y�W�A��i�;*�x��1w���|}}=�`�v�3�닲��8)KW�Q�>�QF�3�*a&���ֶ��4m�BQ�����ڪ��ԋ+]C/}F-P��RBp4�'TF(&����г#*���ʵ5Ź;��㏧G�������1x��5���WU�T�T�������b�V����G4���s{ �7��Ua�RK�ʴٶB���ʕ+q0p㑭������ʲ�}H��M���<y¶d���IH�c��Z&����3��*P�P��J��mmm;�b��tڱ>�(�r0Xt��[��G��>��������7
�7�?���l�8�@u���o�k�>���@�ϴ(�W}�ղ^~%��{1�5'�q)��i��$I�V�m�{8�b#AL
�`W?�z�� ك^��E��;-�n�e��f�ҖP�Ӗ�N-���R���T�����.ky��#'�Γ$��I:K��*��b�JG�r[�N�ZU�[�Ngc>��D�w{�'ՓD�^���YM�v:�|ҞTyޟo���[����?��-���ב��� �U��c��ϴ_z�ԍ?�����{{��c��</�K�/��hT�:uC|���k��ֵ�aG֎�G}�bs�ɕ�G����op����m��`��;q�;v�w��[���o���3<��g�ǎ��jrE�$�(���L�8�����9y~'#9�z�x�����"�S�i���j��	��<���8���)���x�}��h4.
�P���W��y.�q��W�*}ӽ���[����|V;�Y��W\�J��������t�k⸽v�ʕ�<���9�;����<�&_���M��nG�EbdT�;-#P@��R���a��y*Q���WJ�J�9�f�.�L}/cԿ�ʑ�V������[X�l�*��L�x���Ϋ�q�J˪���"�2F������g�'�\�����^�V� 1���'�k����� �%�������t:��H��</�Y��(��(��|�Y���]C�Q�~�@Mxű	u��ޞR�-��*�Y֭�Mc"�<�z�$�CL����l1	Z_3=h�	2O�^z`k��X����~��?\bN�	��Hp*�ٲS���ړeY��Jh�aO��G��b��s�(k����C1W��_���`b���n�+�mca.Ea���A<��e�g�I<�LM���m���8��j�!,�� <�v<��Q�*�g�@Vxz�_,X�N�mJ:e�ZhJ���N;�X0���]n<m���n��'IR��z�,}<Y��6��T�N��}��B˶�|\�����z�(�~ͦ���w�\�W��a�n�&Y֚��^U�$��dY{;˲Kq�\���b��,'q+�fU<rU9q�V���s�<Ϧs��ؼ��/�D�����f�w������,N_�4����s�>�%�{ݽ�ޫ1���r��g��[����h��o;v��w//���ڵ��3goi%iZ��?�_z�u��	w��E����*���s��Y��Oژ�9L���S�np�z�8y���nqq��r�6����2~֘�'Zv���K���nr����D'��#��o�:dSC�vU(O(�Ue�����p�������[���e���c�^������ǡ�	M���Nq�ߧ��.�(��2�����C�;������������/{��O�Վz/�������|�D���t�<[K����=��mnn��j�o˲4Ue��gϖ/�˕x���(��mw�w�~���cy׹s���R�j���Tq���}��]��v���f�Ф.�'�p��U˪��g�O<n��.Zy>%����4��������n0X�Ѕ#G��	�bd,�ǂ�͓�U���塔���SV�`�`���p_�&�e@P>��o%h��{�Kصfa��T�~�C�qQU�,�$yu��{-�����VJj���DĪ�Al$̵h����HyFm���
f��ĸ݃��:8\qOzpB����c����Z��(�Oq��u�j����ġ�E}�~���g�<�A$�����-�������B ����>$����ޣ>�Ng�]\\��]��P�Oy��¶��}�]�`P�Z��]}m��X��7�`��a���[������	b߄�y�g� 
B����ص�5��xњ�G`>��Q�Ċc���R5HB���w�w�b(I�c6�u�{~��\}�lc�\�O��^���L��u�waQw�(R=�:^�`1P{������󂰮���Y�{t�����Tv�ݓ,K-c:����d�¦{�#��e�x�4M��E�4汋�.r�8���$ُ�h/��^�ZmM����*�QU�q�W�عj��8je��s���y�-�E�ϊ,˪��A�yUe{ډ��I5�v4��c������*M-77��8]�<y�ZY�*�~�����~xn��|�����'/��/�G����y�`���')�x�j%����N@�e�V�B��l�E�l^鼩Y:�#v���,?������z~llͳjEek6�f����:�v5m������|�1.�k�M&݃{o�'Q��~�錿@D�8�g��c��=��iԚ��Yke����i�<�R�·j�X5!���������[U�5�Z���Im���޷v�I�R�w�q����+��;���R�����(��s�>]��U>���"��O�������ޥ���}��_\�����0���[��l�����ܑ#G˳g�Ə?��m�klO����[M�nnm���������ܹ;�r?,ϯsG���J��]w��Į�Q�V�Ú�m�w>s�V�}�c��;n�����7g�O%��خq̋l��k~����ˢ,��͍�7~�7,o��U9�v)��[اnL�'Kg;d�6Ԏ�0k�K;̃镩����Nݍ7���[�'���?�귾�>����W��_1�{����d2�vV;�ѵ��8N_q���{����$�B���q��m��f�2�������-w�q�����*��N�(vS�T�˵~���9���P���x��q++��ĉ��Ť��j]���/_�l���_���K��K�/�Օ�R������|�ķ���N�nu�J�^{u���V?&�%:��[�Cj�=;�!Ճ��]	3�W�^�I��ջ恬's��lIgϰ��m
���o�V['���-.zqP����gW��z���G�j�Y��D���e�=�M��o]O��5�Щ��{}�Aܒb�l[Ư���Z9︾\��8`�;KP��ыm[�>#Y\$���������@��{�9xsCY�0�����^�\�O��h�h4��}j�S�/!����(a��� �O�6(�&x�vc��z#a*���lץ��y�5��Ff#zA*{V?*VZ�݉�^���>FK�J�hů���P�Z��}ɓ��B3����W5��^�o{�칲�K ����ņ��[5��mmm����g1pIl�9O�&�_��oj!8I���Bb��kaKݟ�]��w <_%�j���p�/��6�\������a1��e[��EL�_��'+��Tj��}�cгE�_p��O���Z��a0;�b#��L�DY�}B�j�\����Q���;��p��v�T�bk�S�0�:�Oת&�i^�y�β|6���N[�e^z�}���X6yQv�=ݺN��z��W��'I<�YY�8N���W�m��2/s��)�ٝV��Y��iEQ�ɪ��4ɪ�|j�5�Nm����J|�ԒoK��~'OY�dU�đ��(ɋ<+�"��?�1P*�Q�Ω�S�F�%U���W��_h9��/�Y�¶؝i��/�K9`�|>��H�V��,J��2b�<��yYUc�dY:�NgC�[Wj�5�Og�B;�v1�N�Y�M#�&�y1��,�#7��|��'�M�v[;�U���·z�n�]>�fUU�V�vUN�]Ͷ��Z���u����nlT�kk�����������(�����ҝ[[����;�\���?��C"^�(6~�����v�l��*���ޮ%liӘ)�A�Z|�Ue�sy��qKZ;z�yv5�v�}w׋_l�Y�l���	�v�l���~��x�V�A��:tя���_ph�_V[*U��P���z׻��K�]n�~^x������o���wm�o�՜�-
�|��_�x�	�q�j>��oz�7��{���?��|���
^��� ����%�I�:�:�.m�YYy�'_���q_+k�yɋ_�:y�Dz뭷�흝R��&MGj�g�%Eɨ�=�ʋ�.I��ڲ�!���r8�Wɶ��c�T�,T��f�<��4W��_�'k�D����i�[�u�%��cǎY����j*������7�x{s˟�����߿��d8&�wv��U�����20����`���i6��}� ��B-�}�\n���0�G��n��~���3�;��*[�eR��8���ݛD�ڥ6�-v����7ݣ<�>�IIj�u���g(�3}F��8H��is��{R�G��Y�ф��&�Z-�Z�r-�B��/���9t�~|=n�D`�	����WՁ<�p�1�����&s��b��$]j?����D�v�YɄ
	M	b��a��~���e�j~��*_��B�{BK��b���bD��gDqc�~�@1�ynI�O��Z|�m�+Ժz�7Q�P�C��r(��=�~�d5%k����=3�=���B�>^9,n�s�4qFaa�(�a��O%�la�nY��`#6I$�-$�u����F��]���v��vdG�NH\Rey�N'�΍���ښ���l�]��P!3z��;]�۠�,���*,�$��@��ؑ�m��@-�F/y����A��g4��ł�F���P�y��Z��,w���Y������Z��=��6�S��z��[+ܬ�yf��~K�'�J�q�s��K�kl�c���|Ȕc�M��g�:���F\|R��r��d@��q��󂗫��河��cٵ�#I�E�Ï�4K�{9 t�zqe����um�H�W�D^��|6׎�A������(�?�N&�Y�a��R�9�N�$�4ǖJ~�L�~gS�d�����vi�g�i�)YK�Zy��U��gu�^,��t:1��������9��J��J���*�~�j�QX^]��4=�6��ŕ��Mr@��Y����ͭ�B���Hĩ�L'6��eY�'�����f�r����</�QU���t6�t:��l6.�bE�$��8�6����h8��,i�:Y<��I�����D�@t�n��St��ߚN�?t����n��E�Gܤ�+^����c�{��^w���R��Vn���ډ������S����#��$�._��n:}�yx��N���n��X��q�9�ͭǇ�{Y�ƒ�=����[-���V��a��9*���>�H6v���/��S娢P������'Vh>�g�.v�~�ؿ�Nfx�un��H�$��ċ�;~ꧾ�;X�������k~���
�_��_�>��ϦKKK�s{�<�W��u���x4������0��VN����KV22��K���"/�*!��5���K�M�u{�-�����hT�J��<y����N��iG�N^��e+��c6m������(h ��B�Y� �H���e��zo��;ku:-y}�;�t_J\�
H�OM��M7���8���V|��&MF*q&Q�kx�n�A59�^,����%�D�y�Fc[�x��� &t:����'i��������=�A Jh�E}�{�0�6.~ҲrjÑ�z�R��)�L���D����*��� �T>E�v�s�G�c�uj�x8�IT"�DW��ja�'d�S�A��jF��%�)��(W��@<_`A�{��K�x!`q�
��g���l���-��V��]ha�#�*�d6	\]C�ӄaq0���������U��M�g���t?����'4h�$��=�~�֓���0n\�n<��^�kBTv'&�d�ŗ�/�Rۃ���p�P��4�Wx�~g���Z��N>��8f�~qbBV���~�� �k�P'o(�Cu(}�H�B�BF�ۈ�x�{��_���O�p|��-O��I�+a<�aW%������a��g�o�w�W?��{v*��V�~���|�^��>��/��4x���Vq��{_�ӿ�;����[���� �-��(��*�}��d��^�܅�	�-}i$%�&u�?���^�_����E�����?�j��Yy����yĪ���u�P��{���P���;��Õ\�;��kB�����eu��o�d�agF�ճ&�	�pz���摐��2��v�mI���)+�:q
�    IDAT����Y��z��W=O�N�Sja�C��c&,p%���aGF�=~A�j�&ZN�w���7>�� ��~��>1J�� ���\����V^�r�Ǳ��5����Va&��v����;kA���S�N���-s�h���!ۓ��!J�ʗ�;)�Jz��*��vR�zE9��}v���4����I��2/˲�&���ӓ�d�����V|��[�����;v��{�k^S./-ǿ������cv�k��B��ɓ����Vk���f��h�ꩧܙ�g��ή;v⸅4Y;j����oq����������OBQ� <�����w��ͦ��9�<WoW�}�zhṵ�e�h+T�*��/��/���.�s�.a;;�^>�Z�Z�_�@��x�FXP�vy�k���{��SU��������������7��q�ϩ�}���M��^�S����֢,�-=�ą�������������a�N���$�bN4�����D�]m�?��S*� �mm� ����z-�q���d237�ԗŲ��YH4@���Q�s�����Ah����Y�vJ��g��ì��O?�t|��q���W,NW_͛�Y�����+p7��(��2��	sm�j{[�;?H��M7�d"[<�:��f�'O�D	m�	���4��B��o��ګ��ݑ�O�l٠���'�6�מUMn��U��~�^^���Ԏ�&�ڳj����:T!�����i��U�&L4����щN���$�x&�U��ϼV��ZE���յڛ�aZ$�dGj��>����(Kk�a��[[�N��ˤ{��).K}�'3- �	-1����O�Q���D����q�^o�=�v�L�:��EJ��'�N׽�>m�V"��	�d��V�u���G6MZ�2�{��	���݀|n:
ێ�y��Z�*�#����l��*�����8� ��=�0�á3j�1��5���:$�� �,|C���	���>R_h�!��d�SH��5+5���	�S�|�1��pr�eJ��|ȅy�����v4�{���[����N�_���eĞ���h�@m�݅�L��+���/T{u������Ņyլԟ<��4c�,�<�/��������3Ʊ��L���El��:���Ś���K^T/���v��ߛw���K�Mg>!5xHâ���!�%xyU�%��aW(0��;"&tK+8X��z͹1��'[(QY_�k�Ì�B(�v]W���˗/�Yc�8����cA�	�^xK��yAs���b��
[�XZ�{	�4�T�<�د�Xc����;����x��ֳv_jvtM�lX�����}~'G�-�k�)O�2�g�JI�*�?A�����gX���C���ة1G���X��իW܊��,1+ɕ�"�8�Z���Q��i���D�M/�23vU�Z(�[�}�-KKK3��j\�t;�B�&��U����s7�xS)�����;݋^t�����L4��\<��Wd��SO?es�^�B�ҷ�rf���:9a���ٛM�j����v@E��y�t���k׮����W����ܧ�>#�>X�C�hüb��`W���z�v�~���=�ȣf�g}�=��{] �:$�����P,�5��-�9��gϤ���!�?�O��~����;�ę���`U%}���ϗ�)�S�����篏��ߺ�����)}������%3i%��U{ȴ���>g+)J��	�?H��I.CN�$�V��gӀ������L���(,�O�B$��+w���vwwsy�%x�W��͍�:)Ǘ��Jy!�3LD�xJմ��
�taKO�S��&ۦLӃ�^�/-Kwd��m�ol��+T����ow�.]2���J��r(;��VĵU���ζ=L���[lҳ�ʺh��*��cڠ�Й�^���:x�o��%�����Sf�AK����,�����R1����@����1�A�g��C<��,����%{���?�~"H�7m��*���`[Mcl�EV�� ��PIh�y�b][�C����<��{�h��P��A?�#�~j��@U�Bp�n��X��~>���7[��4��w����-O��c�v�b���Z=��}/��A?��M"Iό�B�>�0��޳n�
e�v�dbq��;�B<��U��S�E���=E�'��:�Z�n��A�t�-7Y��{˽w��o���DK�|���$̐8�I�����{|���[��x������>��L
����gܷ< ����`������ɮ�����/�� d���:d���{Y�7��u���/���b^�_�%b8|�]Z{�$��,���z�+g�>a�ě����}�R�����z%ԭ�h&��%�h��Wي-0�0"�OϺ��: İ�!o���%�󃒑֤�;���(bK,��� sbԡ�U������^{�C|y�M|�bB�l�{��d/�b���5,D��Z�ڡ@��BK,�B�d�I9�l�\Ϟ����|L�2�C��Ⱦ������Ʊ-f�i��k�{��3�{ް���B��V�Ǣ��0�Td��[B�G��6�~����#�X!/�|8N_��>�ּ�
]p�^�m\�p�k�n6��If
���׳��������h�Q����B��Z��L���C�|�����A�$�l8�4g�z����bg:��
)[_?��O�~؝8��������?���VsW�3g��m�/v����'��+��M�	^�5��O��PL{njի늙�;	�GyĽ�k_i�Q���^���L,��r�n���,��������D��x���^]����=�P9P���a^��E�9�*y�˳7�U���SO�Ν����u��|�7h!2�#���v�&D���n��҉�_���~i��uC��}E�*4��O���._��޻���O���&v?�яzO��оjPTb��?aF����m�۵�&��A^��M-�g2)��q�j�q���O>�d);��FK������@��'6���ñy�?� t����ȑ#��1ඍ<�"�J~[Y]�%�����GH����uْ�5c�˙�|���cs�V�a�NBW[�2\m�ϡb@%h��J��o4������&�u��䁓a�_6�E����U�	$}� ��������y�*�V�I:��%0��+�V{/���D��K����\��O�yh�~����v^`��ĵ<@��~����=�uHB�h� ��lb0qh����:	}a�ǻ�W�P�,5�(���O��!�A��{��V�ru&��!�q���r�?��>F+�;�\�pѼ���b���Ja7:NZ	�����먅����F��lL���^�5�t���'ݹs�,3X"M�y��	[T|��pǏ��lYM��{̾��J}�c�?�^w����>�s
T�DL�uY1�Iμhӳ�����?N>L�{�CB�8Y�ϡ�-]���S���>�W��X��ｧ?�0��PB,�y�,9�{4�ת=�A�A޶syX��K�:���{���[�_(�v
j���g8�ə�X��xe=!��J~�P��~�8����x3C�v}�p��}�u�"�\^z����m[_���P'�p8�~/�u�{��Q虰�x�"���������4O���q`�Z*t_�����R�E��q0a�g�3��� (C�Ex��(=bX������{}^]�Ǉ��~{�5O�:�]Wv��7����ٝo�	Lg��U�C�tȑJ��H�w!�"��汷�z2��K���£�5��>��':��%�`U홗�A�����M��V�Sdi<���Nz���C�B>,<��N)��3�ɤ.��żBq,��Լe�6�� &�ލSm��ص�)m�o	�v�]��/�X(���}��ti��$��*g�d2��:"������{�|����㛿������>����,�W�^�m\;�U��F}�X]h�����X���7���7�t�U[q��/������~���_�2i�[�<���۰z�`�o-)ܞo�{#;�Ї>�~�߾ׄ�6�j�Y���K=�>�~�-�Ü)[Ҏ�W�WYy�K�.���U9�W���e�ݶg"�)�nA<�O�#G��+��O�r���������}�3�������9�umƕ��?}�K_�-o�ѷ/�G������Y^�:�V{JVS����2�+W.[�ݰ�J�@�z�݌\�x���gY���w��]�%�]�pa��'��x�қ�$���y~tssS"֎��jz8Z��:�,��z���g�ɤUO�*7��	��`�K�	m#�D	��%��[�a�P��젆�'BH(I�I���Q�v�A��_�X�G�'ݿVg�:��]uf�	��}���b�>�&�:s]"��V�y���P�A�Q��W����4��j�ı�C�_��g��#�����?4X�3�U�2���mnnF]'l����8�Y������^�x(G��B̪<���t���AI"L�f��2�s�}�ٕ�<��Ӗ�xmc�^D�ٽ�:�O��"L��<���9�V	����j�dC��hP����:�m�{�%����}i7Dm�HW|�&�n�5� y/����c���>C����c��� ��#���؋�����v�Z��=�.zo�����a:~B����@��P�j��'zI���e�!FU�B}�Ŕ��W��{O]�:x������۝��A��a+7� vW
	W�'�{>�Vs��>Z�;2E]ø�&�V�]�2�����>�&������Xz�v4��D� �LI�݋0Ä�yur��s+��4��r�>a3��p�R�0 M�����-�\^�:V\ai�CLX։MV�^������8n��8��]{0}ȄّF�"[��"�	ֳb��"(̹��i��{aK[������"&�b����	�ד
���l�j��]?\���y5�(�T��؂E|½(����y�1�:�w��g���%��b��*(��i���f�ĲU��Y�hŪKR:�u��V��|�,_������l!�z�v�Be�R#ǂl_s�v�R�6�h�Q�v�4~*LO}l㴅:ڂ�	1ǡ�;���J����٭vv5H�8��}�Q;h�[����}؜E��j�x$����I���/%*Q��~�aw��Y����n��vw�����׼���D�e�0N�/������~�m���*=�q�r`��-�x�=�!�浢t�=����_��<�
��s������Wi~������S'�������ߖw���x�Z�j���㥅E��`�MyXu5��̦/}�P���������{_p���~�m��͵�s{-�A�w]�|�o�����s��N�k�?�'2{��[a��^W�^�%�|�5��t�n�����|6�t�8��v{���������?���ċ�;�����t�TU������f�7����^4��u�8�M���E�����z�`�*3����A����Ǣ����m� j�nirz�
M<�� �B �8��S1�*�&C� ��!`�=�}�Q;eM�C̪���VW��:���I�<��=��^M+k�7�z��~��hҐX���nw���Į�lR�>�O�w��V~в�k��Q
=xv��%`���0����Y��z�V���c�g��e��M}�Ŋ����y�ud����i��`{�δ����I�[����������I�\�SB�&��Hu}��{����'9L
a�>q�Z���ާ�k�6�S�	L|e?��:��W�~�[��~��WF��
�I�y��(�'~���u�و8��$J}�}��ڢ�+�T�m�r��bA��[�V.��6[���n���o��be���Bu���-��Wu�{8�1�>��Y�v��������o�9�'���q$�VO�Y�CW�]����L�#�h���u_��2u���xӻڙ_`�e^��`������O�����S	�̨M���)��3�m����K`"ӄ��5Aja^h�f[���F(QX߷��m���01�1�!8�9����=�S��	��&�r}R�����;�q>\���5���WL�O��]�L<�Ƕ�1(�"��ɍ�$�:�ل���P.J�5����B��a{c�A�G��x�=q-\+�j����#T��p�:�Zs�v�B��ƌP?��-KK$�)��V�u�;�o"�s���*{O�r_$Z}_�C�B�����>B������IY�܃0[8�B����ϗٹ]}-YUX*��\UL���iU�E�ƨ�W��Y��zs��c�Y����7���-������p�b�yV	��!&;�����I��m�m��n�ɓn2��յ5����k�í�`%��
 A��m��c>�w����`P/f�ck!Hv����.x5��I�-
O���w��-�|%�~e���
�/���e!����w�����ʝ?����?��}����p����1d��0ֆ�����p�/{�ݿ�W��M�u�ó��}��ߝ<��7�y~�|>����;�$�s<���vm��m��򖷸����v��g{{[A�*�*~����o��gΞ)O�8?��c��ŋ�nͲ4�?y���x�����?﫡?^j��K�������v����l�X��EQ�M�7�ey�,������"/��"��y�)��2L�U�X+��v��C�a���i�mKiwo�\Z\�A4��CB�hH:��D׬=F�B��-�C��X�~n�o"$L��]H��u�t�zr���ղAP�e�֓�ek��3��$�=*=3�M���b2UZh{g;V�j�X�O�Q	9y��`���W;8�N���E��vS�r4Y&t'vh���U�Y\$�4X��tm�l0���>�Ė���� |������/1?|`G*o��uyֻv���)i�S2�&U]��>�5ē^�����MVqDO�)q�W�PuA}��ש������u��~��{�������~'���kK��vj����$�c��y@���rnIo�F8�D���xl�Fؒ<��jQd���'l�}�~����Raj:�N��A�!(����Hq�:�Ӌ6ُ���[�WI��vG��Y��$%�~N��Wo��Br_����ra�~nq�
��L���l�m�y�$��*�;��hѣ�$}o��u�q�>�Ӯ�
�[t�� ���'a��L�䅟/�e�H��ض{
��2����I=��8� ��sۉ�$iz�.�-�/T��$Ϻ$�a!*n�zM����PBc�� �C�Cr���-*�m�N%FB؅��ק� ���uBN�<���M�-����� ��m�R/���z�^�g>P�[�����`���y}5���vT}�B/,`��aa�� tCIɰ���,��-���Ƌ� q�*E�C�܏Ma�/�؄E���ױֲ%�ݺ�Gإs��{�1�w8Bl�?�����0���b��m�3%��l:�-X��>Y�v]W>x;u�V6.���RK�Yj�<��z�!�0P"�5+'�q�ۿ�;lN��?��n4�q_�9ݗ�=������U̶Xh��SM��yr}���=z����X(���w���'���ͻ��='�ˇ?�Aw��;�j�Bj&:l��N�rԵ��\Z��s?�c?f���w,��6������p|�-�?C�V�Sc����?�G6�������t�����:��q_�u_����5;t������Znye�<}����[���B~�W~������'��}yQ���r9/�Ţ(�W�\�
�sébſ,,.)���0(F����[�F����+���X��{~+���_�ۭͥ��O��.}oQ��>_���k�]�]*�Fky�w8^j����n�+�j0�'K�8Y呢(��l1���i��̦�SyY���|1/򥲬:q)%��v�ݲ��|��n�b��(N���IT��lނynɚƓq)qy�,�������E�|4ZT�V��Z�R��G{L��v*��7��y~�[Ž�����i�qQ���h�/.,��N�D�&)/��@����Bb�2L@u��	a�VP�.[d��:�p��yO5�k^k�ߟ�Uonn	���>}U����H�V������5��3��    IDAT�'q)�Q��r����Wv�&����PX���������C���Dq�ڵ����kfξ�ުM���jwz���A��h�0��T�<�E���u(4�q\{�ԗ�_[�{{�୦�� �<��3}]��`啔=X-�y�7�v�<�q	Y��2yu��B���O������N���_�
[�����(��{SMt���bM����]ً��*J�a�G_1#71��>dM�W�i�V��uBdJ��RR����	� �\�����v$~��
�
e��!��x*�e"N�]��>�6�	�i��za��p�������DT�(�B�%�ڢ��A��8��5��mϺǐ�瓖�(�t/���0�@�Fa���0����Wտ�3�1�۲�P�-�<�V�d��|��Õ!4.�8n	Ͱ�o�_��D�-@+�~�?G����U����S%�+xB%����X�m��_B%To�/NB2�Ć~�qG��}�̓;�}�{<Ǯ�Q6�*a����-���*�s_&R	����R�������&������~�����
B��c�M�-��sѱ�Z{���}թ�
���1t�`��
�FJQ��$��h4����ߍ&&/׈�Q�DAЈ��RTC�u�N��w���^�1��gC���H��O�n5c�5�?���?�^sɱ�l6߁<����ٽ��z��&�=��#�o{��s�w�� �f<�p��N�ѱQ:15mA�ˎ�S{�ҩ[��xF��������իג�����hFU�s�)'��������dcp�@�ə�m6�PnUGf�H���BQ�e2w�Z�dC�.��2f�?�	x�5dKQ���_�4�;��A��O=Ų�ۮ��� _��ivv�9�X[q��}���d|��ѥW�� ��W}M�Z{_�Kc�K9�$��J��7=3����պ�kQ�C	��Ɨ/W�o=�'xS_�����j��-�c�:2qe����՞��뺻�����^��n�6@���'��|��5?�.tw��F�U��뚓��.�N�w�$���4YM��Q�t]JiX��Wk�M�>�,g�h4�l6��Y�@K�`R���9�#@�D��X���P��q�����bҾˑ�H��._�w㔟D�%��}q�j��"�ʫ&&T�=b&��_��3��9ڶ�`�
*��2�t��LX��� b�1�N~��Ȕ� �
�
��e(�4㈇�l@i4N�^��b2D�m,� 2 �Ť�4�$� �RRF�ͳ�u�ܸ��cLm����:�&��-�[E��j(8!��UI�B��4a��bF��`��ƙ ��d�)I�?�ĵE�`����4�x-�/C���hA��s�[@��m�C�T��H��3)��{�^0�1�7�j�Uin���4A>��eH�� (��2���t�v�@�
�@j#�(|��Sݔ�4~�����B[�c|�H9�`]:��<m��(��s�����y�9�ŏ���}pT�d3��1� ��	I�c|��h�D�qS�a�(��~,����t	��8�+QV�RiFcZ"�X����J�D�ؘBd��.� �
p�9�om����l�:�	�9�S������z�(6�z��i���'JC�?㬆S6A��q~�5��p�q�Ԙ�?4�a��v����u�i��6�1�$À� L�8�(ж\��0� H �A;�e쬢���l+<X��h�s;g�F~�,�_�CqLZ����qM� �q^Y���	��ctw�V�t�e�q0㡇�#G��=ŵ��##��Yͩ��"+��t�t��={h���F��h��M����bz��J�����K)O����t򺵆&�m�m��"�#߳4P�{z��=�^�Bi���KH�g~����xqN�tw����_y=z�G8z��fh��1z|�ڼi3-[B7������b�r���[N�r�Uk޴m�6S��m���c���7��߈�dU�ă�r�� �N������l�ru�֭*_(�X��+�i�����$��>u��r[`L��уC����8���d�߼ꪫ������{������f��k���������\=z�YN��QRq<�墿=T� dP��=��W(��$I���f�\G'�II��q2�l6� X�CݵZ�����g�z�-d2�����r�V�N��,b�@���ӎE���l�hGʹ����� �X@D:�X꤈Ns7*ȳҢ\e�C��p��3�Wn�X��-}�%��w���>𹙼��j�|!��i"j�c�57`G��׆�E�Z\��ڂf#�:��ϒ|%�(���B�, &4\�N�E�Wu<ϒ9�ET��q���ǿa��ŝ�`Ҩ�@e6����-+������]�\���(T1ϝ�,��Dlq_�-�	w���g"����\��GD8�iS���Z��+Y�!����=Fď�
��(Ѹe�
�)�8��c�D��9�Fc�a���d$3"����i�(p*���%׾��t�i�!� h��J$Nl�4���a	(��J�u C�7��l���9�XXę����� [�k��� ��gqQ/�4W����~�,��q�Fi�4[ިP&�`�o��I��D��Kj#���H8��]Ÿ��K� xI&ׂ{��5�^�wzj�����8O��=6�=njp��Þ����(:E�1�97�g��A5@\ L� r��Z�A#������Y�j~+ �-�F�nV �s�B��]R���1Q��5�y�E��!ٯ���	K�2��v�c% Pn�9v,Aej~����gG*8۷og�P�(� M���3u� w�t�z�V�Ɲw�[�M��o�Hh�f|ڸq3)H�q��E����}���E�֭����tp�`�B��(.x6ca�!#C��7@���P�M��rn5�ez�H�ϲ·��|`���_�?[p
 ��4148@_���<O�q�t�_7L#'�Eψ#�522��_�������2ww��/��u�֫�8�K�����SSp= ���1��B��.��M��P�
`�Tv��]]��T*N���-ǡ/._��;۶m[���;���/�P�8::����"ʋ(�R�LV�� J
Q��@�p\��]�rǂFcyWO�x����LO�J��oƥ��2J -\��I�Y7�7VC@Q^�� T�v�(k��9�f&Il8�
�#)d𘮀�]@/k�FaZk�X�#�ŋ��n@V�۬�:�[C�(0@8�"%���V��j-��s����� `�c� �X �hS
-Q�d�l�BA�jsw-���=�.JU�����p3ޙ2!<nȈ�!��H��\��ɴ((����51(��b9��/�Z�,�	E;�P6��1�e"ͦ9�|�d�h�<�����Xd�0~�I�ֵ-�"�(��9c����I�8.RD�>���+i|�!H�����(����������=�,WfWY��&d l�� �6�� ����� o���Ie�c�l�	J�d���pі{#���Lx��"P�ӮX8��[�U� qA;R�o�L���Vj_�����>E%� fӍϯ��G��Ǎj5�@Yʃda�L�v�9v8���R�䜰�Y8�ss�,�%t(�|N�8��3�+�W �P`	3vlL������N�c��F��Q����T*\��U��7�g�mb���B7��8�.F2�.]'��	+�&���@޶m7�	�1�8!��a`{y��?y�A�=�u�Y���*R.\{�K΢rw�ܹ�9��>8ppl�F�ڽ����~��d$:��q��=̩�O��Rd))�r�Vn����m����ˈ﷾y�]������"��Q�_^i$��Ҷ��4hAMD}�#�Ҙ�������$��Ȯ|�6L�t�?���"��CC\�=2<Dw�yk��t����u4�b^4�a&��}�}���q�Ҁ��A0w�B��$�."rr�N�ayy^X��
�B�b�
�e��w���U��v:�x���������=<�HaB�!��֪�Î�>_,���7��xa������	JT�����=�W͹'N$�^�h��T�����@e]W��f�,U��hl��HGCI�i�9��F�!6;
��A�aA�6E#���ʂ)IP,�E�)����@���)�d8�*)]pC����6c��l���V��*�qQb�j2��pÂF��q%�U,�~�"#rjd����>�V��*_[&��
^h |&j~(����8.2���!�q[�-Q��h/�%�!I����av�%�`9G���2iRP%Qi -5���}����	�ߓ�$w�s��Y!dx����f��qlt�;;�R\����I,� 7 �5 �E��w��!�g,� 6bo��.B'B
�p<����,w�4z��g��p>�7�C����lIQ����(�dQ-ʐ�NH�؇���".��8?�A�3���a�n��G
Y4�Q� \h&�2c��X��}�1��QN��@Q-٭�0�Ծ�Z�����Z 9KC�2�UDI���
���9�:� �2�!6��
�%��.6��YD�%c�6��4�`�̩�L�g�E�h.$�yD8,RH	�e�z�y�Y�L�ų�j����1.N���t\3�
Md����p��8@���m�-7��E+���[���-�m�Pi�����B��؆Zţ�-[N5M���ݻw���]Pl��:��s8�g��I�~��'�������v�߰��(�=u��-*gU�PgZx�9��wҚU+�l/׮������Ym�<ԑ ���j]�����]GO��e;��A_��[�?��C{��}6ҎFK|tt�~��d�\ֹ�M�Sf\����0:�a�ݰ�pw��Y�H�qS����W���|��۶m32P/���4|���홙����l�a�����3HR�����ڲ�T����s�qN���Too/��喯����%K�T�X�K��]�F���)um.W���o}��p��]v,��B#��R�=�玌Ī��7�f�K�j��u2I=ȇaҕ���j���h*9�"j\)��Ѩ�SJCQ��fɀK�<��5�x�Ş��6�	�.B0�ZL`[�WC��].R+2�zl�ִҙ��� �� dtr�+$�2��t��&H�!J&�a���/�I��  ���J�� �T�s��m�"�6���cQ��#�.86"���p'�(�yƈ$��(q@���/�R,�(�Ĺ�8�B�aY�/�J��D@ �� ��jժ��2"|L�`�R��I�d'�b�k�"��ַzٰ�I�ǭB3�8Hq �Q"k(�d��3�upF� �*ԘΉVZM"���}ʽ��6�� c|�o-� �{dZٶ��)�2ET��)�b��Y����Փ���L{z��J�ml��1��8l� j�41��F+d�Fb�����@�����2�H{�Z�q] �8�D��N`
#��d$��x��~�(�:�n�� �A������q� hp?3���p4}�q��W�_�0���$�viKmlcim��L�z.�a ���F��?CxN}Vw������y�F��Ғ �?��r�ѱڷ?��g��̰�U+��nQl޲���>�%���ldd�Ќ.�)^��كw��H8�b9��5�WQ>zGJLW�)� S
,M14�-Ow|�Nz��YK:�IwG�;�L���,2e�K�Dq��O���5�\��433E����l�Y�����N���@��?>u��8ԥr	u's�֟�t�蛶m{��/Ԣ���Pg�T���&"Q�N� a����}���������	��k_��ڻw�i(�G�g�f�Z��]�v�=�o�b>�1�r����o5nng�X�c�����t��ܩ�(���W
i&�t �t>��b�2��
��Q�YiECav+W�DQԭ�����(sss^�\V�>�2B��dy(�0i\�,8³��2�Y�GS�g�!I!�r�'NS�h�%������i��E�������sM�� ��\ +�OI4`D�-�}n�NX�ܷ�_��q��U� ��yJ���F�`�s�x��Q��c���x�ϋ���������E�
�m�/��[I�\�iD`:�=m�е���hc?���*X�*�����t7$`-o��N(�_|�.,�?���1c���Rpi�Ϙv��.�4��5�[�_�"L��k�����P_D��&Jk�D��k�'n��%8��4���j
�&&(�H�[��]��4���mw�l/�Pc+l�A��ka�j�j�Dl�����7��}��ڗ8r<���&]�n;\�	� c������Md eB�0��#�I-�A��f�c��9�ڰi�}�1�s �����K+W��@G����G�+���}���QM
na��k���?�7�m����a�y
��/�⢺��:mKg ^pxW�\���Q[n!l�w�7���B�������w�G���o�k�f���v����j�?ae��k�m�1�P������M9��j?~�Q:p`?m`����/�2=�ē�y�YNA��S�[صq�7��uo��B-p��~����v�|l������8*�Zz�zzzZ!�r�S�ի��G��-o�C�2�Su�}�� h*�	�^ !ɒ�͑��g��ɹ���������r/��;��X�c��� �?��O{�n�����; ��b�����x٬�9.:,��sc{A�\�\/St2�@	���>�SCNJK�T�8F[�|���4M{�8�@_'���G+X�Ez�6�E[�B��P�"b���z�j#ij:�IT�F��i͙�3��ߦ([�#Bq&�(IT�6lT���,`�st��h?(9,�,������3��H[�֒:�-����"@��ٔ��n���DG���RR���k�[K��k�g���g�0 �c3���yxo~a��m\�_�ؗ\� �g�����ب78��,���)�^�߳6mp� C]��m�L =h{�$(��wbS�hfl�5�5)�o�J%Π�8��#VUD(5p��G=6y� ��d��+�3�\4����F�d/��7@��b^�D�\�t��5�p��}��,\�p��]�S(�՘�n���X�N���B��m4��طs���@KPC����=s��e�p���~�X��r�͠c��N>)���{= _�s��@^|��t�w�Ӻb�Jڽk7��/����Ɨ�s�x�}�z�Z��ҫV�a��p���-Y����yp���d̶�CD����{�T,���U'�)�o�Ŝ^��YѦG-�b�� ��#�0�͍t�%���� ��{��}Z�b5�un�t�k^M߿���8:��O���e�^���P����N�z[W��˶m;�B������Tp����]�f�r���GC����vz+��ԛ6n�ӳ3�E��b��:��}A
ixx8DǛ���(�����<����f���ڵ��/���u�;��X�c���#��<K(��=D�w����g�755���\�U���T� �=�O���A�G���8�Z��(*&��Nt<D)��qܣ�.%Z��Q��Q1
#�+f�|	�h�R{�-WR@$�yH�-��s#� ;����q����J9VN��=є6;�X|��X!t�F�� AC�k�9�à���*�%Ϥ�m�N|�����l�8N�CY�)��7	������~�Y93\8;0q��J�v�,�5���p  0o���Y�BX��42]tX�"B|���-_�����ՑF�WtŲ�,;>0�� ��&��s��x	g��0l��e���kQ�,Ks���#tM3v�0-��_�K�j7���+���Z�.���Ǳ�C�d�5W("�8��7�@��R�B}Fmڴ	:��������e�����w���vÆ�t��ws��W^I��w�	P~���� ���o}�;��_
=��NZ:���8aJê�k����:ۂ<�v�C�����G ���u)�DS    IDAT)Xù�����>�Y��,3	Z��=Oэ7}�9��
-�Kk,�D2�ٿ|_���|�Y��Y
���^u�JVg���_�+�/��O�qjg7��x�>�e,�-�#���uۙ�Nz�+�����s����gsa8s����Q��p��A�~�RQC�#�y�fDmibb�=թ�i�����⊕+�|>�jqh����D�Xxd����f3�ޡ3Ȕ��۱@��ǰ @��w��˻��{{�R��LNN:��7P�9i�f
�DU*�!j@��#
�7�Bܤ�
Ji���&ITNSg�qh��8K4�t=�I!���8U&�!�V� �FҤ}�U��"�)&�k��1�$	��G �C�ܵ�-q%Gl"��:X:�I�k�Z�	V�F��-K*�e�L�֤�h�h�0f
,v�2��Dy��2
��{n���h�k@?� f ɼ\�� ����6S>�\���h�f8�F�(�e��'�VQ`��X�l���"�U��­�يV�s�Y�]�[�'�08��]�/ 7
4��g"`.��Ç��A$���/((���x�RQ]�2^kÁ�����-�n�M7��^�*����D�W^�Jo��}��g�I7�f��������_��8j~�9����w���n������z#�$%n<�gQ<j
5yP	������qt�Tȷ�hL�����xl�e�F���� ����t���7h�n��rP�����Dt��+��o�S2�}�O9Ҽ07G�~��p��. u�v��I33��8�����Ü�B ��p���㴗����,�u�]�_�N�j����x�[��/I!;�a����i�ӸB�5XT����{�n]�ꢾ�^�A���zn\.i��?66��\ד�^z�!u��:�X�c��~x6~��' ��MW�\ũ�Bov6U==�E�g|�O��a&� ��E�<_봜*���@F�Z'�9�l��a6���0���N}Ju6b���Z�$ ���m��������B�0E��`D��t�4%0��#��{�U��qc��.hh!XY�����R���B8�`�B#��~V!]my4�x�2JN��v):Et�z�oF7J۵u�3w�h[�h$��r�����#�x� C��4th&�^&�!���C��C$i���Y.B;~b
tJ=42�N�z��׮����Ϡ���raa�n_��ӧ?�i.�:�sSC������g>��֎L�l�@�s�}ͭ�`Oњ5�(��wP��v�	K�f|��xbGw����)��"�����raG�5��TjT*wӾ����چ��q���ӚD��N�X�b������ p�*x~O?m+����w�#S�_���1Rx�n�}���d��o��������e��ٿv]�/<8 ޅ���u�r�w� �{zj���{�r�����484����#:�#<<�����5%7��}����c9�����9D�t,б�z��"4����7���Nw�s~݋"���mz��4]��������n�*����䂉�U9��0��g
n�Y˸����~1�υQ�#'�d2��8��:N�J9����ϓD�w�DY�y��h���Q�j��d}��G�<��Q��6��Z-��a����8�>Q�t���i��u'I�$l4���?����.;iԛ�|!�L-��xs����޾�l�pх�L�K���'v�B�� �ڻo/�4׭[G��'��:��x�I�g��/у<�Ō7n�Nk���z���MR*�^ ^r�A�q����R�C{�즮R��"�� ��B�¶���V����nŊ̥�(��hph�����1�5�FŃ�ö���q����۷r��hX�4��;��;\pרU����FG�i�[hnn����hvf�c� Ƞ�p�j>��]e�?8x���z����x��''������(ʙց �kxOU"~.�^4#<���0�|���s�kpp0���R�uNPJ���|1�����^�tW�郲�:�X�c��:��-�\r�%~�1������w�K�8t萪իt���>�����˖-�cG�ѓ;w1W-tQ̶dl��NLpdzݺ�h�S{ό������L��E�+WQ6��/���H�E���}��RW�D9p�S���a�F�W	�2�_C���s|�j�A������̖�cѭ)
��X�	�Vi6������^8�8i����uk�Ү'�����Z�n-_(I�̴�5�p ��_�HM>�G�n����B��Z=�+����f#2GDs�פ76n�DK��ӑC\�
PD�!@����Р�`�RJ9sD�wV�X~�R�[���������;�X�c��:�X�g��ygo�rpd��s�9w]� =��cMPW.��B�'�[�j5<p�*�ˎ!`�Dr!�5;3K+W��Ch����Rf��OP3@S L�e+Vrњh�t���?����Y�`ux�(l������h�_���2>���v�~����[��+^执�Kb���y��㼆�`��I�j�ϱ�߿��}��J�֮����;�q���Q�����<c?t8Gt|o�Ÿ�
��������޲m۶�g�o��{Ϲh���?�~ff�=����C��bQ�*�h힘��7�󱣓4�t��$���/hӦ���ΝL�.�(l�gs�=��7
ݟ|!�n<�u~ӱ@�t,б@��9,��׽�ӳ3���.\;<<J;v<�*S�|�+�>�Аb��-��G~đ�+V2g���+WҡC����b�
zj�S��h�4==�T��"�;�l9��zZE���� ��8`��o����(��Pk��*<�Fi b�n>�z=��+W���Uֹ)wT�����O�t�!���\>�z�+V��O��'Y��𡃬Q���`����d��&����B�h�z6_���w��m����������W�f/�I�3=�M5+�@��\�<�
�W�a�8>�vD�ќ�W��5H����uk�B�-v�Z�AW������(ow��:�X�c��:�X�y���/9�-)9��7��g~�J��6m�{�<�@Q[���ffgi͚5r���㓓x�FG��ѣ\�p�l���@�^d��]��I�hB�,��h:vl��8����/N5��LdW�9DiA�(��8��Q^J]��E�����0��t42x½5Ňk7�>�z��^�:�"�VْFCT�X*��� ]p������!Z�g}�ۙ�EtB~��A�0rlF�$	�l&�5�q�\jA�ֹ��;^�~�9�{��-���zsm��z��u����^��x�ez~a�/��!�a��("�`�ׄ��Ç>x55M���➞noph(�������|�|޶m��Ǳ��U�t,б@�t,���׾�m�j�����wu=��N�P�@70���?�>1=�����L���	����[����P��r�*:z�e�9.2����.[F�b���"Œp ��`�!:|� �8���A��ǠwQ
�ʋ	tXſ9\ʭ�xk�]��e�˝ۚߴGk9H��f&x�#����q��B��󐑧��~ں�T�ȇ�;����:1�l~���8���<k��f5,7�ynFa���\���n9~|�7_Ā�Fwvvr}�2wea�FJu�i���5����j:�ܗ���I�,,�ѣ�X��Z��͸��K����>���΢;d��4Տ�Z��׾��h��:�X�c��:�X�c����^|��/��?���V>��Cܵ����tOO�B��U�z���!��՝�v�I�Nb�U�92D���8�T��Ӭ���+"�˖-���"��"͏�C�2��]�x�t��e�l���L�4�3��/(SS3�����)N��\���!m�ٴ�6�MG?uTO��9l���*ZF�Li@�������t��E�]M�8Nc�#l#l8���~��i8}}��T,~����_�^�����_��V��,,� ���U��� 4guu��.��e����Ao��'Og�徾�����w����7��Z��C�=���\܉�>��vggt,б@�t,`-�K.��T*���+�t���q��8��GG���!�{�}���hϞ=�!2��p���Gi�I'���,Dȑ����z����4+@$V,]:N��L��!~-�)x�)9r��8���~����	 �^Sdւ����:3�	`I2�̀���.=zl���������"x��k���Ip7�!̞�m�r��Vڟ�uu���.��`?�W����A�she7�]��q�С�����NDw�F���G��o;es��s�7���7������=���.�V�n��(�=H�5�MZ�~�\�����Gs�s4;7G�&'��뱐�e�]����52:�,
*��]CCŗ���؉�v���:�X�c��:x�-���ι�����\r��AWػw�[�Dm��8�����]w}�^v��ȣ�p����4�t��t�u��׼�5tםw��ի����c۷ӎǟ��O9�v��E#cc�X#�be/�y�)7���"iBG'�0ow����pV��sx-45=���u��p4x�l��8��ǧ�o��[x�7��F�1P3��y0�,����MͶo�/���E�T�e˗�`� =���T�����jFW�D���d���0">���F#��}� �7�j�^Ԁ��??459���V��a�>�}�Zoi���ņ��;�Оr s�B#�a�W��J����}�����n�JK�.����ۺ�����7�y�y�v,б@�t,б�/�.y��o����7���C�so�0�w�������y�]t�%�Г;��s�9�u�f^����W/��v��I�~ի8Bz�7����}ڸi37�cJ@������lk�$ǔq=��k/��� �W@o{���e�4pw�]�<�ڡj�A_���|M=��� n]� ����jQ�L�/�D�$�D�YxtϽ��+9����n#�!.���M�:>�:�Y��gx�5���^6��]
���o�-�7�<?�xq�[o��w��£�ssK�MP�����	A���ϸ����@����	��"R_��u__���W/��E���������5��e���w����Od��;�X�c��:�X�y��+~�����������W^y�ɬ��c�կ~�~�w~�@�D��J�J]]%V^@��(*�� �*$������G�j�z�z��~G	�X��~��F��6��J�đ�~�8���Ѿ]��J�UT���5������o�����?�
	 � ˠ1@< ��<VhX��J�`���eI� ��l�˿�1AM E���}/�n����TUDo��`�f��z�Y?K�j���YN9������Z���M_��m��9��^{m���[?s|�}33ӿ�Fq'��Tƥf�(�ъ�/z˩[X:x��/,�./��A�D�5��������?��O~�\n���|�X�������Nǵ��Y��c��:�X�c�_X\�ҳ~wpx���7����RB���_�J�����733���l6�tl�47S@����`)2l?|�A����X����^P$h~v�V�]K��܄� �̀)F_7�#�1ww���#�&(�o˒�L��������\
D{ҭ�~�~��G���tȖ9sp��ܘ˟�R�1 .su��͘��j�#� ��ۻ�������G>�a�H4u�6M3��wV��Y� ����3>�)ͺ~����t钛�,Y���o�����ߛ���h�V/�H����I�F#�(Lȵ��1�]�����cG9- /inn�2~�&''������}����_�%�} ��}wp`����w��_�y�s�t,б@�<�8��3~������|�o.��Bu�豸Z�y_�ڭ������RWw72�t޹g�$U~�aZ�|�ؾ�^��8z{�ofY�C��Be��L�z{�h~n����|�#�Bi ��tx�l��"�ۮ��x���B�����(�P3^���۾~;M9�Q_�Mњ髶���@j� ��f��
:�sx�>��������W�����Y�"_����,y�����Ӕje�����)�=@�vhp �S���w��׽��_�y`����>⮿������WU���A���i��г�W�
^x�"N?�tb��;�#>??�r ��"\~�gқ��&ڻoo��_����Ǳ�%_���}��W����گ-MS禛nR���*533�tuu9N�Xu���L#��O�Ɖ��|a��m[,�I���߶��&���Z�Ժ�b1�{�I�V�W}��ժ3���$�T*9�|�I�57�.�Q�8��f� �l6��� �r���D���D��?lA.h���*��
Z:�F5\Q��)���2��1U��ņ��J8�a6�n;v6�L����������������I�5�hNe�9}J����J7u�<���{���6��y?���tV�ɻ4Ǡ��~+�v� ������k�1z�јH�����8'���۳TZH���ڟ��{־��p?�����t�n��Z"�����MOO�����g���^�w�Qq�o���7]N���_l��Ӊ�!����ްasǎ�M7�d���s��W�gj���S���3>�;v<�&��fgl��o��3�km�oέ?��_���t�M �ɽx�>��W\�p�m�����:��X��g����ĥ�^�C��#G&��������~���g>�Y��e/cU��/����X?u�q���op�ђ�KX��?��
�>r�������t-_��x�'k��Xk���ː���*<�����O�'���J Z��a�����~�V��_`�+���{_қ��\�Vpl��Cm�8���� ��K/~�$�G��@n�
:GD�z�J�n�#G��׿~[86:��F�z՛����C�y�8������N-,�Uk�Dk_;�B;���
X"� ������-[���E3�3t��16�� A��\�����Y}�i�х]�����}�ݕ�=��R������C�Ї��� �^s�5��<::�lߞU�穱1Wek%�����y���*�Ӛz�8���@��n��r�v�$MpS*�IWW7t�u3lROW�`���T�V%RJ�<1P��
��@t_6�u�A��j�f�k�z���C��`6�71NC�2��͐�Q�I�(W�^#hdr�\6
r�L�l��q"����3:�b��L6u\G�@g<��~�[�R�������(vc�F�����92I���AS�������0RH�tuw����j�%��=W��ϟ�ku��2(8�z�����So4�B>}C'�"?N%��y��d2*�b�/���7��X!�����2�r��(L�z{���
H�2<?b���Tx��AS�ge���N�֍F#�}?�V"��
yt�I
�B��J�$�i�FhONi�Xk�7����8n��e'MS�����\�Y(7͸���D�4��0
��J\�&�Oy��� [,���^��J)��V�Q�vK� ���7�͸P�QGn�Ď�p�f��l6i4Q.WH���8*�bS�I��^�ѩ��>D�1_�$��^)כ���q�Ui�T�B��n��ƈ����-]�����̶<c,9��\�j7Ց�S�M�ȅ 7~��
%!�㩔��s����K#/B~\���$�x�`�*�B'ՔSrh� 91��u�$r<����x&�lj�HD�x��b�9�G1��D�r�a��e�Y�Z.��2~�fq�4�x�(�x|a�<�G�����2��8��0�>[=��0�Q�����H�4B
�J\��Un����x�^�g=?Ci��b��ԫ���0Iu��|^�bc��Iy�
�X&�~�i:�������|>
�(I�8q]7�=RJaHi3�4�q�8�I.�m�1��u�</�y:D��	��DI��J{��?v]�T'�#�s5��U*m����A*4���O[���p�$q��*G"Q�	"S�����:ѩ	RyG�_yY    IDAT1R���qL�Ps�i���K=�`����T��Џ�J2Ik?�M��|�� ��"l��l�O��Z��eSE|����X�Mgg�i�\�{��XJ6h�,=����������y���,�8�%[�����_t�E���aOo���S��[���m��LLжm�8+�r�
�����yƙ��#�pQ��@?=�k'}�;ߡUkVӉ�i���e��(���Dx� �*\D��С�n �J�c�-�0kpL��!`�`n ��u3v��d����n�� �f��N<״`���em�p��h���P+z�������e�v���@]@qZOw7U��yM�9���SS
�����]����Ë.��je�w�w��G?�����o�������s�s�A�C�������N�֭[ǭ���╯$��R��fff�/^c����l� �7n̝}��4>>^߻�����S�?���[�Թ_�x�r~v��5�L&Ӻ�l��D��l��r�y ��֔Uq��X.m����j���\.��0�fg#���F��]|�X�q�a��@1bΚ'Wh��uY�8Z��j�h���2$פ  �\N�Y_�����wvvF{^FA����G�K��(8��А���c� �I�BŤpt1AZ�D���Z���ˉ�X+������/&&"�k�}B��[�������f��`(p��?F!������rڴ8�`�G�/~#������,lR���$���/�4 %���n~~^�㞛�S�&#���V�� X��86�cBDS�\�`c�؟|�{ �{����wao��|&x�'t������u>�W�8u86�L�&W)]�U)h�v�d����Ts�uh"&1����mp�`\'������a�P,h��;Ʊ�A��1�1�(��I���	���-'ͤ	�&�W��9fi\'�>�3�����m&pI�{�a&_�V�o�(e|
F��$ &
*�X��F
萟�4�}�u'��y��p,D5\קuևN�p��㷉r=7FL�]tH�ٶ�<�0�	�P�+|f��0�1`[&m3/b���O��<'�B����PJ��"/F9�݊�Ɨ�V�q�T� �_���Z���DkTO[Qy�2�1gAMp)Ld�0�����>��+���1�kP�V�k|B��,���Sȵ:)� ;��|�pjI���Y������)��B�)�k�/��8!k�z�BU;�m��|H!E��'G�p>S 0;�M��8~����(�v=�n�WEe����	�P�DǾ�����DgQ?�G��Lv%I{'��A0&��h&�uS�N�&iC5�r�:��䪦Gn��;I�LRUW��<'��V1 y�P���0���i��@��M|�Q�����F#��siVt����رR��ۛ"��� ,«�����T���K/9`L�A�'����_�r�韾D�r�&'��W\A�B��
��Ɨ��đ#�i�&��룹�yھc;7d@���D1sz��-23�7M4Gr1v�ϑ�ё!�A��0�����Y��kR\�v�=���w�N�ٻH�0��v^j��_<���6YG�״�!��Sb
�e�]��ׅ��c<g�o��
P������驩x``��N'��>�Ğ�^���x���o{����<��Z��v�Nܨ7�Z�Ω���q	�$[�T����16������=:1���D�a�Mؿx��1�^������=�:E��r����~%M	�o�$ �]�.'%]��|7����ӛ���.�s��(���cjvf1�Pk�cp䴧�'�Vk>�En:� �Y��a@�S8o����yH�R7[#����A�ׅjN��B�@a1�����10aca�uXb���\c�(�  I= �b��2����3$SG�@
��:q��z��TIl��� n������>����>r�g����Q�i���q. �A"b�Q3 S\�ѣGi�ʕ|. �x@�8R �x pM��j����T�9�罰P���0p<�1��ax� R�;�'�/:���{�X�`W��{�,^�"B�}�5��8�o^��q�����)C� �s�9Z�>h|?�!�n��Q��g������ ֑�-M�����#�+.�2l3�d%ep\X�-%�3�c���up��
�]���[�W1����=���&ZT"���{���7D*��k�fjR�a�l�g��g�r �Rw�Zx��\�_��M�L�y��l�$�ϠOY,9j �r]�qj����{CV  �ύ�h���8:�+��U��&�\� �1΃�S�9Ž�����:�N��-pfEB��u����E!� E<a�u]��u+���'�2S���-x�xqƪR�Y|az�'�)χ���ր���(����4���
qAsN,~�hvg����MA-mPܛ���u�����0o�;>�D��	ǘ���|����1pM���g�JF��i�H�i���XX��H����Q�^E���|>�	�?w�=W��\��<�C�qJ�~r���N�8���")Ju���G�JE)"�C��D�$ҩn(r���T�(�%i������8Z���$qY��٬��l-��r�J%��d2Ŧ�9�_U������ew�u^}��'h�m��C��
"���'m��8L޸d�R=;;��G]{�����#~q�m�1��Z�K_�RZ�d�׽;n�ˀa�`�Y�|9
�鶯�Ɲ��qm��R:����U �\`�5��WC��������`�Q�`
��x��L濖J�)qd�\�b�m9��-_���wP3�����Dy�)f.��(`k��(r�?�v�"#�-�4�t���N���Ut���;�Q������6p��R���P�(�es\�P�˗��4=�"��l��ڿ���U��w7�pyF����C�v���.��:��3���.�s�=�M��{w���ƀ���zsa~!�ROLLx� ������!ꈭ^oh 'Dp\�Q�����I�D̿�A7xfz�#f�yv���!Z�h4�v��M�p#��a��[�Th`p�$&3�#�!n>^�:� �Xx�� Z�Y�!@�  ��7@"?�k������:G��m&o��y#�h�F���@�����+B�����Qg��I����(��<!b;�} 86b�?�M$7��X�(@���x�s�B'dx�: ��a�Z����ʈ΂��4~�- �b�,� v"�D���7��Qk�e��Qk{�X�%v��
:�3Z� �����"���`rCd�͘�t�ᨑ7�3�|\�7QM�"���Y�)���G�6�@ �A��<y��k�aq���d����&Ƴ���\@��=5�Qx[8^&��� M���OaC��#g�1��s;���@���%�3�� ���X|��j�v�bW�[~���CZb�/�0� �p��1>d1n �˜�~⶛jd~$R��$�v>1�d9� m{�0�����Z�3��`��-��B!�?���3
C[�#�A�C��:"�fnr[c��?s/���p=�^!� ����DtΤ�J�����c�b��=���NII$�S��Ea|ǟ�>�XA�}O̀iRr,� ��8&[rη�n�)�vc�\������pk�|x���F&+�`��e�`�x�A�Ü[�Umƥ�Y��Z����3�6s��x�1k�#g�Z�_���e���6���=�S1��ԅR�4�r�US]]]�V�*JAڈC�z�X8�����|N7�D;�Hx�Nk*'��0���zEu�uq'Q��䲹j5��F�V�sٺ��CGU,�&ݦD	�MW9L@�Zk�?��Q�1�U�J3���0H����UiQ������I�D�S.�I&`�T*E�%^&��bɇs�IR?L0���Qty�$��r�
�"8�����􇆆y]��;�eN/��g��Gx��K7���N��c�	��u'����iz�ǏҺu'�S��r
4�����]�H��^�k��ݻok�/c�)��e�켉5�H�Y]]dM��!��%�혊�2����:��4�[�1�]�Z����Et�8c�4_��$�'�8ñ�S4��N�y`��6�Hg�c�9p`?gI��������n�˥�����֭=��/���6Po�ᓽ�Jp�\��j�ޥc�!%��y���*���)���e�_N?��}��餓O��[Oc0e#�J  �u�Vo�~&^d�ZC��J�0���p� �k�׌)��8�� ਏD������J��f`fE>���(�@�pG-�e�gB�&����)]���	nnn6P<DXP�%�� =bDD�9������T<���"��Q���QE�Ϥ6L*Z"yv�jE���_|�S���We� 6�"��#��1��F|Z�g���<pD4��"�!�G�# E8w�i�#׆�`�/S�Ώ�q5�R��Ga��op�v&�ց���q]x���A�rL ؖcpKö�R؜��&����^��/Q�Z��)S�	 @����G���Y���"`�Hv=�l�S@��l���:;�n�k���׀q
�ՠ=ʅs���	�b�c�&�3�]a�f�'��Ǒ���s�#���#�^���xA �R���3#Nn&Y���$�+��+�hk��b"�ߓ}��D([��ǒ�n߷L��o~�G *�,ƥ<O�D�1��x-��a8��z�ڑo*2�g�����d�-O~'`��ff��xk%��~�G�ni�H[�O��=m�^��aGc>��yv��4��g��e2|���sC	2�R��,��xN�csD��5)�Q.,��L��`˽�h�DO��Y0QM��V�S�~8��~qdUz��Ⱦ|�s�(m�z��L�9�Uh#��k �F��g�eC���K���xʹ	��Q`�/F��$�/�L�I�fƺ�k��u9Z���PC�!dXN
Ͻu� ��,�0;�1��e'������p��j:k�r���l?M������#�)i�-7�'&5P������`��u`_x�ڝ5�Q �{�4�a�5�y�L6C
���?��b͓��������3����L�4��$MsP*�g�F"����M[�����]�����]�d	ϝ���?Ӧ��	��U�V�w�^�^�@�����N?��.�	E�������"e`���S{����e�\�"l[�2�M�Lp�k�8��F���{�����4q��薵�X��v�3��k���$�]��81&�������^.t[�j�����,نc��.�,�����Sp���qw��ozݶm��Ǽ`��Fih?C�y��f>177�J�qLf���GyD��p�)���3����ן1�ݴq�/�8� 6��̴j6���hÄ�h4b��x�\nh6�
A.�Eڇ9���3��J���L� 8�W� %ȼK���r��O���D�o��5x�.G�lAJ��	���nY�\��h�/��-�R��SƜ�C�� I~Rm:���^���P�S�QD+ ��"� E� I�pUmO��x��p����
�pē&Hh�4��V�v������x-�@"�8WL�f�4(��JTGƎ'-��0>�lp�+�PNÀ�������i����j�ٴbl=Ԟ�22؏���/�͢�ץ�-`�� �x��8�k�3�k�M�{��X�5cc�A��r4�'<<lP�Hg|ԏ�D�'m�^`�=�����0�#v�')V�vP�}D(DBj� ̀���<F��o��D�e�2�C�Q0���#��ޤ�o���4��b�t9���sԓ��R{�K;9�͸�n�QW.�8��Y
�r�s ��A���Y�J��3<l��4R� ^ĕ����|��Q�W8>���S#mڈ;-[�=���ϗBy����&Y~&��R%r�V�OT�!���3;�XF�8���iv��rx���07ro�8aG�5� 6D,�c�T3���T+�l��P<��|��&cc����aZ�(�1S�%������1��v�q&Y��SC�O�3�!i�g��e� �<W�a���# ��2ob54* p��tXz�����`=0��3�U�'��uq��
�ǜ��sЈ�
�\��533e��c�|��|�Fb����	����5%v�6��ƸGƖ�a��8(l� �KH�	�9W����5܀��8ˆ��q�p��Pr�ɼg��mI�~�^3�Z|�e���d�l�2g�,w�t3N��`����!T���1@������	�q1����"������Pxbjʇ����XX.w�?K��w��UA��T�Hm�X�=�0w��#M���M߻�ڴi� ���:������]���@6��D�D���=��ъ��Z������)�hkO|�������r�w``������&�Ʈ�n���Z(��2c�k�:H�c��~�L� 6lhQ&�?��zz�[����P#�,	Е����\6o��������,��Ol۶�S�zA /��O-�����'�f^�*Յ" ��^ea>��8�w���-[�z�7m�`����zU.�tOO�BԴ��wZ!b�IX��� ��ˍ�dc��M�� ��*�yR�d�������HE!O��� a��1�0�W ��m���Z��6(aDCp�"�� P �.<���H��2�0�u�5&_��?�\�VL&�CHD�D7[��2�.G���v��#E(_�Vc/U"	�� E	D\m�!��,�uM�!�"O�(�G��ky�dBC-��/�t~-��+[p�#�-�2��H.���-;��5��O���"	���`��`
[��L4 @�/�v�04���"���f���� ��-)H���,� Y�`#�_*q��D��Z�Ţ����ȍ \�`���ļ]K��}�"�i�'��� r�X�%�K�>gM�T :"�<����8yѱEY�d|�u�)���:~�J�b���f��@���������0-N������G 	�*�-ֹ�g����m�D��B���8���م�ŒC�y�yq�P�}��m<C�{0��K\djsݚwL���T(T��[,�g�����)<3Zl�[�qq.����#����0N�M��{�t)��g����1C��g6�e�)�1��8Ѽ�[�,�n�<�� �/��gF��b"��$��(�E-@�g�(�1(�4.��费>����������ɺcǵ\/� Aqh��Fˉ�G{��y���2�8�:V�Q�)x�H����1�����4�uDB8�L��0u�=Cd�D�����1=5ej&x�4��m��α�� ��
��}~�(�����^�]��i{�#�E=��F+��G�:��f�5<��Χ��ź����(���� cj||;�w<��0(�}���� �������h�L/
%��m=u+8x��ȶ�z*�������AI��dp�h�;�����r�:^���(q��ӷ�����l�Moo?}�#JP)��mE�-M��mm#T��.��-�+�
۞�
�$�O�[�����vev�<����K:15E�J2���e�=�z�%�.w߲m�6+���K~^� ������̆���7Q��(�ʾ���4�''������s=�."� ���l�������
*<�x� �	
�.Q^�Zٺ}1���bB�F>Q��h���T�D!�1 i��ǖ�?&�V��V��,�g�|Z�"��V�E�T��4�]89�b�D���k��X� f
f��*@�6���n�C�*�:�#6f�d���V�(Y"�]���t�Pc����Ij�������MմQw�M��ߘ4%2�E�B<S3��V���U,J� (�s��5`R����H	v�	q?$j�c�|�V����ʌ�;�K�'������s��7&L�����B������VH%=�O"r1�{�N�����Xf�    IDATB,��(>�B�g�h�g@�����.(����Lt�<�o{om�u�w�sΝ�\�j��Je��ɒ,��ellc���lpҋ��:��������0���Â`��4s�n�-![�JCI5��7�������w%�4�ut$�wת���w�����9�����!Z�\��%��,�ƚ]��_ǵu�ְ��3��b��l�!>�}��:*�x����v�k�8=m���?�u%�z�_�gL���ř��ƚ����B�(ˆ�AV�Xh��x�htp��[�2�ɭ[��UH��b4n���݅r��2��V�g��r�B�u\�DQ��[�J�xǄ�4-2��&�v��VKs���wu�
�*�hz_�ww��(�3q�+ޗ���~]�L^b��Rӊ�tm�@��/��/�X}��_�C1���9]#~ݖ�;�q]:c����s�����6-�qAnBRYl���ן8$�^seu��]����\�(�ğWj�牸���\���r1w7�=�Ŭ DO����O����Ҹ��N�t|��GA�>n�g5V�G,vEF�Q|��ƍ;xq->W�8��\z����wB&��̜�g�1���I�'��>�P�U���;\q+����~��*��:b�J�˦1�9xi)�|����㧭�Þ�{�̸q�}����y�P�%n�B";|vl�n�i�{�X���J4}�+����K.�������̣�M����Y�#Wm3P�9Pׂ��vm�ύ(95_�<W�Ţ�m��?������>S�]��)���4�}h��Arr'����c�l�Q,S�������c�?���֞|z�<����"��Mo��ܵkwPZ2�{H������ڵs��+.�^y���s��;�y΋�yx�2�[
��W��=}v��?w�uE�_"q�]8w�%�p���̊���J����T�&W0өS�L�3~Sh�d�TJ)��#˃6M�fEP`8�V��bj(P�IG��C/�rsj~Y�ˇ�����rŜ6�h�Y	R�0=Z�y5�Oi��#զ�D��}�.r��۴v�:N	f����(��V�.d�y��sT/#3��XNPv(���P����ɧe�ln�k��E��h6fu�*=V,s�IȬ楕5�dŭ���]��x���A9�r�1����������[\���[�YTu<.�􀈮)]˧�mk�^�	��B��z�^�~��9L4+\|`YPX9��"I)��m�8�]�?D��Bښ�-���~��J��/
�!��8[�8�U�o��[��<��-h�a][|K��J��͢�nA��syϏS�x]uYr|1�~u���a:-��D���/�������E¢̞1�ϺHt�eT1�b�����K���/0���,���R��a�VH]G���HG1눻�L��޾O��^��}���P��]'���-s�:���<������%���� ����2��[\ ��Pב_#Q��	���[���5�1���-�����[p�~�.����N4x
9�>���B���7��s������]�;W��4g��S�E�ZL��7(,��(Ztyl�_�f�/.�bI����#=��nH\tLΕ�ciTs����vw���W1S����;�:�F�v�Q�<�s��S?m��<ϡ*�mGf��ֵ�{A�V�	gϝ���'xb o<n�����PZ��1�4Nhg��p�j�Z���yRsd������g��}�tұ��&$eT��-���W������V�l��=��˯0�{��m�S-�&C�������y��A_��<����n�)?~�D�b�$�/��rOYh!)��m������4��ʠ���y��m�z�w�����0ޙ�����l�����y�tD�9�M�o���w���/��̀�h����-����ѣ�ʩŃ��׿���W����,��e�3��{�}�鲱�iX�2�?z���t{��w�y�_=�\�|�W�����_���ܹ'o_]]}O�߿!I��|�w��ևgΜn��1Bzue%��-Z� ׄ*����:�)��y�t-��DdLe-�0��y(ߪ_(�W9I�wܺ�?'���V��V$JH�ߛ���u��ض�����$z��r_4��օc��~�Y@]���r6�SZo4Q�z���*�ӑX�m��d�*�*��L�T�;�(ʭd�J�����+A���z��>�>yF�.?�-�LX�[��>��K����e�s�GD?�迬IK�ī^�O���=�5�㼸m���'M���)Mރ*KȆ�\r�%��A���8y���*�r��I;V�ww�q*��ϭ�jC���C�����u-�t���-��z��t�J}��c�����H��E|00��]w�e�P�G�����o���ͳ-G�^ѻ%�-�n�T?e��XYO��˭7�a�<wC$�~��ȥˏ>#��ŋKVvS�0	�����t���N���D��5�Ā����lg��tK�k"ָ�z9w�\�=Pu#qZ��,״G-��,iхE���?l�j�]Y[�q�������[e�"��P�ndSq�}���1�{~�1�{�_�.$}^���fv#&"� )�?.�ݲ�g
���c3��VMw)����j{��8WO���0�Ϸ��Z\f�`tK�ϑjӯcbޯ�����/'���5�~���&�]!�Ϫ/����ͤ��B?,�]��n*�%I�q�DڄU>�=,}xK7;�-e��s�廇�bj"&#���e,c�Tt�YW-0ls��2շTBV�w��k�\�.L�j��w��5^22�F�M�E4 h<d4�	07E���-p��Ȼ{r��i�F/�ɬ]�nx������lP��_��_�ڟs���oxc8�ȱ��s����%��n�a�,���9�H��W�'��_~��$���+C�XD�x�8ȝi��=vL!���^e���?;V/�]�$�}2�ٝ�
{^[\�(��6�{���?��ٳ�L���-P
�I�.|��3�Cl�nV�P���8��-���n��3da���f����h�"�gΜ�D�gϮ�������F��?�S?��χ�}�6^�[N��'?�sמz������H��������I���0I���5-�Dɱ���/>\{8�.8��{7��5a���a�]q[����Ed���ߊ5���mY&�m'�m�̳��k�����!l+J�\ʠY^<�I}LB�D���Y�K_M�ԕ��v�[	b�-}��X\�U�_՟�]��ͭ�:Y}'�#��[���J�z����D4�O�V���$��#p�d���rks2l��E�ڗ���Jɧ}�1�zɟ�3]hB��dM�-��Z�����6q��r�>��ֶĨ&p�����+M֞{W��{��J�K J(>|�xk��
\Ǡ�H�Q��OA=����A�M����ک����];�,ؤ/��������Շ��رc��k����74����W_m����u-������>�*�z@�I"Y�ݷp��-V�Pb���������ĉ��z���UjG�� �-}��-����xL��U�S��D����4�%@�b�_���zU �c�=n�-�g,ǭ�D����8�=�����gu�zi,_s�k�g?��h�EƔ�w�6�g3�yh��3$f���x�G��9x������*�#x�q��е5kSׅ��z�)w��O�K��S���+���Y�kUף[������a��/��@�"��ח���+wAr�>+����9�~�ˈ��8�A�,�b�J�T��9_$�x��r˦��ntA�F�p��Q�Zs�)���lkm�v�&��n������v�h���d�,�\�eY�\�Zƞ�R�����wOI-�1?�^&fʬ.�'^ގ���y��l�Me%�������J�/
�w�ww�p��s�,��h��f�w-���\F�De�Q���������3%��+n�ǌ,�J2�R`�L��l(c!�~���E}|h�V�ŏ�TϬ����D��?C< ��[t݈s>�ls܉rk�� LҢAh[([<I���ؖ�Wm���s�ȑ+�G>�1[�J��������ݻ$�����P����s� K{���"Ӝ�*k�t꙯y���C=������4�[Y���C��tW�,Gץ�UG���E��i	N�'��>�q�6!!<�򅖿�\��'??@<���w��Y܁���rUd�ܹ��H�c�V~�QΝ?o��Z��ۖ9ix�K�_��oz��]�z��_J�g��s��	^��`���w����{�ћ���5!)�O�9=����ȟz�D�܄�V3_]Yk�"w˜Z�����s����mq[سw�=0v��m=D�ä_���utA��~��٘Gtl+�t���0��ߴ���EAY�l<BU�	ãFu�e����)�ᴽ�U����շ4�F�mD�4������?o�kb���Z��ru�Ь[�����/��>K���IQ�cYQ*�L��Ԕ	d��S0�Y�إ m���+z�[@[�e�B�2�`��'M�B��C��A��i��,�:w	<Mb�c��$:�Fc���$��a�F�-k����\L<�T������Xu7�Ճ��-gsm�F���Rol�*}�t.zp��ڲ���6ӹ�U_��ﾵ���B�>�1����B���ks�(���{'��t,v}��r=���d�}I�~���]�-��&tg���-Ϻ�}�X�j�}=Pe�ѢD����>��1���g�9eX)-�vߔ���`Ό����o�~Կ�[�����~���c��Ų�G�)�Zch����:�.��~�]/>��^׻�CYc|��=	C-F��,��eT?-�vi�w�d�/�Bom���*5-]���ţ����t?s�kQ��_w��_k����_OT���Vh�ъ]����]�.-~n�0��2�_��_Ǥy���S�Oٱk����RbR�Ʈ�=#�"�s�J�y�ͫ�[g���X������b�|�����x���Q��8u����xf�4�,�ʲ����,c������k���8Ǩe�m��e��vsA-~��t��Q^_:�]�:O��L��j'Kb.�~*;O�����y4BlY�yQ��>6�-�_Z�=@��CY
ܷT"L�������߹��]
�O��_��an��E�풕eԶ��w�,[GL%g���4`z�]����oy��m?򑏆V�T9�{���������l.���v�cc(n*;�����8h�Sc1��={���n������<��I4�)h9�Ceឿ�;,�φ�ϪX�eA��J6u���+�r�x���䘃~hk���o�x��&x'-�.v��f>�#���������ʵ�N���fS~�������y�a��WVqe�Ю�ⱔ��'Ӽ��d�׾�+��[n��g���o�����u�EQ$?��?����tsw���N�h>�/[^^V-k�:4N�<m��*��A�o߾T�.�h5h6�ۖ~Zf3��Z}�0�OexX�[ܾ��)����+�X�ȷl��oc�\�2?;M��ߖ,��o2P̬����m���m:^��%�c4!�L���3�U�y���/.E���M�p�ҍ�	��#�tg�����JKC�V�M�zx�LP�Rtt�ɳ�^HL��w��Y���=$��rV�D��G�}�p�t~�6��N��[=�f�MaY%�eD?5���W�b���hb� ��b�Wgm���r+�=��C��=mY<�\�>^�iV���1S߲@�
]�v����tO!�~�Y����b.��#�V6q�?�'V�[Y��>�#����,	:F�'4�x5=O��[�n��1�!/�ǭg�[�����-�-s|z�.���\zJ�L���U�������l���w����d��>���2�w�P�:o/� ������l��(la��Ec��I�.M�:o-�t�8{}F��u�Jz_�k��0;���zW�bm�O��$77���5BN�ܭJ�V�������HzO�D����t�� � >�7]�z�o��ѱ���ެ,w��ir�����J���u�רm�x�0W�zk��9T;z-.n7��}kS���:�/���b,u��()c���ÕZ�w/?����<�?�,���{n,��4��v��RV�3~kn�sG}�p���v1�~-��J���w���_ϲ���]e>�HǦs�N���̌��Ug0P�$���W�,,鿮)7.�*�1Y�Y�g��OB�}��[�=�(Q��P�����:��������zF%]�����rn;�V�3�����������t|���|r�t��n�U�ٹ��P����Y[�Yi��9��O�3KZ���2�>�S��{��{�/��/�˚+b�c��M��o����S���ǎ=jnO�8a.�_w�vm�ܙ�<(;pLK�3?��q��w�������J)X���\�]��?;7?�����'�`SY��m��o�wLp+��|�uW��ƶ/&v�}w���V�=�o���H�շ�j�
��~�~(��_����>��%v�X���m�w���ݘ"�>��c�#G�h�|�+�����>����c�R���Zx�� ?��C����{�-/�\�5�W�{��z���|T̮�������R��������0�RS�&���U�}�4��u��2_�X�(�[Q��)�*�`](^>�� �"�*5I�e�Ge�������v��*>�!��h�T=YK��W)���IB���Mě�d 0�[�q��+E��]�eZqp!f[��V�nz�cY|9������ĩJx��}�qUQ�Zݕ�n���kR�O{0�����������z."eM�skD���#�݇N�:���\}O���w�"L�S�׶m�zl�Q��]�W?��ǥv$�\���19}����Xsk�D�Y��̬�����=h˅��)����o.Z4��X�����#e$�]+ed��׮����������MO��aV��,��6��d]�z�Sx��q�_ҷ�}�-cb�������������x?DN޿[�l��}��g��v~�]�:�()=����`�N�[�c��6����u�t�Y}�m��,8�O�m��_�>���/�|�s۾m�xLtf�*ŋ3�w=����פ/6&���ʷ�}��"B��x�r�"��5�1�5�������{T}�nZ�E���ݶ��1K�����H,v���v}1��k����Ԏ׽��"��*2�Y�4O���c��zdA�]9�ta,k��]q��|>r�]۶p*s��X���L1�9[�-г&����Js�Q,���E�Q�y���r'Fj+Ι�O�ˊt1B_���ǭ�z��e���ЖAȪX%��A��h�p��]v�+IgJ�[�p���p�ˌ���UHA߿�Х6��H�+͛�o�>;��ra��[����>gצx��L��o���Í~���1��M;���E������X��ҁ�zq�c-�*^�by��U�+�#ǂM+�}����oyk���Q ۹kwx�{�>��o�Rw��Kh+�	^ϝ�u�b8�WX��Rp���*��`8��J�R�=���&S��X)���=�n	����޳�Q-�6���z�ŹK��qn�"V9q�=5;��z�d8s��Y����f��I�k�T�3�0����[�Q���������}��i��M�d����3���1���:v�t]�-�ma><z���;�x�/\v����]�x������>������D�����|���y>ؚ$�ֵ��-�V{g��q��j_s�̙}�Q>��f�$�|Q�������j_��&�D�~BJ���U��:[�M1�0�c�v<���fi�Jː�f�e@�D���z�J�p6n�mr�"&Ib�T�S��`�2��o��o���I[	ŵ�V���^�%<��^>==ee;� ��2&~�1��8!7-3��Le�¦�$Z�R�����=`���|�����ҫ��*����"l0����.�Ԧ/ZJ_QY���D�T�u�\ ��ܢ��Ē�������N�*׹�N?]�4������_�
��Rȥ%`�I�
@��׫q�7���?X9j%��5W�+i���I��ܚ�|;�?kQ�V.W�TM-V>ڜ��"fr�N�?��2�22t�q���%��JZ�<��U��7`    IDATTn���Ϯ�mj�Yב/�4��t����
�o��W����%|�`�����-�.8M$�/Ll�\���LG߲T	m���Բ�j��s��Z+�Q
G_x�;	{��uح�~-y�=-���;*x����˒�c�M�/����r��Z�!�uݮ�B;W^f���Js��LT��r��S�^�g�p�W���'��Ɉ�v�"��>-�yOx��q����[��=U�,}V��JQ@NZ��Zf��M�g��-v����8~�E�Ħ���� ������[s�[�\H{NaϦ1�H��c�JVef��R��4s_���](c;���}>>1��3S��+Ziշ�b�.In�йĒ�Q��q_q�\�T��*�s����x��C�?_�y�js��w�*�[n��3���g_�ճ��Z��.���~�2팜8q���(F�=�Y���xl1�h���_��E�D�}{�~�z�)5�D�������jO�%1�]I�᧟>m�
e�P���Xڴ�R����<^�ʫ�G?�1����C�,����D�3NCtG��TL���������v��@m��{���u�]oB^�x�F���ʬ�ʼ��6Y��ϚK��OYNc��ʲ-���R |S�zLA:Sڦ���.��������X [\�yp�3Ӓ��}R���c�.�ߋ��;v�P�"+r�{p~~���dY6����R�v_�Cs�v%4����͵�Si��m����?���ɽ�����JR��n���0K�E�|�C�����g�N���v�V���ۣf��o%���l,v{����b�_3^��vw�����P�TuMUsL�Z�r�h�[��r�V�+U���*=����l�҅�A2�k�U="�Ys���A%s�o6���v��EI�{�)�`�(t�0J�T�]G���<��N��rJ����~���ٙ�p��G��pmu�7;7�k�Z�S����z�z��F���;�3K����W�͢9hLgâP��~6B��!�.�%�(���Mͦ]�tVdYZ���os�Y�=�7���!��hk�Z��Z�D?C����T���d��L6���,�K}���$n�m�E�^S��Z�_;6��+.^�1@���r7MG�Q��3i�\���v�Y�	!\ظ�m�/q���e�;�N:��H�iVdô�]+���x���'�����NTF9曵ҟ�\�������e�$mE�ɽ/I�F�!A;lE�%�Dk�Qk�'ma�T.�)��B2�b*a:	IgT�Z�4�������C3Q)�����*�1����ǅJ(ҤH�������E:�U9���H�z��f:*���]�!��D�I��yG��H��DU�:���*��Q��jTѐ	%^�#+u�hC�CR��onnvf��J~�o�[k%�Wyo��%DTe�R絚��?̛�F*�[�4�����t��d���_[���1m���T�d�XZ^����Q�������^�A����/ŢU���8s�-�T��,`���x�w$�=��]E<��d���[��n#z/�����ʨ�q�R{�W9>6/a=�F�B�|����YbU��h�����Z��E�[�Է/R|����g��"�틴r!���H� /���
�%t�kf�S��Ō�a�(S������S�r�
@��/�|QMT�ڂ�$��(��՘��|2�2���1��lĩ�]��2��U� ��g�Jx㦅l���L�4'n�3�ڥ(w�<���[\	k����)$H�}��+�+r��w#��}^�O�$f�P���0a�;T�R{��X�/w��r�K��K������I�ƝΘ�ͅ�D��(�+�/|�N���bi�o���[_p��?�Z�-���k��淄}�C�{���G~4|�_~��r?�9ou�ˊ���<ށPW}��w�ɧ�UW�+�&�o���4כ�W1�����r�kn1��0�w�L�>��C���,#����z�^��\f]g�[\�)fE��&��j��:�(x�i�k�4h�������'�?)���S���U��V����t�33�U���}�7!o{�m��ɓ6�g�>m.�^_s����W_���#������A|!ޏ����g�2�E/ˏ=�Qb~��wz&��;��~=z�ɽ��29q�D�w��bω㏝ܻ���x��<�m[����,,,$3�����l��a}}6�gݹ�͛�p1mw;��^�gA�f;Z)��Zì(�Z04�Qa���ۑ!�F���lT���QZ�2���,ϳ�ʾi����?��,I�N��I�I���`��nt{��Զ�,l��}7K$��bX$�0
i�$Y�5�Ծ���wҐ֗�i�e�D��̋Q#M2��V��h8H��<i��m���n��4EF��K�d�b�z�Pw&E2i>e���1�HeW�[���lŔy�3��|���X�!�Z���&�^o����N��.B��w{Y�lHh%덙X�:�LO�.\�E"J��4Z�d4� ��{�-[��p(�?HF&�m����,���2X�!���E�,�ZtiG��!����p*
��l�3*
mq����Fh�[���t�h�������ŋ:[�Xv�Xj��D��d���G�53-r:�{f�-w�L��~�h�t�ϺQ�����/�Q[��KHsq*��t�jӫ=����dnn>/���̒�U������S��-��/��|�-Զ��<���|�`�e�RX�]��[V(�z}��R�iG��ve��B�!6�ev�}.�eE�^�LX����"�\t���--����:K��3K��<������3q7/�|XI�T"5����u^�.ow��~b�����*�)�YY�c��8M��l���]8	0����|Q�EF�1�).'��o�����w��ѱ���+���nw�b�\4���Y�]f��T��/���B���}�Yxc�t��{�'��O}<,��ąg�I�!Z~�2-f�3e�u�F�����*\��d��7����d����e�XU:���I���?l�2>�=�}+G�{Z���G/���KOܭgѵc�)���~����z6�g?l����G�ѳ_����y�������r���j�r˚����ͥ���B�$�����w������G��ӧ��33z���ַ����v�{������y��x�[x����J@���>u{*!=y {���O�<��b)��o�������W�������g��$�7_SS���D�~v�SI��Nd����嶗4��DBϿ���As�w�~S���%��	�ì1j$��K�a��v�pJ�R�Qxˏ M��m��Qn�)L4�R�i���6�JJK3���a���(��`;4څ�Ң�F��I�&�`�Hv�T��|=M^�I^���F�ݖ�F�r��e͞�Di��eIQ��F�H��aV$i֐?��xQH|g�^��j�[�Ѱ����I��y��,It���&m=o��A�!SY��`�i{O"��ng�~���(&��N�Lq�
�]���	]�l��eh�A�tY�A?&����Z�WC������V���Q�{�Vk+��?�ti�|8F���r��q>k)�C"Z�����+++���֬��ڜ��MW�Wr	�&h�|ii����&Syي���\�Vo���P���2L@��g���F�,��@cZ�����m����t&"Ʈ3��	��kA�
$m7lZ�7���X���GAJr����&�jv�-�L^�e����n��y�]�������n���De0�������ܜ��ښY'�Bx����ŃvBe��L�)�9%V� �b����D�V���������K�zr]+V�bM��%#���mneNbY�u�X��b��X-S�(�ۑg�e���윶m���7������-($���{�7������D�ЅeB�G1�R���׭p��m�f.b��#�̟��'��+�:j�_���C1�����^�A���p�����}��,��g��M�T{�V�����v)��d#�A�ԯ�F+�&�g<���q��������}�ex�s�r4��ۭ�hϞ=���Р���/��Ū{�ϟ�%����o
������	;2]��w�z�u�{�����o��o9��~A�>�0i
/f�z�m���=��{ｉ��x.�5�p�	����h�>>��_J\�KlOMM%SS��qv��DB[�~�%�h����������]3L���R6��|C]�e��Q�XR�����,�����2c��~+�VZ��YMi(9g$1��Y?�5�ͩV�8BY�sY�cE�tFi���F��9Z��@���N�Ք!\�7d5MBtm�ﷳ,I�a��2�����3�)Kvik4�Gj<iHi#+�Q��p%��6��U�\"4E�oL#�jn4̟<kFf�`�W���oj)�M �#��l���M�h�-�!���Ĳ���#%]n4ZM���5[9�#�Czmu��$>��/qZ�L��F��^��W,��&(�b86ܧ������eY�Z���ж��q����%��2P
��>��J�
6�3��,����Se��q�]�$
c��,�+�N/�^�		�I7���S��A��A�SFf�{'O��u��� �M�"���I�k�ko�+wԎ��]�E�d>	%�w��ږ��9գXnM�q���b�2��Rc�ٴ����Y[hH�*+���'X�Q���Y���K�:4X[Z��=�~̖��B,�b��2���.3T�[���K�T�1Ӊ^^���sS�+�Cش.�VQ��y;�Yrԯ~���·}�Ï�؏[�	��w�w�O~����>:��g�ڷt���6X �,�s���'�G^qUx�G��W_c�ִ����W����+`ӊN(Vd���ea.�>u2��;?�� ���Z��8F2g��C���[�&���?�n�d����?�X=�_��"x�w⽤��fc�m۶�.�]�w�~i�ݻ��c玖,�1�b���T�~-d}_[]��[ػ{����u_�����}qϳ���"�4|qrK(��	)�[��LN���znn.�p��ff&Y^^���ED"��^O��e�Y"{�7�(�,�E�P�z�DZGb�ݞ�PK6�ҫ�\cؐ��|*�a�)����5���a��I�2њv�4���$n˟!M$^����iV�O���L�vai@���I2�Y<.=��,��D+w1,�"-����FSA��6����E֐WI�$�|F�Q�h��� �L�O���?=J�$#�:OFr�)�&Fy���F��,�xC=�KE��Fy��;-�6�C�Hd4O%�ͣ]���TO.��6
wh�xW�g��N�L��9�m��Zn�V;�wM�6��^U4�?׬�E!��R[��+K~�~G�o6��jhA�m�~LAְ �F�w{=�<�z�*��,m��ޏA}QM�W��/��"._Om�JJ��Z�P��xͩ�k�K�xK���#��U������1wo3*�y�cY�c ��P
U/�`ŌJ��R�����=~&0G�qN^sk1��\
T<����`bq����������yY���AVͅ�9�ұ� �����[Au�O},u\����ĜҪv��m��B��ԗ�M+�Q�����L�hbw���L�h�W[1�_L��W�Vۮ	D��=��7���_��ό�`|�?���+��+�yے��S�fyy��S)O�*�������^z�p���a���K/��W��e��
��Y�𷴆�����fg���b�rլ�e�������Z^]1V���K��⢴d����v����=iݵk~�b��5�}f�e�9��i(@[����-[t����ez����[�ϟO=�����ss�z0ݹsWسw��{o�{��t�M�Ợ��"�4@�� `��o^_�r�� ���cǽɃFWY�gf.$�����YI��Q:̥��F���J��n"a.WQY���F����y�dyޒC�D{c4��4key!���Y֐ی�HՎ���yt�ɂ���3-d��"���h�����9��N���.Ƚ�(�NQm	a�3Yċ����V�6�E1jgY#S�Y#k���Ei-�YCޝqA1*F΍"	�"�a��n��._�X������E����n4tN�"�(�߬,�E���F.%�C��E_�I�GA���-�Y��g4*�L*!�6<�hH,G?v3s)��m
�Y.i��Ǣ�%����3k����L:?��JL�}1P�yL�!Dw���K��*�y�]���mk�,:F}ʟY/	fw���}��&�=��D�e�?O��J@�ݚ���,-�(������ܪM��ĸ��������g�tt,�빞/\��>��qc���yc���,����Y��O���`;	Z�^HT�8y�����2!��X��Ñ����F+8x0�Y3\q�	^�:"���t�`P��O<Z�,,]���U��ҫc���U,5F�ې�����I���/�R����Ltm�T�.zM�>+z�����Ȧ0Vi�4���T�;vl...��~?]���6����v-e�������/y��ʵS�{da~��w���ۺ�����߁�}!�@ /m�sp뭷�>�`�u��dv�T���;����\�0���C�-���ES�M٪��Q����������Nw:�N�f�kk+E����F�ΨH�`4T�4[�a�ʲ��e�N������ز|�!i'IҒp�F�BgMY��C�@˙W��a���(�I�����N��6_k}R��{U�L�6���~�f�E_[����huZ�zɵF��̈�V�/��F���ʉ*���ʤ��%��\Z䴚��F���7)����c��C�����;��\37���͚܌n'�!A���e6s�T���(�t�0��h%DJm1��MJ��6�r�_;
��<��.�������]H�>s�����p�}X壿��o��oYnc��J�+��'O��z ;vl7Qy����کhay|�*��Z�W	�+��*�˜�7�� �"?�D�hm� ;73mVj�%7/�|(�E��7f�.˖�b-k��T%�_�w�]e�(+�>C�*���}.�;Yh�fw�����O�puu%]__;s��e�^z�%�>==�SSS���(��Ԃ��E0  @��"0�2dM�u_����ѣG�S�N%r�{r�ېķ��h���5�66�(E�OYȓv�K�B��4Y���a�-���[BG�|a4�
�Y���e����9�*_���&ic�����z�n5���.Q�1�%�+Ko����7�l�|aG�F鋮L2J{���l�j���Q>ZN��B��<�&�p��G������������;[��u_}�QГ ����g?k����[͂}��-��|�e�ܾm����b
1�?���v�5W)�:�3V|�K)Hqx&�hZ��?y��p��y�V�ܻ�k���EA�Y�cA������T��?���T�Ĭ��hi�15��<���Yܦ/x�rb)�
�0�g_���F���K��^wM#I�����+�\�o��g���w���u-?�� x�O��@ ��s���ߞnݺ5ݻ�Br����R@ʃ��;��h�,e��ߞ��yb�ư�]����������O>�R��9|�p���YY���˂`E,�"M�^�CE���!�l�p߶}G���=�|�[���/�ܻ������=���',�,/��ki�$h�2��r%��,�^@GbYrUA�n�5_��(l߶#|�S�����%
�ͬqh<cų2�����<Gt��Y;�y��;�<�///M�޵{Y[?����_�����_�� ���8*  @ ��������{���n��Щӧ�%ac}��w�ގ|vϝ?�n�m�kz����S��b~c�;���۶{b���;w����[P����Z@J��������}����\�"�NO�v��D�W�p[���W�KKLO&嘮O%{�����%�'K[��]׳��@:�&}}�~���.�=S�|����p���e��=�u^��[���~��i���܋������   �$	��������_�8r����_��U�ۻg�e8}���H�_	�X0�JG&_��S�l����հeqф�`X�F��4�ڳ��Y\-G��y���~��)�E�J�zF�f�ҠT~�[g��*�    IDATj��dM�o����\*���������p��3e��{.nc��zvj�I���p�`�W�a~a�iQ�n����?�����w���/�ہ��   @��H������W]��z�C׭����ΝS�B� �VW��U1�H���U��zؽg���]^]5�l	������7�(!W�Ç���W�]��Z^�R����φ�U��lԡ�̻R�Y�X����{�*KJ��Є�$x�_��J%������r��!V'tW��Z��gա��i�V_/PQ�1K���U����|zz:�ۍյ���}�g?�����Cޗ���9A �  �$������o���o����OR�������ť�&t���Ξ=g��JC�������׭8�\c��-[�����0=�<�i��W����L +�Ī���*A���_>fg�Cwc�,m�f��Byn�+K��TS���&d��bK</n�~��;�;.�٫�X��ڜ�/��O�ޤ�߽�]l#�B"*��\�y�7ff���­��z�[���?��[��'_�./�Q�  @ ���n}�?�����oݺ�Q����|J��;�7..-����}��s�,{�
+(���ʊ��X��gf�ov}m�R��:��ewP��ѫ���7}N>���h�Vda-����ga떅���b�˗W�T��$xU2\i┗Y�n�Πlk��EB�_+7=ZŷO�w컱����1K�_�^g� JK�hq�J3��g� �o�2�ڠ��,���)Z�:�N������}�9������xѽ�/�!�  @ x!|��o��[o}��R��;u꤉ə�١�J��W��ٳVnqq�	_���+a����l8�B���&�UiM��
�������*�m~�f5�-`M���O�$�ܱ]%��w�I+c83�kn-C����"�ʠ\�r��O�U�)����󰺺fyx%�%f�Y��[>�`gkW~�zy%>�_���w����V��f�|�����s�������������_�q�R�@�~)��  @ /yoy�W|�[������]�p�� �����K�_�Ғ�W��KKK��V�rO�~ڄ���\.�;��}{������lu���j�ʯz]Pel�hdV�ق�Ҥkk+�����V�|s�`&��>a���� [n��(�3��>�)��h4T�m۷������lY���7T-p�}��n�
v�G�T�^�D"W��d����1����9s͐E��(+m[����H�
ߡK/��k_{�7���/����   @�eE�n�q�Uo����?��|fkž�]�v+�lz��/�*�� �������رc��,ʰc�sc8q�tX��l���|qێ��뇯��׆�ьAl*���1KC�ŋ���T�N��}��y���	W//\ZY�X$Eѐ����t����LMO��K˩�_�,lyu��V�6�[�����^~�,����:���,�Ibnr���~*��Rw���y|ǎ�ǁ=���-��������b��   ��	�y��c�u��~m�H���l�v����,��t�;����ì�L����Ç+����C�n�ݳgw8t���c���ի���!m���7�l���DLG&���'±G6�;�����z�^黛�2��,��(7��<�����ư�pvv������Eq����͚�{��-��t�z���T�����\KץJ	<5�����F����m�ۑ#G��?��O�D�Ab�����4�   �痀������6��_�m����o9w�l��
���E����7�w�u״ґ)PMY��p�5ׄ�����f�ݻ���j��۝�p��W�$m�?�	LY[�/K£�	O=y��|lc���j3�"�,K��n�͏V�W)���ݓ�z����RC�U���W]����;���}���15��;b�}�!x��x�i@ � ^��������־+�^<��n�}!�+���z^�o��q��?/1��Z���뙛��e�5����m
b���a��u�
O�$3WY|'�<Ν=ڭ�X��rk��@�C��m�:V|B�w��zP���Q>�*�U׿����[��|�ϗ~f�/�߄   @�eH@n_��Ow:s;��͡(�>���I��nwv˖��F�ۘ��O�a�ܽrT�L�4�0;;�GE�k���c�nZ�~5�[��<��p�������Rò��,�2�ʏ�)a[�3��6��lҿWAnY�>t�-��ķ��[���pH��SB�~�i �   ��+�:�pfjaa~feem�Ә:�5�WdIv�����<��4�23;�j���VVV:�Q�P���������5Zf��J�5�����1�[䣘w7SڱAh�ZV4BAn�\n��|�%�Ub��[�"�h��y����W>��w����r�/��_=�@ ���H��o�=}��Ls}��f�/O-,l���jLu��Ő���$y����W�$�)w�v{�̿��X&X��f#_��=�"
Z��U*2�+��!��exdo^xB?%��A���)�B8x��Ƕ����}�{�������z�޿+)>@ � �E�(����Dcjj����ص�����<==s��tzf&��VtBb��A?��E��3�m��e1�������������d�xD���[��J_w�u�`˖���w,1H� ����   |���{������ݛ.,-�`��y����r�Z��3(��4����҅��qA>��Ao\B���U�wg0���hI�b����*�ɏ8\w�������<�����/ۡ��  @ x!	|��?7����Ϟ>�}����NMO���ZtI0��,p-���Z�V�W�Wi��%_�~�?.8!��\dٕ�D�����v:����_y蛿������R���R-��   �-�����ei����K�0˲#�vG&�4W��4�;���I�6�4���X����+Q,Q+믂�$j%��RК`�b�=���{�^���ݻ�<p���|�C/Z85����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@����u@ �   ��	 xk ��   @ �� ��Z��@ �  P3o�@��   @ �@�V˗�! @ � j&��y ��   @�Z�j��:  @ �@��5 �C �   TK �[-_Z�   @ �� ����{@ �   �j	 x��K��   @ 5@��< t@ �  P-o�|i�   @�fޚ��! @ � �%�ୖ/�C �   �L �[� �=  @ �@���� ��E   IDAT�u@ �   ��	�go^J�a�    IEND�B`�PK
     mdZ�  ��  /   images/b13518ba-21c5-4f60-a735-1d8041d11d7b.png�PNG

   IHDR  �  �   �lC   	pHYs  �  ��+  �MIDATx���	�m�}��}��g��{�M|��$Se;�58��Īb;M�D�#"���v�N�&�ӊr`'�؉I��h�6���7�[���R"QI��||��<�i���k�s/i.,:���Q�;���k��^��   �#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   �4/   :��  �N#�  ���   om�����^��f�m#�  �I�z���'�X+���~����������޼u+�0��mc�6��<�~���~���7~�����_ϊ"�ײ�gk���ol���٬��'�|���[B�  �
��_���֭�'��_o���t>����Ai�6O��㬪�&��\�W�7R���e?kB��7򪪎���h�յ�?��ß���?��z3|Y^  ����3��÷n��=G��?d!�鵽��ˬ,�UQ��~��/��d��8��:�ě�Mo�x�����<o۶ʲ^����,��(&����x���������7ڿ?���"�  |����?Z��;����U������*�z�q��ZM�/�(��i=��Y��]�[P�BUՙ�ۙ}��{=���Q�������e��%^  �ߦ����_<<����B��Ъ(���An��Q�BS/�'c%�\�������g����Z�/ϋ,﩮7􊢲/���~���e��!���oVWV������4���?��K"�  �6����g�I��Bm�����r��i�[�m���c����d��,����&+�V]��U[�i������Mn�lgw�/)���+fs���   �M�鬧����l�x�f^P-��=���IUƐ��zv��k�)��~�Z�f��z���|6��,/  �o��yV7US4e�_��N�k�xo�f_h��w����(­�H���ח�*$K(}8y�V��������?����w~�w��W3|A^  �߬��SO[[[Źs��~��Z�_�{��j�r^ͳ�*��,s���WB^U�n���+vn���7�W��!�?{���Л��vM]��.�f�wX�^��Ex  ���~���W�d�lw688�Q�$7��}�/6O=�6�[��/��h���'�_|Zӈ�f��jl������ܞຩ�����tBl����\�?TM������}�������i4�o5���<�g���  ૞��2�qcp��-6k�hi���7KK�j2���٬͛���;�o=�}�lv�eg���O��;*bț�ݫ�z�כe����ŵ�W��GI�-�N&��l4���J9�g���Tڛ��I���4'���ݪ��S!�/  ���҅���F9m�ނ��ۺ~��ҷ��m�մ�-�֓��e�����6ͥg�����Q1)�v0�NV,�Κ�n4W��djwSIC���r���x�A�7y V�}cϰ���r�DB�zz�5F����+��mz���	^  �U����h��=ɧ���7V���l6����b�r�͎����?8�c+�;�yu����a�w2�~�Eэ�n��ӯ��e�gYӕ��aV��{Ku��泬Q�-GY^�ƶ���e���nz�}��ƃpS���|���/�?���a������~����ֻ�y���t�Ak]������o�u�|p����}4���Ν;���J~|tT-�,[+j����ٶi�)��O���G��۫�������������� ��zO=���p�����������Yx=g_XrU���fVգ��g�����h)+������;��㦗�%�|���R�n>>>��,{(D(��g��d�z�S�͛�߰�:��h�ݽs'[__˪6��ka;+����`=�ا0����j�ťKK�d2��~问}���2�&�Q^�����������������?���]���d*���������|X@A����V!7;::�,���Y;h�4�hgw�Y�X���[ߡ!���5'��KK���Q��<�=�ю��μ��t���qc0|�v���yu��w�굳g7�E�]U��+�i�=���eo2  ����|$?�^yxm��3�#��Ł�a���8Wa�J���PU(�1�KK�����zV5[B�ܡ���d�[8��1ΖF�L�������y�Ӫ^[������R������WYD%3�^ӫ���-om���g7S�qv����|ns���������7��n�������|4���5��᰹y�f�՜I޲�Ww=������ǳ�<�̿���;;��~�e���U=����0{lavTE�_�rn�B��<�u�x����o�7�픃�0����7�m��;�ͼ����{zt�է���}t|��{���+n�f�Zb�֒{B;�Zj֚S�nf�i�!
�O������w>�?{���,�fmu����W�.]��F���2���=*��~Y�>s���t2}՚�;�^{+���v������?�Co���G���|Ŏ������-�׍s��(p׿y������ �Uɮ����K��z��n�X]]����Umn����a~<g��;�p0���72��f�o���e�̮���77�fw������t��-#e���m����3�̠̠���x�^��/�ij\.b@+B[x�p�����:W��`0X�498<x��>���[h�S�ᰜy]�L/��n�����ן�f���W��=�y��f(�+p�c�Gu��?����_�/~%+zW���گ���?����
���_��}����Ɲ;w>�5�K��G� �l������Z;�3gΔ�q&�
h�.--��յ��T�«����V�d2����t_�gZ��s��l'k�ժ��$�Cm��N��d�^�\E�����~�M�w��W��oŶ��lln4v���Z�y���奕\j�TV�uo�w���R���}�\][Y�Lf�kCA^�~ǖ�YYY�4)I���>j�{u|���vs; ���+���|}^ǉ�u �k~��U��wfٷ|�F��o��������r��g�Ｕ�8� h4$s||�����sc[/;��t۶ǡ�B��|�(�;�|;���֠_nU��`0(�Ӊ���F���͢>:ڷͳ�\��yW�T7n�h�\��~���m���w/�G?�TK  �Y���w�,���eQ�X�X�'��ں]iu9-<SL&�ll�T�Ӫ@����׽�=��욮lyw�N����=����:��gh�#��J�_��g[��5���RM�{���@��!4�5����$�-�F��|f�?���eZ^�"������^�>V���������G���+������~��o�r�Fѿ�����ǰ���S��~������=�ؿ���W������/��W5��'h4�;[����S?rtx��1��
�]--/����}����m��6��VWV^UF����ª6�?�ZS�h�hXB�p�Zm�����ڛ7ox�T�nU�=���j�PJ_k��k�hH#WX�ίC��󐫲��`�߼y�_K���F?�@�{ܾ}�T��}���p���̛�4���>G?����M�[��,[8��ݾ>�5$b�QP��������8�?��t����W�ּ�9ф�^�W�W����U�3��|���,��6�Ѱ|��K���K��Ȟ�yĥ�b��`��]����l2�����F����ʹ]��a}V
��x����^���\˥u�����}�Y���
���+�-�Ϧ3��j8�5�8���:i�Ț8a�ƙ3�5`*�3k�Nl�ۊ�����ʲ��n�g�O�����R�{�r�k'�{�Y1����,��vЯ�㶱�^O���Z�\����hu���[i76v��͵v{��OP �����|d�����G~��۷�N���e���{[�w�据�*��u֯+���]��:�+�Z����]��>�E���;�߱���?OZSX�(U��/��<罯*wPi�����j��2�84���k��B���v�]V]��}/�pup�k
嚦�~����C�����V�]}]��������Q�E��X��4gp�k���v��C���ã��3��J���<}�����\���O����y��?���S��o?�C�+�C�n2i����|����F�@͙�3�ŋ�K�.U�Ԛ�3u׫��6�m�VϓVYCi[9����L��;;���ʒG��\;H�`����]�T@�Nt��h����Y�����zB*s0���gtwwW=���;;;�B�\�v��p��x�k���
h����C����*���Y;0tz�܂�����F��i,
�^/��@��kGU�����`�֚'H���k}�Ν|�B��>[G�Ϝ=�ˡ`�K=��/ߧ!�|پ�ϧ �kk�������Sdt#���¿
�=��z��6Z��g�u�v���z�ɵ<
졆����=�s��]k%?`���sv����j.U��L�c}�R��`�@�7j�2��<=���.ʰKס��N8�\�g�`�l]'�<����`0��e�G���@R�I�!�o��m���������>_9��`��U������s�e������F"b+=<QGډ����!�g>yx�����NB3[�֖�f9(��ر��=;�G���|��k��5�����e1<��I3,g��R5NڪZ�ٲzy��S/�G�q�������j{ܠ	��SO}[���_l<a�,��S---��AL��޽��2A����E�f���k�%&���� g�����<�ݹ}ǯ���|d״��N��K��9ш���ƙuz�wKu�Z�!�4qF�N�3��[U���m�>���`>�t-*u��=�N=����da�v]�N{�e��"�&�e������&��=�vͶ$��/�K�o��'�}�G�ҳD��^����??x�\��eǫܾt�^u�?���?=�Gkk����zr$�o��o�X �l8�2���zGU��e ��-���V�a�S��A��]�����*�Τk���_~��L��
R����B�Zg�A�a����0�]�ND߳X�֭��0�H�'}O;�>�!����I���r'a'�eP�;�?Ph*�8�^z�=������X_W�To��n;z��R��}?$�,[��(��k���^%���F��}��K�E3��o�;��Z`��n����u�C7���f�jh
��E=�
�)@��˗}�=�&�{�%�@[��D�i��R��Myhi�g��^��w���ݬ�y� l�:M��tOu|�����˯�@�F���Nj
�
�z?��n�����C;��$�Z^� l���9�󕕕j6�ض��ZFՖ�a4��}��z����~Zμ��^��*G�5�����f`�W�Jhp�g���h�{��m����=��^[-p�R��o/ڄ�L���_���g,������}v�zٿ��wf�K5;�~���	N-
�e@^*����Vi��7F��c�KCv�f����9��a�m~�6�~�k�{�5w�^{�~u�a���~�[�o&֒�l#�hTU��ܚ�ڰ���a]j�<�loo���Gk[&�@ڭ?���zO<��/q���nj�V��ƍ�����u��n���3�@�åAs����u��n���Z�S�O!uem-�X��D]�Bn��묮g77��x����]쭏f��A뽬z��ŋ��۷ny�,�گE����5�����zO�O�m�kr����놏~߻{����/�>#yu���K].�Ƕ��pWGX�#©��Թ�^���,u)�������{~V&Q����fŲ�'��w��?�goa�c�7<z������]�z�+��ї�������>d[j��C����=���{��^�x��֑zG�m�S�_��Q�廟x�Y���jc�Li�sptx��d��F'�tjV� ��"s������]�
C��rM���7|Y��^[{]L=|+ .�F]]]�҅���Ǟ�\|����{Ҵs(��z�L���<��*kM���li�d�i��v PY��·|��>{yjv	m�M����ܢ�[�u�U�hZD�յ��a�k�c8Uֲ�T����g��k�(��u���~'�zC]o��4��;	xT��J6��p�<��f˰���TC��Zh�ȧ^S��������I#O!6,˒�Nx]T]�<��'>�P��O���V^����(�$��캣6���u!��R�]om��t潣��k��^ʢ�W/�zx�84塾V�x}����C�I㦊�a;.���^�]���>0�����s��A��N�<՘�9�xJ'E�(`����5=[1�K���ė�i�x/��[�;�1dǓ���dg�N?~z=���!Z��A����9􂍖�ΝG*=��X��h��sȢQ��|ړe?�>��n.=�/�uh,�2"���_���7~��Q�n�O4z��1�ʇ�>ի�QjD�+���5�T�f�����S0W-�혽#;0���C���-ˁm�[����+k;�Gv��7yy�ֵ]Aډ��qoП�2u ���Zi�~V��Ю��6j���NG��p�N�#}�fi��V^c��jk�Y[�/�9�\�5�/�hϞ�i�Od�<��/<�{=������+��ͭſ��m�[+C�>��p2Q�'�A�l��(;����l�7�G�����Vϛ���k�<����ʪ~�X&�7�~�o{�:7>��������Ǜ�l����ύf�v:��G����ht���~��X��pҋ�-��h���p6��ً?�u��N��`6��{����?[���Sf�|� }��>��n�\�ˑ}�}�A;��b��I�ŗ�d���������x��Zí�z����hmۨ$���~mڶ����rQ.���ӷs���Å���j6��&���Q~�Ν�������U��6�p7�s�nJ��;�~�[_���^}]�eG�@������B�v���]�����|��9s6{���|�j�������ݺIDm�vm�lvəL��S�׫/h�s����ڮ�S�R��������>��x��"L8����c/��K��E#���d:�k|虾sw+{���s�������}zx�c���{޾tns4<>�ٰ����_�C���;,��-�>����c�|,;�|~�����^���4̬�������{��M!:5�E6�����A���w_So�BV������ܹ���x�h'�x��B��4��;/����[���u�V~���|��f�;2��~��������W_������e��m�.8���
��S�������=�+��@��]�5��z��c�a��\=��bn�Ƣ�>Q��Ϫl���S!H�A�⁨��X⯧��%�ݖE� �4�љQ��/˼5�P�����5T���3)+P�US��H���=���4���e�<-��q�׿��O�iOX��
�)��=X��逬Ю�S5Tt�����i�S`����i��ZFՆ�v��P=�gϞ�bi�Fr�?!ؗ^+��p���S�J�6�u�co!�~3�����Z�:�����"LK�]�^ �稆��2��y��We
�ڟ�?��F�C�Z�J�!�嫞�ڷ�\w�wz�PH��^S�[ˣ�t����Ν[�?Z�0�I�ˢ��5�-U���w��i����8P��֥:����M�N�~����'��¾����kT>��z�QZOZz���ԃ?����qR�+������,)��i<ݐҺM_�>�I���t��Ok|g�����wSǹ���⢥�'�R���p���7��gZ���(��k
��?�T8g|��S%Q^w��֫�le�f�sϏ�&\<_k��4�G��8<��Tk�㣱̮2+���C���lZ�hZ;i�u��m�FC���X�J��X��f�5\������E�����Vu�m��]4��� ��7+zŴ�TX��	4o���IQՅ-�h0��~����m�ׅ�O��DY��U~��l�h������lP���t�����>泽�-��R��
{�fسw��jM�YQ���O{sk�i�򺢢�E��X��W��04����h�Q6�-�,��iE�0U6�-��zM3�UYU̧����Ӄ��W�Zc��G���p�{VG�dz<:��e���j�.�k3=�`e8��{��[�ɏ}�G���U��ٱ1��u��'[�v���hǃ5��z2k�̦7��q�Z��Rê��6���6�O֨�k��Փ���onY�>w��M���n$֟q��N짞���������_k����^�u�kUϩ�q��V�����Pݨ��o��M?oZv��aP��t�޶�c�Zh�{�nv��,��
������<��*?��`�e
�:����xٮ�:g��E_ޢ���Mm�x�E�z���}��z\7Ξ�nߺ�Y���x�UU�!�|3�΁�,�|�M;�Z��;��5][ԃ��8{�Wl]ݭ����[؛x5݇������+�����[�ް����ի�߱���M�����������wd�{{����ZX~�v�#�����ga�|e�/��[�HK��:���Tb~���1}��,�>`�R��h��T���Y�'�.6?�?�kR镕����������677K]ptq��������vqU�TX�0H�M7j����S����Р���̃��o
M�����Gٚ-�BT�I.L`��TI���g?�Y�W�/^�ϧr�Tޡ�l��B�&<�PaU?S�d�u�����{�z�=oZF��omoś��x�����3-�NZ
�
���!7M����&-��kZ���4��'I=�
�!��_W7;�eW����b�ƻi�$�ƞY}O�@a��'?���z�0%]�_ײ�w��Z/��C��ֳnrX���~�����k4����������P>��׋�/��AK��Z�z_��<��%۞��b�y�D��7x/���?��;K��!�R���*_'MzPx�Ի�&AW �6PcR�e<����Zư���XU�ƕ�᳅�ƍ����.i�FL��"9�7s�O����ÁOѣJ�~1Q�@���s}�.6�Imw,[񩆴�n(��z�t�֍��M$a��d��QjP�z��ު/��'�6�dFǺ7�bX�bϏ���+)dO|_������Ko��Q�آϛ�#�2���S/`i�0,�2z�U��������N�q&[�����u2_K:6��X��r���~F����#D�0к�s\܆���:7��L�Pu��F��ױ�-��3m�,�M�S��7\�9)��d/�-��tПv������>�dYx�)T����y�r;���Ըj�6T)���C����׫����M�&S�J߮{����as�������(�y8����U�3�FeQ�m�͛��p4·j��m}��W��GiT��.�Ւ]!�H�땦Z�W����h6(f����}֨��<p.��T~6�k?��+?77����%��R�u*��x�-Ν~ޝ�f��Tg�:�����sQ���S������Jĩ��t���ʶ��>�ܶ��ř�a�Y�)W�M3�Mgc;O�'��ض˼�+&���^�e�l�_���z�/�ǣ�5(ʢ���{��Y�������ѽ��?��O���e{�Q]����w�����.zCUYD��>��Ғ��};g�!��\���S.\��y����^��5��k�^����ϛ��s�ƞc�{�pX��g����Fo���y$^=���o�G�y3���^�L޳����ɾ�unq_��o�-�[�����7*���5��|ue��r�w|�������OngoAoj�|�r��ϖv�>��s/<q�?���w?p������)Xz��s�=��d�Чq��i��6��mٙ���ÃR?��N�
mv�kbU�`��;MLG� �a؞����d�Q�a��]���	�NB�:
�*�Po�B�vv�"hH[?�״ךF��J.�Ë�K�`j���Ԕ"^�z��������=�-����(������P��=�}�%�:�ؓ��)���7̾�B���O�vN�y�M�EP�8�R�n
�
C�����S�{��K�hi[�$�C�v�N��Zn]L��T��?u1�����n�e$C[�TG
@Z}ch�xAN��0uJX~}�<����Sϥߐfj�*�{*O�.볅p£�h��!M��7��xE3Fh�J����z+���*�IR�E�JU!P�YW���S��^�>�k_��r�n�X#�ϥ}Oˣ��'>�Ҷ���G����}ݶ���Xʱ�lZ�cR�zZ��� ����x��:}b�:LA.�:���C����ɔ�:٧}�P�<�}�R��|�>=N\Z.�ꩌ���v�´�8�[�z�f*9]Ýz����}(�ظX&���y�k�}R=4�N���X��+K
���I7���9��,��./��xcdK==�KqtF�S*��c!��7.�K��^�D����s���-6�I�%Yz�:��X^�b�o�f�^D��,����Ư��zzuG�F���ì)�b�$s%���^˩�;�}�º������b��m�v��Ξ�����֫�R��w� o,��[��*��B�.b�Ow�k�N����t.��~�T�Mׂ,��~Vewڷ�N|�2�1��l�:bA�K�4�����`����:ɨ�>���j�������u���f�I3�����a*�C*J��d�=U������c�k�����,Ko��q��U��a��x`�U������Mq5���;��^��]�x!�Y��ͫ^�wo{�;kf��I8�z�Y�O*k�WN��F�:����Ѡ���M��,�_g�č���`8���P _]9�8ZZ���Uu�W>\�����ny���gׯ��]�t�υZ���\��G���%+���צ8���F�λ>JcǺ��Օ5o��u^ZU�({��>b�O��l:	�A�á���h�%\�EG���(�k�2�*�;;�'-���k��H�����~Ly�U�V��LI���|�C����õ��?e>���/ފu�oj�={�_7�?�����~��X-��W^�[��+WF�����I;س�=��b���������^}�U�@���Z,־������v TK�`k�jԍ7
ӈ����
m:�h����NT^{p��'Le�9�d����ð�@�)mj��F��ի�� �_��_�/�wIAp����on߾�ꤳ���l��<�
,�f��p���^�u���{T��.��,$[8V/oO"�㐲z�ԛ���iBv,��$�n���t���l}^����B��G������^�rٗMR�j(�X
u���+�� R���3g������X�����&�=(:3���P��4oy�3�G'f
�j��B^����Z�\�ԯ�z�x������FL�M�O4ڏ���룿� ������w�?�������Б���O�Q��C�V�b������GK�<�k��'�T^����E�~Fvq'l&���z�N�k�nݺ���Cxn����~��/o�Xd�E����^�12�]id$� �3MMW��8,��o�0�=*S	ʪי��>��O���X��آ|�,A�?g���m�!�67N��_����;�&�Tc�?���-4����,�t�JB ���I'j/�-zHO.��B��h0��JJ���F����:�<.w��zī���˗z�㴈Y
{��)���n�u��E� �2W��y<���������a��b1�H��K%L~��p���4��k�}|6��)��eѺ�q���T���ŹK�����0b���c���˴��频2����/\�ؤR��˫�]�p���:I���oW�#PM8g�͘޹1�&�w�Ӻ	�V�aw�O´�E#�v��U�S��Q���Sǂ~���<�@���.��E��okk����M�/4��?R��W�d�̦�ڰs���/\���l{�:Q��^O����ԍ���;NoiT�,�Y��̏���}�d<�o��g%��j�	K��O��_�z�l�-Νj�k�L������fב�xcVQ�#�;l�u��u���z�y�JSs�/a_׺����Y��GZ��Ml����"�~�4��api���i2����ꩴk�N25�l����gWy��Q��&3?G�q���0����p�ѳ�׿w�xo��0��s��ѵ�	�65켬�U몪C��v�����������c6fH�����5�pi�/J�|�N!�z�eo�4H��^��zx��.t�y��c#,���s�=?�iƲ�虧���7��~�/��_����h���>��3ӷʃ)����䓟���ő�����|���M���ֿ����y��K٧?���I����e��~��ϫ��o��ڥP�Y^8w^;V�D�"�^�Z� ��cvrZդ�
=vQ�4��.�z�ّ��y��FAHñꎿq��~+_�Bq�����P�·n�Ց���5�t�bx^ʃz�;==������A�N�]x��<$y}�}���yo���*��^z�j��w��B�-k�=p*�*d|�3�Y\���w�ν������|���}����2��L��؂��Q�Z=�['f���-2.��^/��Y�լ^�F� ꤥe�t+��b8�O�#��7��sj��� �gv4�3]�p��r�pL�'�xh�r1�ً3>�Z�";o�]aL'B�z����t�J!��g�3:��*F�?�s/��.��t�K��ԷeхFu��	9Wl�$�Y.�K����RxJ�o��ç����׼�A�������!�pTOp�e3<h�`ɾ��g>��VￖA_W��BR
���F�P�P_�q���<��t1�{�����m��c-C(�Q���_Lg��n����~�>�,4'=�����l��3�Ts߯�p���4�3-�.�jx�ѕ0u��{���=�E�C׋��`��K@�����|��=?��m��c3��bq:��^BzG}��8cI*Yx�>$�~����I�j*�H=�u� �=���i���Ϟҏ�w�X����R�tSlz�r}�E���
q^��=Qy~�?����S$*X�a��T��4����Ǜ{�h�s�=��T���|
}�~��Ҕ��g��pt����w�Zibi�OU�כ{-c��=�&�fִ��I�V�M���Z���k<�s�]�
f�Hh��-�f؎t2�ci���j�_ͨ��kD�=��o�/����E��⥋�vwv�5uD�>O���J�q����l:��Ԩ�yR��m˘�ȕy��`uQ���d7.{��ꈽV(��4�̭x]�����!���5�u}Ӄ�,�g��G^�����+޸�y߽�UǛ��>K�ܷ�,\�.}��롞�����SE�횽`4�ٹ��������7G:w���F#���/���r���k{gVJ��f8��`׆�����ً3	���06d{�8�T��A�Щ��R�F*����m;Cb	�ɱ~rJ�
���rx�p�_�z��{VD��p�iHei���ק�e_���ܧt�3�}��;:U����-Cͮ_�~fk�����~Ys�?������ޮ]o��S��-���c�Go~�����a�#7�ي��ȏ��o�����|�{�����~�����r����	Uh�<������?����}eeէ��2\�'v ���,-[эB�]��l�W�����g��qc�ñz��*��_{�5�F3.�e<�)�gO��	���l�+u����������K4w�nXe��'�L�a�U��"��vB�3l���VQнs��7����D��"p������&����ʕ+ޣ��jY=p�ƺ����P���~�EH���u�ࠡ���ʕ�f~!TN7�h��6R]�JO��/�^�>K�Գ�^j���>������	7ˇz���.���^��[��Q,IH�d�*gi���$݀wzhT�A�vP`T�������FF�6&�&�����Zq�:秧��z߲��^�k���C7���}��M�}W�j�ÂZw�X������������v=�j�脪m������?�r���'�𰩐���ը��_�{��|t�(C��5�vo�K���k�w|�wf��ԧ|��τ*���|U�<��:�ҷǁ-����X&���򗁇�����׋"�i��,�b���i'��*,��������2z��wn�2hY}z��Q�-b��A1����.zX�8$�����4|���p�Hurm,MHe�ϰ_Ws�	��o��A
ۗ��O�/��7��S?�z@��Y���`�u7n��r�´��!4��+�����kR�a���e���4�P
ӄ׉=�gR(^T@�龃8CJ8O�Q�S��xc_��s��M=�>:�@��ZE�(5H�݃��h�F����'.f�y��hAZ���L���=�鳝�?R������Ϝz�&���|��\S�h�3��59��O�a(�����5�n;�>w�\������������^X�[�}-�X��q��~7��xՊ}�p�I��q��Z�"�J���z�z�LGz���G@|��ҬG�S����z�0R5H�:���uGjB�sii�ܵk���Y����4�Nh���;/j���P��_�p1��qM*�Pǆz��������zGr�P����a��뭪j�����凉5P��>^V]�j����S�p�mm�񹺺�S�.����,N�Y�V�Zeuޤ�����554�c9R�ao�ޢ� ��P/�OE\g:/dm�q�"���{:�∠OY��|����ݿ����>�n�/n�tՁ���'�I���,�L�*�X��,����ܡi5Ká��h����:���7������?Q)w�=s���������G��}�7��Doz�m}nƏ�}�W���~���!��������T��=Ԇo4�9�0�؅m�\�@��ӆ�?�`�mۑ|m���O�����?���_nYtݍ76�j����o�1[�o�s�ӟ��B�O�a���`��RM���6�,����*�ܠ�����3)��K��K#�D�p*�A��f�~
G�~�L�a�j�����`w7���Uk/����x���ih�[�
H
��_{�C��O?���"�}��E��իW��vҁ���2�J{�$���e�^�س���V�~fgw'�\�'b��zb�5���B�.n�q&�4��!�4���~#K��N��>���u���ށӼ��Y�C��j�o�����x��dšv��?��gRo�/_�����c�z35|�ى/����Uk0�f�{[۱qΗU�&��u��K�M)k��'΅Ϫ@�j��Y�l�xhR�Nd���>ָ~<�춳��
�j�h���mg}F�tՇ���Ϸ���������~�Cpy�ԍ�M(�2��.�v�[��������l�{����	�a�C���,5:���Lge�Sc�Kl�j?W�O�A�]�z���q�muˀ�}Ɗ�E�b�/zC�,	U�����J_K�P?��rS�9�3����5>�|����tꦴ�,3�4"�P��YM(og�p\�a.C��h}{�y�/.,��gQ����c8�}���X����4A
Ⱦn�U޷sk*7й������Zg��4�C�}/�Cݡ�����9�{qyb@nJ@Ky����|5�Z�x�T��9γP����ң���K�TF�3��ЋJP�y*�ᓐ{�(Ќ�G_�Gקra[N��Z�
�i"��$�4�����W���9�O-K�<i$���ף�<��4�}Ҳ�O���у�⾘k=����NN��^���WG�-�p4����`�e�-�g��<=�Yy�*N�XW��k���j����+xC|3O��׍83�bV#}v����h�^K���E�S�c]'t��2�U�����qM�fi��u��Z�\YZUO�ȇ�/��Ӎ�>\7��w�F��5��7Z�䲋�/�yH�#���R�'�x����C�fo��:m�E�z������]�[��R��A��A��2�"��)�z�/�Eqj��GC���5+ܯoN�ſi�*n����=
~3o�d
N9i*�C�_�5��]޻w��lZC�o�.G��e�E��j�R�ؚ�W���ε�v����Gٛ�+x��������s�,;�������}���?����{����6w�wsk}����
a�5�B����co�?�ܳ�|i��5�5�c����v6Z=c;�߱�',����0֑ܳ�~!����[����(ֶ���ۆ~�.�8:8z������Ajg�l���@7����Oeѝ����'�t'��Q�eRo�����&�p�V�p�=��$���n�X�Z���}�{��:9�"�C�
7�9�ހ���z��\:j�_e$zʚN��fUua�,��߱���I�xN-�B�[�8N����G7��	���Ah�ۅQ!k�J1K��i�R���xײk}�b���,����~|�Z�D=�a�ǞA]$��6�LH:�O�g5$���f�:�?�֝�N�YR�`?>�yb'���O�##�;�y���t���UϹ_��w4#���W����?�����y�k׮�6���_�p��n�)h�E�X�Z�:�Ʃ��������K//jm�}��>��؋��*�Ϸ�h���𶎴}`�yE�OAZ_�y��"��k:��=��P�H�[�8N���R{�d�7��{�E��rORR@��>�������_|�?tv�Y���,(��~{33�%](�$o���z�:��=��n6I�e��Lә� �z���)���>N�A���\K{�5c(ܲ��+B�.O����S�ԥeN�M?5�N��Ƀa3rě�⍘�7@�ϖ~�V�4L�T|��7��M#X�҂<�P7�S֧fr�O�Զ��K�4Yq�C��������>O�/ͪ#xT���,_��'��T[��C��5�?�����e~��{����>_�nu�}?N�φ�ºN�Bi*¸��?_o:��=���p��#�c)Zӆ^>�Vp<^�ӝ��mo˿��ɍk�Ҩ���_��ë��ڷ����~|죊a��8c��w��i�K/�^l�?�dȽ��_.�}P"M'Z���F;��7͢�(��сT�i��;��>��:DO��9�gc�Ǘ��y�]3,5*yШl]Hӈ���z�h����/�����|({��+a۝*�K7��c;���i(c��ڥ�@�y��W�˛t�kR�R�q���ٺ/��TB���E�|c��j�ziQ�U����<Ue���6���+���"�T��#z�mg0ibGђ�����*Ubf׿fue�{Օ�V�W�V�J��k�����7�ƙ3��.ՙq����or��ޏ��ŋ/>���^�����m�ǋ����x��t6_y�w�~��G�o㓺x��kʦ?6?r�T9�.�ڡ~��{s������^�oݼ�Cۡ�/��/=x��?������M�8�w��������>��[�������n��d,�fG�M3�P����d�����v�<6���Ps�.ښ=}t��]��T�g��q���"�y�t(�̠Q��h���4����ׯg�iX������0�n:Jw�~zY2��.�:�]����$�rx�}O@���v)��O\�w=��+�t=M�[�k��O����Y�LS�LgS�S}������'�&�/�v�j�8���T{�S���9#�g��Q��eA�M��3�%~�p5����lt�F��EXW���*9� mM��j��6�Xc�;j[g:�鳫�F����ۗe>���#�� ��w��i��i�ܯ�k��y8<0���c]����=�y��w)ܕ����'̉��I��q��t��͍z��0�����я����O��=�xͨ�m�7S�k��.L������y��G�%�	�7�~zXI�?��N�8��=z^FT��S}M=����iĬ���@U�i��>ǵE�~��:�����=����pmxl�����&4:�z���
�!�����|رi7�itf%ֶ���cT�S=���{�^��x�b�:N�;֠���)H���ѣm�3,�^��ӽih5�ϼ������E��Eu��A]�4�v
G^�Tᩄ�t"�w��".��J_�<_�y���5�>�2�(k��IH��P�J���T!=-�d�����5�8O���+��Ѣ�$�<��W�MC����z�oh?Uc6�]��[,ch���NǺע�0�|qæ���m^/�A���&3��5��\���m�q���� ��X���Fc�Z6�W��C�چ�75�2<;��Ž)�<��G1 �M��.� v2�LQ��ԙ�$��r���X�s���<�h�)�)0i]�b�Yz�����G#gi&���5&�z�����T�WqE�K��e<��X{�������T�f0	3�.�K�(�+��G��]��ty�z��Nu��k��
]>�X��J8�S=��>����9�#�?�i�w�t�ZwGǇ>z��a�L��8O�(����f�qX��X��s����<ͦq���]t�f��ͼZ������0�r�6�ꉍ��$<��/V���c6��//�(boq/K�C�s?��|9Z��ry��m��M�]}���=�?��зյ��iT2<�`���|d������7}߯H��{�'�_���?`;�v��g�LU����l�޽m�iF#�^�������T�r�����_�������������p�m���g>�3
��p8ؾx��g677�l]�/���5��K�|�I]������W�u�褅��[[[�wxttk��[�W��~��j�1o��֒:?W�u[��Dtv6��_5��u;���oG�f֎Sv�|�.TM�]�K����-�X�(U��'�褭�����of���N��¥f��k�U�_������^�S����u;����/����&����`�T릇�4��y^���i��b���x\��G���4_f�}��{��������X��3u����p"�g'���:��p�+��]��G~a]ZY��>�oo��i7�ז�~,޼h����Lei(=�(�Z�<x��-�I�5��4Zjz�����BO8���}�s=���T?���O���2��u���ڜ=s&WӉKӔ��['�]�z��ᑇ�6>�lo��C4M�Bp��M���M;�o�Os�څ�. �d��4�K�����z��N� ji����q:�0r2YLI��LAV�5a���������
�?��0�F�Z�i��zKfވI� u|��8�z���>����v�0s����Z�aj�P��!i����� za=��Ƃ��nj�ǯ��c9�Ɩ9�$�@?�!?I�G��i��R-������x(�Q'=�1>v[�'�N��W)�����H�L�������n�Ұy����j�/�ZOa֚c�)<�z���	��r��R/a�=5�Ҕw�O�i��<�_U�Ǜh�0k�b�t�����Yf��<�Sk:.�?+h��~�È��Ã\TG굚�}������}�Nx�Of�9BC���������4��0�@��F��p�r,'�73k6��;6��z�4B5�fa�����"L���W�x܄2�����l���\�;�1͋PJ��~SW�1�z8}�U��*uO�}JSօ0\���|݌,���^w��H�lј\^.c����W�Q#n��řw¬0����E�|
���J'���1�*��qs��㾌��fu��7���8E���7�@Ϯ�[���p�\����9{��}����p�"�i],��4�G{��7���ł��{��L���N��i�[����ec;�i���{���Y�㩝W���wըn��w�W$�N��7O����[��*��:ǫ~R]�z5�76*��~������S�h]]�
 ?��~2�ƫ��s���/��ľ}�~࣭��AܟxS�e�?�{�f�_���3�.��������N�v���R�4˳^�ԫ�%���|�-�����;F4�rɂ�Y;�k=^��|:#;I��gRǓ��(8ߤ�n�y(�b�!r�7��ԓ�z|��Z�:ع�PQ�H�S��YMOǉ�!>�z��O?�XA^�_�~N_��B�=�i�m=�U�r��Z����h��YY[���4g���X�^X`,tr�3a����·>R��*��kě2�8�Yx2X��-�"ΙY�i��~a�J�c��TU�Qp��$D�gni��fP�k*&��$���AM�wY7E�gS��w��w����u]� �O�K-�z�Ğ��?��\ܬ�j��v�T�&H
����B�����wa��T�aL(5>��PW'Sť'���>O?d!�P�BT�6,]�ROc�b,M�������M=��җ�����O���0�9iz�4[F�S;�����S��y���,�\��
��{ol�u�	�Ϲ�o����T�R�ed�m�8�1�M1V��h���p��A��?:��#��+���S`A��*
n(O�O��Yʔrz���;�a�^�Z{�{^�6`)�vq��~������[k}�[Pq�c3V����j@�ʼU��)�}����~�6����U�	g99�¡M����<i8���2{�q|�Ț7^ x5�TC�]1�J�Z��J��Q�ٲ�b�`X��F�~_�)������)7@Pˁk!����W�f���֊�/�}�~U�7���0P�Ds�ה9�[�f-..p 	X<����R|�ڞ*q4s��pf�	1�:x�G� 4�xv��]&��!����mܧޯ��80�5� �h�U�g��'́��y���e;O�Q[���*��yJ)�R|!Q��R%8�34�N�h��	�؋�T�-�xn����&"O���%SiN�89Wrڕ�Z}��Ca���8.�\�����V�&T�G���=H�2fRWZ���"1�%�%P��W(ϗ$�c_t�!�ײ�,���I<8��'f�ֈ�����s��Q�.��K^����9������׆�7I�=�w&_����y��uF���L)@~��Qs�˿�y��_�ܳ�xP}�?ŋ��ܜ[Y]�w'K�^��U]��k�"}@F�+m ��z׻�y�q�T.._��n��[��X��o'�h���آ��Y����;�^_���M�y�봉���:GR��Y��~# +Z	L6��bm��@�c/;�@�W{�L�#
δ�P���mӵ�;�ori\�p�*[*-լ_�O�sJ�u�zI8�}�ɨW��p='�Ђ�j>�%��%�[���$S�
&|�z�V ���>��"*lkvs���f�͘����1J2�3,/-��+,ZK��t�\ ",��q8��v4����B#Z�W=����lxNP�7�c�kA�/�V�҂8���)WM�	�0�l���ޮQ��PN����E�*U���Rx9����I
����$!iF2��y����z�-��qQo���c�
_)�7N��w/^�Xr�q�zp�<��S=�
\5��EK�Q���^�7����=P��h��*�@�� ��Ӱ��2�z��>O@����ڔ_�Y�xx6U�k}f6�cƱVyse�7�<sMfU�]U��rQ�QC�")7�V��R&�����PVVy�{{ݒ6���}5�f�(��V3I.1<YH^��oD��ŋ����{���~�O?uV�\�'���H2>뵰1��D{\��dH�E����H:E�1 t�6�g���~i��!N�uK1'��H�e�~����$&{~�xMlDӪ�p����J
*�x���.��3K�M���ø�{�`��Z6�d fHN��8�X��aH�(���;5��'N��H �ن\��/<��P_"�=�0���4[IA�4�W/릆0{��W1UϬx��F����5\Z�Z� 	�(�?��=��P�]��RM�?�� y�)�o�M7'�6��3�����K�X� E����>��瀤gx������S��U+7<z��/sw�=�ȱq�:(cZ�{i��D;/�M9�䄍�̙3 �0�����ş�&�a�fD`��4���N��z�w���A�UX�cڞ��s�>��D��\Q�6�0>pdm�Vwas��4/:�w�Y�������px����8���6�$�F��]�E�C�+@�hH�����h`�D����n����]C�܋(P7�e̘��Qšm�*N"�����3�"�b����ӵBV���A�t;�!mqin����k��H{67?9k�� �ܺƋm��yjX��e�
�W�.���no�y�,��ڹ����>�hU
��Z�,j��i	�xS����hcɳ	O3��V:A� �S��z�8�륅XU�M��G��X��V[�=�5M�2h4^�K�
�|H���~?�<R�0/����qQ�׌M{qe��r��Z�s�9�
x5��@T�'�'�K}�Oi U`�T6Q��@�ЄD}��1��Q8)$����+h��Ӫ�A�

J�p\���{vRr�(�CP�����\�v[��Ā��}K�G<|�m��u��e�(rB8�D �/�T��}"�1��+c�G(�������<��~��kA�/�zww��8 � ��c�vm�s�����m���R&�i�$4��5/�F _x�1O�|B�ի���D����]dp	�ױ��q�x�ɲ��5m ��$j8I��0����A��y��x���uդR�A,����zr�l�������3A]������b�&�ӧO��	����F��u@��U�ڒ�¼w_H?�5S�����M��,�_$����_��z��Z"�@���}!�\�N��{�����|�ڿ_�^���R�W��R6~yV����؀���*s��V���Κ�H���ws�w��ǡ�UN���-����Q�U��}�{�S��8{/M�������&�]��h@�a���Ewms�';����>��rg��A�n�:
�I�ץԞk��fڦ��|"��P]?4x��S�������	� ��׮��^�����L=������ţQvSa�L���(IeY���9������~M��A�D>7Q:b���O?����d:t�l3mj���O@�����yD�r2�C�UȢ�\g~ց���ȱQ�H�q�Z�v�[�+���,�'��m.0��A=�hL��Jf��A����U�1�����G�d�xʂl��#��� R
��C�� A7P�8��*g��݃@|Պ[b�*jx�)(>���Q�)�
�4/��$ԹTR���z&��(���q��^��3x�po����7���V2� �;xmk��Yl�x߃GN�pm��l����S�����m���C�&G�$&ڀ�I�{fwo���(�V��~w����`��-W�	-���RP���1�?�+�O��G%�E��mP�$?���:<G_i&\�+ҨB�״�����)�� 9\�ܫ�TC�Zښ�9�m�"��ɒ�۾�w~ 밖�N��R(��Q�'�\TP�k�6���q�kԾ�A�C1�v�Ǌxnc.*����JZ��Ӓd�R°�`�5��̫�.}��3�T(c��$�:I�D�5�V(㟍e�O#?�r�c|ćK��Y���b,
,5)K�4���F�^#�>��{���o�u�O�n�D׃��~����ί� �v�ZZk�z�>�$��q���c:�Я5`���=_*��ǣ5�A����[�O��T�|B�*������f����>V�B��]>�:�ޭ�k�)��? 0G�F#6����#�0��'Yr�ԉ����|������^ॉѦ��L�҃_���2P	mtA277k!����F�?����g>���CG�"@\KWo6B{���%�6m��U�*����������F�����C��C���- �hԊ��W��=��Z>7�$����Vo؟#�ݡ�F+�1��M�����*mlmZ�;^��Ԯ!0����?��Jy	$�j����ı�ʍ	�3u�����̳�`ۋʋ�&#��j�2� �>{\A''��r@�^��Yz!u/�B���׶Z��$Ud�����q��+��A���1�@Ze�'87x�
j"�9��X�,W:hv:�86~,�ic��Ƴx;E
��y "�AW�
�X".�$$���|��7��4
�@F�u�W.�A���M|�������^��d�W��5�L=˚��*�(��Ew"]0�*�&X���Ox�h��c���6M\Ԍ}���"'ꥮ��YEI��2�ArU�P��(�
^5ζ�%����a�!��Y|��5vz�lRJ��T���T������'���0D���;��@�4�T�t�hw��\�П�:�=���t|Gx��q�M�-d<f�8:>���^o���S�c,`���	E$�����z{{YɑքG Z}��)����no��9X>n��fN%A1�ʲ��7��zI��ƀ7���z��W�0Hh&26N�9�x���2�Z�t�*h����O�ד�ÇLg� ��,Giؘ"���7��8���駍BY`n<���+��V��͐��Jz����x~��/�$aR]Q��C������f'�-�޹�����/8��W�+�R/z�ɖu��%����M��c��x$C�s�a��������P��|c7NF�;9��G���#�?L��ܠ�� o�lE44�Ӟ��4�z��<���j$H>������?�y~�>�gX�-d� ��(`1���{�'�x|���g�ɂ�h`�O۴Mۗl�?l��v=_{ee%
77�B`{�ZE-M]���a�k�i��27C#C�h:�V�z|�6:T㙣E{�֐9�z���(���QgfF4]=���e�j�Є����K�߱���{RLtq]��|4�c勢i$.6����0t�g��$���^ˇK���PY�;３�� `u�G�z������W�{���G\+{��6��^$�b��r{O�r���hm5�7.��Ǐ�=����޴ܭ~7��ZXє~���E�i�ޛ"�n�i&|ܘ���E��M��5�T%��r��U{���%�Z)n���eR_G"����ꨣe�Fy.�R����'�D����d-|�:Ԟ��Rm���V�D�e߈W��/ޣ��%+����.��0��=*��8v�'����%Ƌ&l+e���&�<�LY���c_$+��|vf�-����}I`��d����Zjzݤ�__/'?i��Ѡ}ǥ֋��4=���c\�Ӧ2��$���]��&HE�Y���@=����k�C��1��)dp�_��G1���9���] 	*�-�Js���s�uVr�J�n�V<'K2�im�vH'+�:�T���~�+F�P�X	$ �q���@�̮�|~+Ip_���`{ߗ��
$�W5�	ߙ;n��<���lH�y�|����%���G�Diw岔��1�#ǎ�PZ�Wx?��G�?�Б<�F�}����RR�b�8A���h��v3�:�"��h{{�^�|�B�Q"�i�DI`�����Z�S��K�]��3��N۴}�/��F�aj"W �{�#������4��v;�ȣ�jQ��jP�D���4��f�x�4BW�¨�j�e���w�Ȯ�]�
�B[+M�f��y:�����8ɤ8N���f"�6JD��\���L�&R�̒:�E��R�(!�y:4I�	�0i����c�^q��bS� �?��<��D�#O	�d�J�aɳ�u�� �i�a�z�������Ϩd���{��r5T�K��a��߃r�a�)�W9�J����þ�ɹzg������&C��vv�����G��֝���p���k�����xDcӺb_�9�H�
�7c�"_]�DP{��T���o���(�o �N��">���e�� To\�`4������jVc������SC��B��;���l�#t4o(�3p\�C�'@wDt0��Ƽu�-�-ơ�|��ﯠW���oL�p�+�c�_ ҌK�3J�wv{{t,{�葬3Ӊ��q��NExƬF��=n�|�I���#<��#e%�mI�f�*ԫ�^��pv}��$�8����"g��<^-�˰fxO4',B]��`�8�>2!�B�Ъs��%FUA�z{5�
;*s
*K(���w�h <��n;c>��O0=f{k�����c�s\�7���=}��gb�hҮ_�}ŀc��&�p�E�1�������l7*��L$��\�����h�9L"��h����g�=�E��q���p�] kk
x�mڦ��l���%�n����)���s���kbǱc��mnn�,����l�vhi��qL�?�#?�����dY�L�L���<ws��Vi�] �8O�w@I�5{�'��'LYa��(zߊ���+��M;&���I�V�d��N���95N� ��z�y�mUjO5���t�Da �� ��=p.�vW ����*l8��MTu�o+F_��y��H?��F)�����.���@r2D,��d+�M��ـ�����������_�@X�/�j�T"�S_;�;\)K�i!_�/�<i?�,Ss� I%8ǔO�d5�$���p�cP����CN���@nk��*��Gu.��uy<$��R�$I�'�
sR,���,xԹO���'rĪ:�h:�g,U�f���T R�U9D4��10;$��x�Rڷ�-���B?�m���������due=�x�"VgΜ�P*�D��p/@��C��Jǁ���U)emY�4"����e�Ī�U@�$�~�M��RH\ ��}?)=�q�y��Z������ �˹T�u�]�����zn�F�4�ZÉ�7�W��fr���:d�~"���z��;;7��+A��o���RTL�Wx%��ׄH��x�@����y�,�ŅE^8�Ñ�ag���Y�ow�gqJ�O�T�q�^�l�v����{>iڦmڦ���%<�����'��� �?򑏄33O�<�t:��ʕ+���af��F@���Z9�n!IH{R�y�&���h����y���!Whk9B�u�1Hw�`Z���'8��h��K�}6_l��}[��dpH�0i���z2��s��q�{�/���忭��
}V��R�Jd�M
>c�������GQH�L����򯪅�U��M���{�Y	���+y�*� �E�G ���&���b
MH�e)3\g�<;��z��ӱp��Vm�jiaX�_^�D�ܹ�mH�E;�e-ẻ��+��:p��.�]2f*�pFCn x�b�G�\ˮm^��33�S�.]Ƶ����ozӷ�'�|J0��܌}�+��9�H����� �r�[�������fsk���x�����%#��^��_��m�C?�GQ)A��O��g^��������FB�<�|r!��]&���)T�_�M����*k�?��sЭ�-��:$`�9dp��`<���l��"BR����=�(
�f��ǎ���+�4i�4!���T~qE� u��Mv��ǂb������-����n�^/.1k�ӦY�6ɂKɚ�J�M۴M۴}�5�_2>��ݾ?�@P�����~��v~>
�4��ZŹ��ER� �I��(&�8SX��$�r��+Ж8���6%u���%iڦ�/v�����5�����*��, �V�%t�R��UU�jR8N���B}h4��}��ta�I��]��C���(9�LJ�Z/?��u�����r�	p5W��v���k4�����8 p�/$Y/	\ P�;��LiD�sYq᪳����B.�[y���,s`�2'W�D� �tc��ӄr��Ѭ��!۳�Ι��6����ٶ���� js�s��5�j�.���Y��Ck�'�4;r�HY��Lx���kR.�*ka	d��Ɋ����k�+��o�)O���{��� �K�4�'�uf�|֊,[�ȨL�/;l��E���4h�Z���t��,A=�E�g��;�Q�y��*`(���Xƞ���uC�HZ�V�-�	�dRW=��;�w�ANj'VI�����K3�>ml��nw��e���sڦmڦmھ6��U7�Q�G�]����{{+��x��B��a�!(:����0�� ���$�5�¬!�S�a�v�՛��~-I��h<��d�HҬA��V�5�]��:�Z�?' 
�IH�[G��p ��� �qq��#�:"aL�w�����zc���I�$K�9�m���:�"P5-���yJW1���q����}�v>�z�VcD�������C��ĕ+-�?�я2��e�v�������+)<d�o}�160����Rh�Ɇ�ï7=��Vp�Aj�)UP4
PJ�>��suE�,�0����0�zj�p���������O<�Ε�U~/��wp+Z �~�'��v��zю&��� hϟ?��4K �
�f�y��F��P0���Y�����6��`�=�������^�VnV�6� � �gZ,�9�g�2��ymɺ����|��������mڦmڦm�^�T8���1+ ��m��[���V�ٺvm������U����lnn�����q���Xcn�+�1���ϡ�ҵL3@8x��,�뙹��/��k}�aMe$��+�&,i���'(^^�_K}�y��Y_%��+@��p9v�^#�_F�W��ޛ��z4�wg��,����K�
	G��((+��8.�2���vv����@����%0-�b���/ԍ����ڤ�r�r��d�CyYS4+�9�^X�w��:�D�2�|�R�^[3�c�mڦmڦmڦm�^�V|���}�<����$g��V���G��%�c��I�a��*�@:� l(����Kc�&K!�`��{gsWېs��8�(�@` 1a�aa]�0)�	�@��U%�PD���TCp- pV�`LJ?��Ja��"E)��t�'O��'��R��oy����x�ݽ=���3'�L ΁�-��iѿ�k�Z�N<��[i�V��S��-.�(ٺ����Y?xZ�\ ��i ����I���S�H5ʮF�F��h4:�jՓ`ZNxڦmڦmڦm�n@;r�p������ՠ[���EA���!R/�'�T���W���k sx�9�V��-�0gF��X3)��vK:�j�2���ag�T�)�$5H�q�9k|��yի_m����C�7�3�`R�������۝�&�K v�S>q�����5��λ^��i�z������4WT,��y����FvPo�����z;�%��P�IM�P��l����^w_*���������:�5s��id�gΞ�gn�ńdU�;E��z��^3m�6m�6m�6m�vZ�ߍ�q�r��q���3����C��7QP����iϰ�W=�3 ��5I3
�/�+%�A%Ș��:ۢ1�A�_So)� F�U<03mT�t�V��6����a+�	�mY7;4�N�\�x�)�9=�W�q����DD��\���e�˄;��Ue�F�in��V~��q��A(�xt��"6d]d�c�:�0�뵬?e�vg4��Ur�F� Kf/�a���p�g�&x(�?g���ft�1�}k#��Ԓ��<�B ���c�w~�w2TT������(�C�gnx�޴M۴M۴M۴��l�F#��fan�m\�
��m��,vqa��wQU����"C���l.]��U�\c�E�<�a��`u:���/'jI$<1��B�!��VM��c]a_�"��1 $�U��:�&�8��zmlVʢ�w�e�3�A�l,�� j��
Y��V�̄��^:�p?�_Pp��´Z3�zb�����3�N�@!��^��4��KK1�d6��KQP�xx�a�)�������c���`GG�X��^��9��)��P<���滿�{���
�q�
?������o8⟶i��i��i���m8k����<��"�v	{[�^��VWW��_��+9����0/���20Mg��1Ph8��`6���J���[���'����\a�e�G `G���?c���Wo�W-�r�}��<��7W �*oq�YH��Z����2��f���d����E�y�9�~�����%p��'�z
E:p�ؼ�+������ݯoxB�c׺ɬ���8�qݍ�#������������g>��;��;���/�������of-����1}o�ߝ�i��i��i�����^j5[�oo�DR��~׭��;;�%�y�Qs��q����j��a�ᔪ���yU�(mE��V�o�E�,��T�ջ��2�CA*ə�M|�߭��5��P�Kx;.F"��	5EPD}��ad4+���*�*�N���\ ?x��/]6���O���~��x`�;���������=#��j����Z1?��?nG�8|)����V\��"T���A�!�q�hL}����q��� ]�x6<�2ommE���������r��?�Q�]����f#�zx�mڦmڦmڦ�4�a�ު]���%��{=�v� �6Sڭᗛ��������[o��<�ȣ��;�2��>dN����~��桇6�[�,www͡��r�|�<˼׵�$�PU|il�Ĭ/}]U_�&�F��L* ��m�\b����J�}��e�H�"|9�R8��L�%��@�:#z���w��W|�����{}�s!�,5�����h����Be8N�ݲ=���ަ~^YyI�/�FQ���$��A?�D�ԙ��"2�.]�dn>y�Y?�n���Xn��6xp����d�������W�q�=���ɡ�`�����}�#?�#�fڦmڦmڦmڦ�ElQN��������7~��̩ӷ�q����>ko��Ns��%s�=�`Ł׼�5�1�|yì>D�������ҧ�~ƈ�C�^՜=���d������h�=���M�r����(,�@T)FzN.˿��x��^���9_������	`A�P��J5��nW|:��h�^툽���]���~����e\�2ʋ��M޼z��@���6 kp�����8�z~~�����7&�����8�F�1�F������?f.L������Q�� T+�e �]q�������������.�?��ٯ���"zoynn�7{��������i��i��i��i{[�v�e�QT��3�щf&l��4s��?�v3�0o��n�B�C�~������l���w@@����0�6���{˙[,"yҬ\��0R8�sЦ 3g%�;���.{�����	J�E�7
"�B��,//���Cfkk�A���q��V���Ѣ�V�[�n乺�`�^k@ �Ԩf������������+��#�T^����"�H@�t���pr]-��t�.�ƣ]��ŋ���\��a7��d��w)=Y��Y� g�z�x�	���d,rgbp�,;��q�b_�������A�ַ�5��w�L�G�QLV���o��_���y��߾9�䝶i��i��i���e�4#���.�3���/��G���UfgQ4K��By
�՟�V�=�o|���É�'�'>�I��3g���>Ips��&K�ɃI���B��eު,��D��J|�a bz^e��V���HS�]��.���P<�"����D��{�C�>���R���;z�$�=�,V@ w0L�����.�Q����C��0��Ȥ�c3���l�%Yz�̙����ho{�ۀ�?�ۿ�o?5j���?����e�}Q�Ui�~�Ϯ�[N��j�I� 8����"H���o������T��w�ü���ݠ��g�~�Ի������uu
z�mڦmڦmڦ��hY�Y�'�h<�!�z��F������-��̃~��梦�7��>VC'c����?~����_ ������g��z�����g��0��X�m��ƃI�"��<}tO �<�ʫWg�Z��t��Xa�˅q�czXkskSj#�^�l�k�����4�{�ሿ/5 +@/J#2�������X"*��vw�\/.̳Q�vh������fL#��:���p�G�`g��6[u��//�d�+��ԙ[~������Ǘ۽ �[�9����`;M��v��t���3�td����x�	3ә1�k���ORG��pk�
�E�N~�{�c���������y��3k��^����O��/���;��$�K�K����hwvv Ob����΀������h\�/fg��a�o�����ϱy�n�������J��u��N��o�w
��������^������}�_P�vw7��d�u��Ís@�^�O>VL���h_��V�=�m��������t�	l��Y��~��S8�jfLo㪸t ^GYh:���z�U9w�>*���>O��E��{��0[��K��iѵ��z����њ�a�9�����hHj��ꅼ^/�z����r�2_���Ö�����2Q��y��KE�y��w��sh�;��bo��E'��܎�������U<���r��^Z���"��[�������yΙŭ�/noO�s��%��^��i��kw�w�q���/4�qo�<�y�7��͋����>�h��ާ6�����/h�E�]\=���Η;'�W����`�g!�����-o����w+�qڦmھLK�6�666�G>�s��haq���O?m����o�&� \xi���������k�N���g�⅋���#�i>���ʹ�s��Es��1�i�>/� ��@C�^ XN&&�t��{0�K����+ڰOnom�1�-u|� �k��s{}u4`5���gt�R}.g@�k�1�x�m:�U�7�Q��D@:�Cf������C���
>�ŋ���������zO�T���"��}��������F�c�kA�'�lX謧�z�+o��EI��������Ц�A�����$�x�+^�������W�^�i������������t��/��/�_IGľ�]���v�뗂��[���������ǵ0L�͠�|���׋t�i����<Ӯ�� m,̴¼��84����1d�Q�b�g�� �3�f��:2v�AZD�*���=��� z�~�zH����d4v���|a}�Y�n���M0��lgm1HF}�3��[[��"&qmi�QO�Im.k���PM�0��64��$M��Y/�"qE֠��k�G�h�X5�9$�FY��i-���!B:�a�h�l��(�p?���z����[2��۬����A��2�2d�f͠�����Z��}���m���`�G�fv;��㒃�m�5�$ٲ4��^o�7�)�-�&����'����3W���Dt���bqa!�wM��8L�4c#��(�<��	}�F�a������\�������KÂΗ��+���lw�b���Wy-�>,�tدS_���y\U��O�-ƃ�1Y"E�0Ɲgɂ�6W�Q�4�,��F����$��|�
I��.���$B��<�Ie(@��0}˟��x0�G�Vkv|����-�[��(g��|8���|6恭����`� CӞ:�������Ռ3��|��t?��1��i2�h85�[a��H��cu�l,�������|�
m�,��5����0]R���K�gR��V!-u[�[B@3yȖu.rA���l�(4p㽝K�G����R�4����3�]2�ji��(��]A�R����-�{���b3�$�t^��@7��F��:om�Cyuz��hp�,����c�^�qR��i��sp�`C���U�M�&޵��p?��S���O�?���`<l)蚨�AP���B�6nϴ�Ao��?�I^�~ż>f���i�]
��4�\�d�cW��9ͅ�����&��&��wRG/Ҙ
��"�\� ���h�c$�$G"���m;�R�2?��r�����:��r\��y�Pk�X������/sIÁ�@h�D�+�Zq��	�V�|J�����p�4��"*"����z����ѧ�s>�9ײpdsפ��
�F��>��A�_4�u�)?��f�h�w���v133��bic� ��yc�����"3m/I��6 ��7�԰��K���ѥ����ի�����x钹��/g��ɓ'���ڥ˗�˿��8Y�}�ɧ�ͧOq��׳�s��8�/#\}��ߥuE��)��M\SE`��+J�6�Af��^ڪ�n������V�_����S �I2.ύ�`�E!<�g�>���׾����r��ss�K��v���m�ms�lҿs�q��̧���y�����K�^����d�4{6%.M"�HK ������{�=�gΜaj���a���o6k��L��v�xx�� w:x�<�N�!�뮻:��w_�~����g���^�|��-�?���F�b�V�!�`�Ή͙:����BN��I���w��Gx���)���Υ��=������3��:�F�6�$�6dK�Iy�i�KA��O�1�@n(^k����6>C��8��[I�� ��cIdU�{���l���k��$����^pv�a�:	 26 )e�~-��I4�9�n��I�-����_��A�pyD:ρo�����W�`�ࡢEa�&��������������v��V��,~b��:�/�N+`с�4�3�����軝]!��wlv{�{7-B����� �D�?����D�A����KKK������8���EP*�$����s繿ѧ��K�'�=6]<[�M�h�~�|n;X�gX�9����С���@��
�^J�!!*p�,^�E�������p}�v�?�Cc���z��
��A]�����y�=S0$�ȩظ.� ��;��˚��紌!ԝO1������u�Ι�./?���s��S>�XQ 3
EK2�}D����,�E�R�ف����#��z�c\3�(�ņQH6	�t����v!C�!VW XR��*�^���H�	�UƮU�o%!��w"�Kx����M�;��>�V���q����=��{��Z����0�����>^��P�%�@=nX}���� O���N&�X�0n$4�ҧ9z'�ЗQE:�E6b���v||�k?��%�^�cر�h!���qGh*G.���2n�Xs��A�K�z��f�̍���,a�a[l�X{�����H���"�_��L��I�R�8?�!���.L)ػY��;�Lc�*�<Ip�YlȺ����lX$6��p�$�l��c���8��5���`��]�A<�o�F�x��yt0ۉF��}*�Ρs�#:�����A�5%�!�Q��g4TpIl0�������"��MC&�U�y�`Ȱm��K�l���4y�mlt
Z{Du��JCX?���;��$��E<'�kfgyo:{����?Kkl�5g��C��z�!�O���������sV1���rv}�{<}��we��jf�}����H��M���礼F^��*p��ʹ&^��oz ������+#<e�a~����e�?��.���u�����7 iMxь{,>{����#��-��{�W�~����o>��Su�#�/�]Y9�I �>���ُ�<m64c $�ر!��k��O��y�7��^?��8`I�Q�a��e����.�!4�|���c�XDǏh�^\YY�{aq�n��|� -��nw��A�-�'jHN�y@���M:�k�jt�N�1O<:��Š�7���s�a��������F��; P�z�I
@Ӱ�� � �0�p�Cyk�3	��?�+&,��L�΅�gee��'�X�>��>y�$@�
���@�gP�@ ���W|����Bf$���2�Zw4!-��y 7	$�t"4&��è�,R�w��'C�~��b�v}�0WUYX�S�N������<ȶ�2s�,a�
x*a�Є1M�l���NCGZ�@ߣ~fapȝ`cv�'��~��C����q%D#��
��� �j�s�^<��~�s��ˆ
�o3�����<O9��
��
``(d�;��k��܏�V�y諘� :�I� !��@����HYF G�%B�5q��G������xt��y�-Ƌd�f_k��X���ɞ���Ɵ��s�8kXN^�}��Zr_U�QMn��13-IƮx�C������M(��F �Ȁ����.5�5A���!B���윜�Z��\�!�I��}��?@�|m#VP���c�6+e@�Z�� ˎw��<Ɇ.�x}9�ת��2S��n�28B�1����u��0�� 0TbN
a(����uG ����^���/F_b.��B�T�r�x�����I��(��U@3r�)V��D�C���H-{�`
��"5f�$c[�n�����@�0?�G��r�$�8����7��| ���c#O >ݧe�Y�2�)�TΊbS��?K#}$s�ף<�S�z�^��z͑����5���;x�# YA���a"ศ�E+%=
2��B2v��h@ڤa��qV�XV�l7�g;�GA/�h�؏~Ϧ&����7�����EA����ԏ[u2�>k��x�[��Gt1Yܳ�6�t4/�o����<�;�w������]���n�^K�`77�9P�ɘ��{���ٳ�>]�z�����H@;rD���?�c�c|ƍ�@�s��ڤ,���}(�T;SO-�:�/7&��M�qTUR���6�և\���j&���<�+�ت�X)r,N�G�-ɯ�<�!�׉�4�Z�] ZM��sϞ�O<���]Z� vaXb�.��
J�����8f�o=~�Xc}}��Mi,ߘ���7��0.������i&�%�qZ�"�Q�i� (Y��_��כ7��������'>i^����[&�`�7lԨ~��'�@K�@�ho�q�wZ�JZ���<����(j�4�����Z�bW����x8�mr4 ٓ�Ѐ���bp�+��4�
b��O?�#��l52�I�/�\U�@�%H^�vw�|�x�����.o\f�,D�l˱2��!  ,�R��ǃ�6X�^[��f��|_�`{05�w:l^ j��ƕ���x�с��x�f�yx�|���7�Z,U[�r�p��=*�y��Zl� ���޴��ҭ���4��5`BC��@߁7
�Bǰ��3��Zx�A�{�H���4aPXCA� q� �N�� B=Z
0�k��W�Qo7�	_MP2���ߘ�z��ClL�s�8�x&X��'aM��Z�Fϋ���,��zb��W3�pX�^w���M��H�x�방J��ȏ�L��% ���G#X�7�	�ɆC��F��k=}A��ê�彼�P��_k�Ðs�ʐ�)������B
Ð_�5W�1�3A����s���/#>Y���To�c�)�E�az�(�<oU\��R�G�aFɲ.�3KZ�q�uB��-���p���ƞ����� �:k\*�q���|������@]������E�Șlh�!�?B�Ք�J����1ck����иM`��Ӌ������g}R�<�&8�r{��a�����Y?��5i.hߋ�RCFrؓ�O:�=�5`	�{ų��Ղ#PG2�\�7����C_k�8퇎D�I�9j� p�g�s�&q��EF�D7�)�v��X'5Z��Ԏ��1����� �����F�����(�8�zX���#��Gq0�PuT��x��1��*f�D@������_�)JV�%���8d�kd�ө ֋� ��̎�#^oi�,.-Z�*���egI�ތx����>�{t����6�9��w��|��YJ�)D�`t�!�L[G
�޸Qo��ɸ�b0��q�>�j1��=8.M��w�٘V��mJ�	9���VhTErUb�Z::=MZ[$�-�4	 ����w� y�3m�^m�u�mxi	��(��}��q�'�In^�d�~7m~߸��K��u �5޿���$��!��U�<���� �mgn3W6�r���ŋ2�i<#B�v�PyO�w`P�92?6y��+Q4o0J_`U��5��>``�j�#���g�t�~까cꭅ�������LQ�<l����}z��	c��GX�(��HU]ȗẰ�<K�����#�nnn43�i\�|�s��̍n/���Yh�{�����4�gi�@�9rđ�d|�A^�������
���ln��6vnx��3������B�xq�!6�~��^?b�# ̅F �(a�#c��ᖧ�J�V�>����Kvd�a@�99وxP���,Z\\b�&!c�lA��޽q�m���k��l,p��{{2��m: ���z� B��]�x�ݼ������� �9"�@��_zW�yx�`�U/��~`�!�f�n�l�t
�	�QO&�N�Ä	�ǧ\<�ܕ���a1PBHQ��B¿	_�xO��>mBBQ�˔���{��K�6�{{6)|G3Y� �ց�x_(9G-K� ���Y.i����7��A2���1�7���+�?�G`��0���X� &A�~�sQ0
@�F��͚=@�!�y�o\k�h�{��!r>�W6�r.��פm8�/�p���GáU{�&�,�F1Z�#���+Eס�RZ��?� �zo�W�&���=K�����t�\��	�W��x��d��9�)��?3��p=�dM��ܩw�@�>���>Y[�9�E	>s��n��AC�'8���E
d�Z���:'����C�xpX�=x�x�1j��'p���@|�1kdf��gãBk��]��~�0�}+�^(J ����2�z�qǳ<���"��r�aʚ7p�� �X�}�=���v�: U5݄�[��O�+U�5ӑ����y0�	8Z	������5?�4,\3��ǥU1��<�l�����U��k}> ������_^�+^�!���꽩��k�衆��8��gI��Ep˱��蜥~���1� ]"vBݡ�v�9��H*Ŧ��Q�D�z_M��q�s����BV�5�#f��}���|�DP��j+�Vi�������P�8r#³~�I4C�����؇��]�s�2ٺ}I ce�^9Fd�Q�N�eH�h�E`�u6Lx����.�"�X�9l�y�is�@��#G���,��+tz�J��"oQ�A�}��L��b��Q��t���me-�2�4��P�Pl����[[Li �	�*�ߣ����xʹ��r�z~�ە��hT��!`�3��}>u�����c��s�Xlx8�1�}ǜ�_���Ml�--.�940�~��U�����������'wx���p�܇i�|�����ٞ>}�}�s����Ϙ��1?񶷙������ʯ����|��쮗�c7�P,�P;rԬ,����M�l{g'"K:�B�A�٤ͮ���g, ,��st���e���C�[Q��������:���V�わf�)��R�J�8��&�� Ā�Z��n*�N������)_�D��M�=R}8��^�!{�ěpd�p	�T ��'T�}�C�9���u�U��N�8��U�=�0@�Z|���CP���N��
�AA�C��Ӽ�c1@bX<x>mx�=o	��>�G@��i�\q��
0����<�lL�YP�+6"zQ�e����1'�~��/���+��fv~�&�"�% S��5�]#�S��s6X�K��x�I6V˝��xh?ʑ���=� T�YZr�b�x��\-��C�ǧ�TDe�5�[� 5�DF�|��T-=�������)�}M�!����k���2J}X��y�EZ<���RYH�A�Cך=�`ת����yO�P%*\N~�;jlc���-R# ��f�N0���Q��r������1`� ��t��}���Q�W>������O��}(�B��N�Ay�j�gؠ#����Q>���3q�QH@&Vk_�;|F �$t�8D2�`Pσ���X��6rm{zf0�aXc���K�~�^/���ue�5R�)I�x~�~]ӱ�g�(��3�^0"u�$j��x��Oq�1��%���3�R�F�g�x~�D���7��� '��B�
=/���4�&�r]�����k��+��S�Z���1��` �b�3�C����W��=��7D�E {�#Xs�{c�-�(�xZ�^1�ZFف���X��l�C��QF�Ұ�x����n�Aǘ/��"#�Gu����Tg��k��<�k7��α�s)��}����0Y���JTC�kV��!���vK��З�%�9?F|B/�K=��2(G�3�\��NO`�>�è�v�v$^��5/^Hh>А�h�y��yL>�䓼?��n?��Cf<�X�;z���'>��-H|%Ɍ�����u,-��s�8��(�	�xM����7���0���.�	0�����x���uLuΔ%�%�!k�_�5AN4���Kd8It{
8B�����w�����55Z��1���M?��^��E��l��ߋN�rj���3<������S�z�/��i��uҿ����4_g�Po��wޚ\��?�أ�����Dw��e�m��'N0�����s����`���Ǐ=�E8:q�x���\c�@-�À�{.'l������̌�8D��3i:���@�
k>6�Q�U#�r��<b�-����}]A_X]o �����]A�Q��L����3JdC���%`�Ԍȇ�q|,���<���p�jL��z:*��S�	�����҆0��a�e��z�>{�Փ���+x\}2Ρ?u�d�k���IڃWB7,L�[[	<���/' ׬�E�sQ��*/��Uk��3Α eY����?ހ�My�F?a���3�{�~��Q�[�L�%VpB�I����C8Tiy��A�y�Q:���r֠���ە���q�{�MC�U�n@,ZJ�*�Aiz# �H~Sn`y|6i1�Ǎ�c5��`I�k�O!Fx���X<��x��%�����&���_/2��)H#4��Ŵ�o�7[oXӚ��%W�t�x壟|l�:�7�}��h��f��Q��_���3l�G�N�Z�|�fʹ/�&�h2SDt��$I�C�m�!�=X�VW+��C�����B�� �
��1��o<Vh��b�]^�z?��s^����C����{�����Hx�<Z3-�v4�������Y�}>��Ng��[�D;�D!3�0Wz���*��x�E�En����p�
��1���Ft�(�K�z��y�k4�����՜	MRE�9�jV�4�9jk��.�D\Y�؋�Q�����ku���dQ���/�*	˨C�F�Q���eJ.�+je�dh�1����(%Ʊ(WtJ����j���N��砋�{O(-��b����5Y���f��G�L�Oi��lfy.��zG�א�Z�U;b�W_� <!r~�⳸V|7�E�@��Z��R#�hA��$�ܿRh}���F�R� .��!u� �9];�?{�9�#ĝΌ�P�Y���@a%uc���,����>�����A��p)��d����j$��K<p܃$��xԗO���E��(%�d�1m&ί�T6�[B���ɹO��}J��x�D�c�̻�}�<D�80���i�w��R�����}��5�T*�;���>t�Y^Ye��N�ZpXw��ř�_~�ˍ�v~m^�y�f��������&�yZ~���f��f7�n�����1���� ���^�:������sL���p�<�i1�v��1CG�)'����Mu3d/2�"�V�n|m��c�k�
 h����:4,�h��W7/����?��c㳊��4a�ƛ�,�)���)���ɒ��\����1Ǘ���7*H�����@M<)��K��� ��}���I�+�EiJ�П�L>������.�[*�L2���J�j��� ����'�N��s(h�ϋ��RfjF�^��5��ϊ���U��hD��R>,�UA�$�L6'L\�D���$�XǇ&n)�C��Ӿ�kF���@��#G��������c�?��$�u�|�O��=�z�)&��¸pc��/j��L����:�X�9����[q�V�A5�X��(��+������c^��p�Gd��g��|���l򘇡H�
�\���e>�`��~U�㓓g�<�}��ϱQ�X�s���B�����D�C���?U��q�י
Aߟ������g�G`�ycO����^��>,��<�ћ���+��B��y�LE�[][+6�I?Z>�F;rO�H�V�Xc��U%�V�(�R~V�������L���]3�؀R�q��,�7 tS^~�Z�B����T�u�u|��\S
S�^x���f�{�J��1��G^��.9	?���:��֘G�+��tL�8f�	���~�<k<���%�����\�� ��Ɛ�[���N����t�@_I?����O$�!�T��>7��9��N�0qXS�����5�?�cpm	Q�5 1���?/U�i��$WxjH%��ΧhB1�O�e�_gf��*L�����h���N|�-��i���n��SH"�dnѳ���Xx���G�!@˞[�̧�/H}�-G-DՄQa��uV���'ޓp,�ه��D:�G�r]+�a�%���Ս`�)`x�só���%?�=�D������B84%���&�����#!n�؆sB I�5�)EM�J �ɧ�6ozӷ�X�؂:����������j���S7���:�g��C��xѨ��o�/����������������Nh�,�DQ� �C�ڼ��bc�����m�ݦ`2Z�����o>��d��9!Yլ�Z�^	�ҁ���x�W��j*�P���E���ˇ˞�
 �b��h�X6Sސ� -����w �� b�a��|�[��*i���h�A�y˽/.�����bZZ�h�縩gS75I\�L6�yo{�ht]^.(�_�ԛ��`�Ӊ�g�D���
{�G�r��f��M�?��[|\��h�ե���5�\�g�,����V7�j�_(i	J�����`<�*��SS���]d�P�00"�]�*�k	u�O�k��E%��E��@�s0�0�k>k}��	7h;;ԫ6���{:q�w��5��\��A?a�`!.AwMh]r�m60����f�Ú���iҕ���X�[�/	oT�虋�g1	�M�!D�̈U'Z���8d��D�]�i�&�2ܻR=0�E�r���d�~P��c���������14J�$,7ә+���1L�3<�S�l�}�P����:?G���\k�w˝�HOǉ���x�l�<�crf���!���S�kb$���ض}x�(ý��f�����))ʓ��f��Z5d��H>c<���������U��YC�r�	�-Y۴�uz��'B��iUri�s��K2�����ӥ&;�^u��á�|1�R��8C�u	kV�g^�N(�`�kQ/���ѵ��^�+��p�tY��d��m�$S�+��j�hc���ń�5'amo��8˫+޸_+4�ǥqt��i��j�,GI����*�P�-}�<�d�>����^K��e?�g�QE���Â0(��wN 2��P���?�Ix�e�ܧ��z�=�Ja���P��S��Z��^���>�{�4�����dRjX<��tF�sS�0�,󟛌cyv�S������92 z��]�rT���:I�V(Fܐ��fJg��t,���G�N9K�n��%�B�9�P�=Ĩ���c/��;�=����{^A{�.+2��;;7�����5�NϮ��O14ni՛7T���^�@�B<���l-����~��+� ��>/%w�ڕ�:���׮]�P3P�mR��B�N�&����3�������ҍ#N��.9��L=092�
�e){#6���۶����>\��5QB�a8��������ذs��%`��\V����E7dp�^$� h*�~}�����$�P�fݣ�1��a"ϫ�P����#�aJ�P"�����.XlPJ�蠖�(�E��e�3I �>dY�$����W��zPԋ��|i(�������6r<�8�"V��	��'�{�Ƀ�r,��OgE����5�ᩱ7�
����.�5�+�Ǉ��-��8 ��4��sĸ�|yC�l�!����:�=�<~��9w�\Y��p�"��{�5����x�D��-B%�K$�ʍ�z���`C=�:��ӈ��1\Y�
�]7_�!��瓟מ;Ϟk=�
����������צ>Ήs��Qy:�5���9�1cR�'�\�R~O�O�����B�Rt���7\q��.���<�xi��+ր7�1����))�O�i���av��5G.W�7�0�����oJɸ_�/+:x�~��$)P7Q��0�)��1����t��f����s��.4}��*�iJ���dMd��dK�>���R�jH�r]�� Y5|�Z����s�9j��a��E~=P��2}:�4�M@��$HM��1�&,U�ᵮ�-W:�C<n5Z�k��T���gS�o���k>��J�$���Gc�V�ʋ|��I��a��s,�h�Q�z)15��Z���1X1��4J���G�2���
O�icO�K� B�8����9
�u}WN���(�DS��Tv�:@upy�4��J�W/v�@R���/�A�i�N<��_w�d"j���l�v��DI�݀�_ĪB����9��*7V%>�nE�xK�40���f2��B��D��Ct��S�?v�8�s��^�� ��D�^���-�� �~>�خ _�6�7������a�� ���G>⣉M^�M ��=�_�`9$���I���k���.ƧN�4���KV�|1�������n���{�{ݸ���t��M7�Po�gghb��Ď��2O����X���$3�\��Δ�#���ox�Y���;l`���|��&u���,<*:���3b�0�ϳ~��\�!��'|����6Nd|���u��o�t�K �7���A�~����'b������*�׷j���\,��� �I�@��b"���<�Ǽ����-@	7�u�^�t�����k�b��Ϟ=Ǜ�t[�,,,��e'PjX�3& 
��>sXݘLh�pے'ڨM��h���`���ƘH �d< +���>��~�S�2�~��͓O>���M����`b��c�F���~��864��) �b� _��� T�}���7g%�q{���뮻�k���.�5�q��O0�����X$J������@�Te��TYU�� 偉'�i�D�*?R7=���������_zȱ0"ԅ^����fD��c��c�Y+H�5+��gq���g��W��|�3�0�FF���E�y��]f�O��>���rB胛����R���z�M� ׀cb\����csC�I�x�T�t��I����xV�*�}5ք'�������/��"��I4��Q
U�P�����@�ȅ�����N��Q��Z�
&{�=�I��jx*�Q���J��MT���R�f�D2�W��0>�9U���AW�7H��h�?/��pDΕQ0�G�S^UH)�:X��,�j��I���j s�>ӨIDA�gB�R�ҫ���k��Aׁ*����^uQ�)�3��y�_�}��P�I8 Y9`q�4��?q2�kyY4G�����&�Z��~��&�iu�PiTT0K��ͽ���س
-J3�=D�ulk���&��L�Y"QՄT��1	�S+�Q��Ј�zu��[�~B5 �j51`����o����W�L������NB3j �'ޟa����զ���"M�D0P���;����8��.�%1D�2��=#
����sV^��g<������/�Y��a��C@�셽'�(ϩ9?L� p����QN���?���E�O������߿�?��7���Kx�p�����@��_P'�H��o�W_���Z�z�
���Y�/\�����9G$?ilL�O�&����^���������u�0�{��8L�_�1��p8Tﳀ��6EGT+$t�Kle�p#��x�`� ě�J���������ڻ�`K����}۽/�6sf�H3#����1`;T*��+q9e��xpbʮJ�R~�S�J"�S�cRv9T��<$�)I�Jv\+8�.$@�F3Bs=��w���Y��Z�ϞAرAF^�~TS3:�}�������_6I���{��F�(s&���a��8���0���a+l���۱ٞ��> 6��{b��n�歛Y&Yi��QV�s+J�������]�^���V|o��n���T(�HY����w18�f5�����H���B�M	u���B��+.:w�j�a�&qYE��vP	��=��(,��7L�񫻩W�.Ӎ��@��O��O�'q�z�u|�FO�es	�X7�9i0����A%\ڌ�����P��o�-H�X�]�+	�NQ����׾��/�(qQ|��P�CRzO=��=�X����Q�c���ey�m��}�x�Q��H�h�A�[��q���N��ޕ�¥:=.��l���}*|j��I��������r�d�4���b5��kW�^��y��V�U�ǟ��!D�6�szm㈼ʫ���D�Wx��%n��8��mc:�(d���_���q�msz}b]r�/�#��������o�@��P����'��N¤P��D���Q�8���_ۚ���Jʰ8��Q�`�?;Au�q����a�/D�>��(k|�zo�������^�j�����9�5R��5Ρ�"|f<cȉ=l���mD?�Bw��".��18��:�~w��W��ܨ�����'.����Ha�k��	��A^Y��Ik,�ҮD#s�b1t'�)��� ��0���y��hn���u|�lp��Շ	ҧW���Y����~�ɔ�՘�m��>�醚v?a�&aZ���~̶�1HǳQ8a�.=����.�ק�d���=�'�q��:����8��w|��iK�xf�7,(3	5��o�b���+<Q׵v�S��,L��,�!��X�fl7hϡ��B�M����~X�ھo��|��]A	Wa�N,g�0�����﫧�B�,~u��
��ڏ�*@�}�>U?'�Nm4uj������7�_�,��,�������C��i��/���KBs{��YX�9e1�����+��>����h��6��>��o]���	y���[������W�_X���8�U�B��o��o������E;�������v;��#o|xr||R]}�Z�w��=��#v&G7�b_�v-,p3{�ʷ��%b;o�!T0�x�'�&?ѭ����M��ߋg���$��V�M$N4�a��͉by���#:���pIW;��$�+��w]V���έ۾,!�f�w��f�k~�i4�U�6R>����?S�#E~2@�[���8
����&�u�|�c�'
q������ڵ�����O���Ʊ^2^Ҋ��C��?�}��&�(pi$*��h���0��u�.����t�)N��t[z�*S�k��/�W���v	ͷZ��م�f���;����U�����kqYbݯՈ�ѹX��Y�`#�a������̿��/���)����$�K�V��m�a�G��Jxz�1��ѳ8j����s'�m���;��f�F����\u�1��筧t�K6�c���I}�׊�NP��jT&~_�P{z��x������QJ}_'
���Y�'�'^j$^:�����#n��)GC�X��B���z������kmW�J?�~�V!j�l�ĭ�Iۗ­�����uЕ	_�1^s��rt��~L�5� �I|�[��QX^;�6��a��Q�8���*�T���g��/��q�7��h���w|�t�_��Wm��VWr����~\����
U�K�ǺY=��J�\���|A�m+�YP�?^jå߻�Ą�C,X�ϧ���KM\�;n�qR��3�S��׿���	�^�0�2^�������,��k��ɨ���6'��	A[�$E+�Q(����]�D�ޚ��:SmwC����N�Õ_?� �K�
&:A����:)��{�	����}����NmUѹ����k��ܷ�������&��F8I��궟�����g�e�����o���Va4�*|m�V���߾���K�H��⹍�V6jj�5;GvuQ?��e5��ˍ��Q��+���_�v9~>Զ[��>��_>{��đa����o#���J�J??gik	�٧?�i�9�֚s�z�q4^����H���Di)M�k/~{舢��W5�����?I���p�|��qYg?���J�]��?��٧��Ӷ/}�+_����C V)���}�{~[�Iq��}�o|���c�=Z��G������k������(<����}�Cϲ�M�|�۸��ov;��x��Kn��v.5�.nܼ٩�W�0��g��;l�èH�T�pcQ{�:��㊣(~���/����T�ee�8���K���j� ���Ku:��;���D��h����m�`�	_����F؁i'/čtZ���:��%B�lv�uџ̓@�W�]l5S����~��jQ9\>�߷��!�fd����HΨ�AO�.�Q:�OU8��L��񠬃�nK�~��^7L����G>��=���
q�u��ӈk���;aM�����G?��ȪɊ#)�Y��`CMX���C<p�v��%�z�N$�c�Y��б"�-���]uP?�p���&�EK�Xbhю-�%���A9v���+����򸽈B`�ֿ�����˄�g%��������Q?�+^���}�k�����'�~U<t�n��)������so'�s�:k����/�(�������]W(�}��k��H�^/���>�w<Q�s����r�F�%v�3��t���~7Lڌۛu/	�~/�hœX=7�S�{���[Q���_�x�������p�>>�8�_�xrq��G����:��Y�"g��1�m-�7�vs��i�镝X��T������5��2���.�dJ�� �ݷ�J�0u�N"l�B�Ȫj^��V�~����X��pU.�N��+�8���u���f���8��&��_lۧ}�_gmW���ye>���C�z,�?�~͎e(��K�k�FI5w����G�?��e�N���z���s��z�|G�����.��D,m�}��_J2��-\ݸq�����:k���[��	F7�~��/?�;�}��7����|O�n[�����0�\�K�}/~M�C�O����ZP�銭x�3�;�3b��xB`'����u�d�	�~���tl�����#����o�ۇϮ���Z���m���-���(\a��sm��F?������>c}v�Ä��H'V�Gw�u���J���Ս����apeN�t;�o�d�����^�GO��a��N��_��N���|W��� �9�>|?�K"��ŉ�z��O{����{��瞳<��.�T
��zx�K��l7��W���X��O�a��7<���#�l����R�4|7�����=ӳ�	~����GݎlV懻�z��u��{g�κ���_pgT=��oy��߾�Π�n��v;��ѱɰ~��`��A�ѥ�tR���Ck�X��3����3���+���bH�*���āp	�VG5bV���Iq�-J| �NM�a�/�]8�*����~)?��
���(�}=��=j���X����tg�����C�o��\<��ã�"�ek#�Z
�7��y��%�FY�vq<sWA�0��wa�ð���~k�
5���QH� �}tae�*�[�!.˻�ڹ@T�	|��G*�}MJ��f�5~�KV�?f7���g����X��YvZ�z��O?CK��;:��>d'���<(b��٪U���W��ͅp��mS�������ݦ�k'��o;-����2�-����t���3���tYX�l�^���u@�I�'��뱆 ��|Zo@��e8?0a;�_�m��9�Fu������?s��q=�6�#�q$9�X���_�X�<փ;c��ڡ���=j��Ȩ.���&��x����c���'�|I����5�Ш66^Yp��mxX��/ �;��+Q:Pk�����o{nqd1Qm�z���"����x99��oN����҆Ǥ�s�7n�qW�M[�N�89H��ަx_��V΋0ڼb�S�~���B�����9���W^�e�E��.�s�+8ƓG-媰鶞�?�='���kX���JWشA�^��*�JR�y�C	�ܼ}[�MO�$t		ǉ.|N��3߯=��awY\)��xa�+w��k�����,�j������-d侖U���������9ƓC?9��P£���s��Bk�5`'���_���'���"�����l�����>��1ǽ�O=���o~�y{\���d(�&i��,,�_�eN/�t#�r���1t�p��3g���g�f�:�\�j<�3��XC�f�_�|<�5��~���x���u����l��n��N*�1B-$�ՀuׅQ��N�����awhWW$O���ҥ���8�� �/��
��~~O�Gc5�&��	��Є�xU)t\^e�{�h���b46!�z���%���v�q�6sk ��"�^�ڦCP��������89�������=���g_N���Ν?�}򓟴En�\y���ߺb�ݸm��u�z�۱_a^�F]��{��x����|~�Z���5;Ij���'�=��������?��r�t�ҽp�����rY6��h�h�|UN����b9������[��Mpr|\�xPk�5�������؊�]��S&Tq=��J�.���<�a���$��Ƨbw�f�ee�W}�{�C����ۻ�~^��X�=2����ޯ�v1CK���V��[��_���Sj�ո�i�d�2@�vҭ��K\^���d:�6G�g��j9o���6�����j�엫Q?ZU���{������=0w<��g��s}8g�V�P�»m���]��]������G������g6٥۫�^��#��)��Y���Ёw���u��ns��r�}s�Qȴأ]ޛgC�t����\t�tv��[M��P�z��/�`�ˢ(��:/��֤�Z�ݸ/W���.���fv��
����n��Z��s���sl�~�/:_=�Ka����&{�2�a:�A8���+w7��ڮz�1�ܗ��������{�
�m��e^��^ݷ�Qv�XW�Ct��{�{���O��4u�����d�w�y3r�o�Q˺n_���7���˄
�]_�l1���myy��.�iF�۶��Z�-��c�%i�M�s[�)��ځ�����)�8~�p���\�B]�t���k�{
ݩm�.���ʦ��6��f�U���sҷ�~z��}u[�|e�I�r�6�Rn����D�4�֭���U��8���V�
�%ZN�\��ں�lӑ���2!�z�N؊�PF�󋹖���2L6�|۳"��"N6s�"�Մi�2T�:!����:��J��þ�SA�t�Hc<8꽉�G�P�џdn+��&;'Y�iX.9�WOV2�\C�+b��w߷�XcYJ<AQPW@��k'���khue�ãN��Xb;�n�����N�4qٿ��R�_~��otZ.z�GӴ�)�E&Vǫ.N�����9�6�P��x�g��#�;��m[�+�,�k�E����Ix��]t�`�p�/��WQ�N����&G٢z��u(�1,
�A��F��<�Y����h����5����2�Ez��߼��m����zrզ��)&��Pc��������v.��cc�>}�ʕ�CYAZp�5��|���mW��1hB����j� ���
��o��久\D�fX��������bw�x�J��uk�廑�uS�S<y8�p��H^|��v5S��:�~��k�yVΕ�?��/�Q�mԵ�Օ�7om�ǉ�9��A�=kߠA+���wV��P��N��>���bv݆]�s��bH}v�J��mđ�XZ{����޻Tq?����~�-}�����N�on\�Q�Y��u�{�*-��>
]]|y�*����3��^Љ�v���t�^���h�X5��W�ޯ�������p��i���}�z|W���~������A#�ָc�O>�����>��ޜ/�W�݃���+��F��.ٿ��_��o�;���b�L�ut�oo����v�۹*�O�2��ڭb����,'Kk�1����n�Xխʹi�0T�O�m��Ա�I��k���}�_w-]�^��o�ѹ�k�7}�[����I����̒;{s7���;8T�Dd�������h|���R�������G��������]�����"�W*��65��K���������;(�y�.��a/i��L�[t�c�Ř����g��#��t_��v�.��q����NW�|T���lk�P�/lDi\�ŉI.�P��'�z����	^�Nd�.����_t���G�ښڨ]>��4���b(}�U�ʝĭW�n�pa����:.��k�~9r[VZ�>�M˾Q���'j��.]QY̗E,;p��N��	�;ؓX����aU�ǵ��YQ����n��c�bY�j�O�����Z�O�����k6�{����ޫ]l�'��R"-u�ޜ���wM
s���׸ڣ� ��wvv�PW�祫C��s!��'���_z.��~2�p���=��ea(��$D�,O�����O�w�"��զ��uA���ɷn��B@/6��ʙ��:�������η��}p�ݢs�>�o-K�M5����RW<�Η�0m��F�����u{�x2�δC)�MDW����=�7�����t�UG��h|zX�dT���bH��]��?������tuz���8<����h�]�!;��,C��pE�}>����@,w��g�TB��c�4_�s|1�Rl�ڇR����U�£�s�����O�։�檌tR�=r}K�q=
W�2�\���N��6��*��	���n%���S'$��7����+a�ɲ��m�K(i���aۉ��"LH/6>���#�����EE�G��<��<X?��ڹYy����v�����Z�?����5	���wf��_Ȟ��3ٿ���NN����ٽ�'��O4��;ww���٫>�~?��ת{��~�z�3 x7~�#����s����t�����.���=�^x���~�7�}�����������Q�r�~����0���==���������r���Q:wy���{�
z��F�:_��!����5��纄��3�&�۲ZW�;$�j�e�rUI��=Q�;�c�]���ծ,4L��
{>.+��]2T�'��k��a���i�B��Jwpw�л�cK�V.���$W�X�}��z�[]����d�k[Ml��\���
�{�;�B��+��t�����$/J��h ZA�DJw@q�w\��P��]�-���Vwi_OQ3`�:ުdF��F�ҥB��:���w�Jg����ۧ�L��#�K�\���� ��
������+�J�'��w����ʍ{�j��G��V��B��=����ۋK��m�y�1b���ྈ��6l=x�E�鎳�7j{;�]�*B��fY��������vqt�ӥ^]
W�רj�y�H�ڧ��x�x_�碑$M��"6�_jԺ���G���iif�V�f����l�����E�ԥR{*�Pē_.��H�a��OG�����+���<􁮺�ٷ��*l��z�G嬃�m㪈sA6�6�m����|~lK��whX$f��b��%o?ү�6?��U�K�|���(p\�&���q��>�k�N�ز�_����݆l��b}��&!�ْՍ_�T��q�3V��(�J�b�����$��ĞĪu�I�-�au��P��+u�%���*�IY��^��
ܾ�&p�a�K�Ha�
ue#������t���m�UO�'n�EuTR3�9��f���m�.�]����¯��j�0��t�pdeV�WX�m�k�s�X�������O��F>,��rN���dT��tqq�̓�w/m#˝_a�Ug����C�{>�����PN�%7n\�>���eozӣ��>�1[����jm���߷]x���+��^A������R�����A����S����~���	���N�>�x��/|!w;����S�Ϗ�����s�C���n�w���[[���x�O�i>��s��A*WP�g��|� �j5ܮF���}誒kex��ܞ�.����&|�`����c�o�������}�`]��Ua�γQQOTR�~��i1,V�z��Tg�ue��p�V�p������d<�pR/�l���Φ#�k��>湝w����Z��.�Rٍ'Ũ�U�ʔ�d\k�߅��p��KK]����G���0��0p�L��²;�k�l�Bh����T�֥򢛸�ȿf�/�� �#-�H�Ze8��ؿna���a4�;�����h��.��z}U�#գ�hv��UY���Q�r����e�.,S���J�p]���H�ޛ���"��ӑ�׶�m�Ӡ���0z�j�Z�=�<�g7ڇ9���+cYHh5���Ia~b�:���F�5�Q�؛��g�C=��6Z�m�FC5ҥ������?9��nv'�����>P�=�����gvm�{<ֈ�&�N�d��Zy�r�� �s���R��Z�.P���.$��F��YgW����Y(Q}�͏9��c'z�v����=����O/ok�͕�V��̴*�,*�k͵�:�(/WK?)�Y����9.���vm�r7�t��W5�U�����3,m���}���;*�aҵ��j�׭T�°/KhZ����	����׼uQR����lXX(U���;�"����FWU�b{Q���~~gw��#[-�J0��:���~�C*E�W��[�I��`gM�+?~y�k���RT�T��*�6?�GV��'��K��g���� �{n�A��o/�dW-NN���#�>��3����Z'�O�:]��|�w~�^���V��<��4��>�����+���F���
~�Bm�,��c�>{�����}��
�͛7��.��}'�>��(T��'yY����'�]��O���F���F�<�����y�k5um���R5E;���ג�������U��u��v��R���^jb+�R
�e��[�B��Ë>w���+{������Ǻ�?�uV��V������
T]�)'e5ҤH�6��f�ە�J�U���ͺ��u�6�r�3˭��;`6���ד���J�^� ƅ6ݗ;@ꅪ��r�kH�R@�{?���!��r<�-gt�`��6���dU�����v=+	���mA_W��
�Z6���v1ua���/TۨI='��b�,l�˼
���^O�`p�L�Z�B�W�%���Z�ki.��T�e�HR��.7�Ye\_,������)
kU�z�[�B�0��9,�k�]��vto|�;ռǉs.�BI�}r���[\���j[��}�ф1?�V�x�!�BW���-�$��;wl�1��j�"I���bxNH��]W�ߋ�=���ua�طe�ʥ��h$�VԴ��:X赳mJ?�����Qͽ�*}ow�����8ʯ�U���F�7�j����0*j���6:���etUN1�Y+��Nq�`���2���g�6t[���okͭ����~Jj�m�X�3v�Ѯ�z���MV�
u񾋎o�=��T5Y�z����DfdԜj�˰*_:����ኇ�C�'���'�d/|{�/����2�*���0ʝYK6��2�v�����U����ݣ����v��:. 3L��	m7z�vw����fy���m+X~��+'�&����6l�m�阌g��sV\�t)�x�~-M�d�0/��p�6�C�{b���'�_�Ǎ����w@��;8�B�����˭���bq��L�Y��NQ�swBP�����U*�즩������U!R���o����k����z��%�Je3*;����|�����Ε.�V\�Y6�|���D�9G��x�\�)���=ϱ��U���_��>�Z���򱆖G�������wO�P�Ne�/�.�+�Vlt`;��*Ս�V�w騮���8��Ġ�:k��w;�;zL�	m��7z�Ʈ@
�Zz��?��4qb�O�6z\�8?�
���n]��l:���?r���e%%K��X��2o�1����/�>��2��5�b����r�T��B���Cªk��J�����:Z���/�+�k�g^��䶹$��ȺE��c��hq���d�Z��t�l[jw����ͱ�a''�]�¸B��&�gu���_:�N6t�7o�*���7�������m�����wAN�.�w0t�Љ��}��J�G�_-a� ���1.��R��[?�����Z�����6�#��M@��ˡ�%֥�:p?2�Kh2�JKT������e�c�m�Fb��]���;G��´�O��}yS][�DkZu��bi��z���5�k�����+jwם9���n<�;��w:��N'�;9:�"H�4/ �%�����3r�����?U<��ӹC��������b:��߼9�U����٬)��	�:7���:�t�|��M&�������Éf�������-���jݪ�{ѭ�z�v����M\�i�]][#�E���{U+���~�Ye䂷�na��*�f����42�:���Z�C��W	mm"Ug+�V]V �]*/�T��jՏ4�%eM�k]�rq\�>�I �݉���g��Y��[��
M�T9L����dT��B��y�W���ڿ��/6K��|����ȯ/m��*���b9�e'֍dVN-�kVd�꤭�⭕�_�S��M|�|���Z�t��4��N��ltZe
�S���*����M3ȭz<�mVوB�F'U�������DA~ݿ«~N����	)�k_�*i���9=�z�P�Y��k��@�b>��=޾�C���Z"�zl_�۬�䶢/3_z����muӮ���ӎwX�_/W��r�o�^\-n{g+{�{�Ӻ�^��p�����^���4�m���>o����E'��Yx I�ʁ�Q2d�����[��:���-�իWs��k*Rِ·��u2P�՚�.�۔@%�X�Y��g˝i��c ���j�m�s.g��F�3���w���~AŮcfGu/���S��e��KW�ɸR�t�q=j]��J�Q�
�#tv�_���Mf��h�����j�jJ��ʅ5���e��W�h|�n��%�;�7���%��U�}�%�G�ܾsх����ڭ�;w�&詎G^��e��ٞ٤?mZ������I��A#�]X��Y�}���������g�J�U�۵��_����_���bP���В1tɇ�PUrR�~��F��R�f�-������s��I=*��/���1��{����q췽�Ym�vN6FV�� ��}����=ԣU�^����}�}�{���U�� @B6�����'�xBu�ťK7�+W���ҥKZN�����=�_�q�G�o\t��ֻ;�`ݮf���/�NQnXU�ޅ���h����u��뾿�:,Ha�.�� ����y���f���}��u��E����r��[8���W}˳���ѱ���F��a�X+a��de����ۡ�����Y�^|����P�j�52}��K�����N�ܹ�}�}�w�����o{��܏}<{"� �W����|D�j�����8��S���?�ښ�vaq_��Z����Y�����^�Z�Vd��tb�RT2bەZ�S���>�h���CDVՓXFP�J}ٰ���n�{o�f��X����5[��:;�g�=Y5o�~nj��C�a���k�v���i����'�O����1��6iN^z������l>����N�'�щ���Wj����  �&UU9���z�ﻇ���r�:��ՉJ��^-^�C����EGf��X?�.��q�Wן�ާ���U���7C�Tm����O��u`P���ʸ[}�:RX?�vm�42ۆ��OCl~��q�f��G��ʆ���5^�p�կ}5{��Kٵk�*u�p' '�����٫�  �&��}u�����J7�U^�eЭx�,m$�:A�e�.��DFg�5��j����2�( WUjg�0��;�����uU��)��j����\�=88��Z�������B�V�S�՟�<��a��F�r�~���k��_��ް��ݵdu�͸�y�{��s�}�v����M������:���U[?O�  �I�zy�ח�syk6-�_�2����=����UX�x2��+�b��jzm���:�e�l[}�߁A�q헶�ä0��R���؊���6�*�H�:GĖj�E]4��N��E���ܲjy�1��:e��yb=�Cp�#���6�¹�����*[eP���uϻ�N'ŭ�7�w���w\�~��X� ^  �T�e=�͔L��]1��u�ڱ�""5��0*�ynm1����-�����*�5�©"�:,�!~�<���6�,�u�����\��K����[���w�G�m�؅j�_�<(�n.�z�XJ�Gg��|�/��������Ϊ��\X��������5��*��k�e�n�{ӛ����UNX/  xMra���W�+��В�.���ɤZN�6«�`
��ԯ��[�#�e
��@}qmB۪�~�}a�׺�s��yc��_Y*[�պ?g�l��kCɄ��(����0q���8<��ϙ�]�ޠ�_�dݯ-c�ZY�������%�7jt�J|���Vh�ʾoK~ےӵ��w��������n��ˏ��-_�߻�^��  �5i4?����ߛU��k�^(��>غ�W-]hti�q�֤���[��j���(����hh+���U-5�;;��Ivxtd+��!HV�-�l��C���о�86C��l�e�Ȧ�6j?Z����Z�p�.t_kwZ�d�5+�]>{�Lwr2/6WZ���N���;Ē�\�~��S���1��G���w���B�V�[,���b��"[�J�r<�74��({5#� �פэ�n�x�_���_��|օ��;;��X�E^�p�J���j��{���P��~�+OW_��-�?�U��=��}����p��jaU6�+G��C�-Y�YX���*��Bo�0�M��"m;�W��teղ���[���!cF/�?Ѳ�UuG��Ԏ�]$4k�V5�[��j'V( �0^�r	�f+��'��mݯ-�<���VMS(�7��m���s�����j�*F�  �I}꩓����o���'�5��v^?{�֝w�{��ᡋ��I�jڲ�o\����hl�4M����|a�pU��nm��&���I���8�,vP���;�uZЂ�������CnKǮ��᝻�����+�����qպ����z��o�p����7=U��Ϻ����ϯeYw�e�Z���h��������t��۬o��UUu
���c�=6�~�����?}�Uۅ�OC�  �YO>i!��O<��ŵ߫�˟�;{��~������mU��Jn޸�����y晙r�xRg/�t=��̭NV�7ͪ�h����Z�ί̦%����*��a��H�3��ժlBAX�x�GV\[�n��K>�-�������j�TZ�򥋿��{���/��ɫ�[�
�  �����~����o����?qt|��.�~�}�Ѿ�Oܟ�������'몢����c������\X�U[lmo�m�~�
�y�}V���eEy�㰺]-={�j�7�]4b�FtZp��ߡ[�Bs�vvv���>p��d��  ���w����'������mko�߯�w�}��.y��駟�w�t{gw�p!W+�������Z��N�[�:�3�(�Vck���:,����wJ�����b̀~_u��z4d�u���md8��\ݎ��WF��<��"�  leG���O|#˿����ݭ��㽝��]2}t{k�m[[����x]Y�g����z<�N�˦�jc-Ȳ*�4�ۏ+�u]������R���&��|A]�}�v��ڲY6j�[�6c���ޗ�u�t��E�  �.B��Q���Ͼy���'F]wg��w~k:����j?��������_w���z�jh�]5�Cז��Jf����%���ٺ�¥-Q����E#*-a����V>Q���Y5M�T�bk6{v�/^���   �z��d�B�Y8��>���?\]�p�>:��ݹ�X6f��}���s��Z�u����e��y6�N�f��J�ٵb����K��:�땅\?��N��_<�]Y�����lo��l���gxY^  �?��a��O�z����z�֢i�Z�L��>�v�FE�/gp!�V9ú͖��|���z����4q�~W+���$6��+{(;���C����~�����/��  �=R��G?�o�m_�ON��x<.��R�V�$h�Zۭ��A_�hnݏ�f���P�n�ZݸR�-F�g����#��V�Oo�^w����u���  �}жu]�#���B�vb.׶k�f���]��[(�6
��l�}��P�տ5QM����il4Woom���Z,��s�ۑ�9�"�  |��=�r����^E�   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   �F�  @��   H�   I#�   i^   $��  ��x  �4/   ��� ���=ׅA    IEND�B`�PK
     mdZ�+s`(  `(  /   images/8a1d81a5-79d4-450c-9f72-108cd2673013.png�PNG

   IHDR  !     h@~   	pHYs  �  ��+  (IDATx��	�U��Ow�Iw��C��" ��!�@AP��EDAYUa�W�A	� 
*02��8,�2�b�ٓ������K���;I�[����w���[U�T��޳�gp2Ƙ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!�[:	�9%��f����Bw2f1X��D�KhI=¡�5�~ww�{�<˵X�D�lii� %$B[��tϙ7o�d���/�����̙�ؐ!C�5k�S��H�A��y�X,B&X�0���c;�d��3g���������D^�����
�::���,����={��6��k6?�zD���s�PX�.���"���ں+°�ܹs[�O�^��6	GmY;����_/B��-��Q9rd�4i�6�<x�xhw���5�7?�B���3��Eh�1
a�18���DxS\J3f̨	�СC"��V۶0a�gAR�+,��5j�:��!>�6����u���X�7��6����/%�',B�V'�������,��Gb!���LS�N��!��tꑀ��z�Ҷ#F�)S��DM����-[Z���ؿ˯p?�r�����٩���z�&�"ԼDe��q���F V����]lK]]]	a�	����Ӵi�j��ՋA��7�,d˙�l�rk��`��r�~#���B��V[��E?]���m4x�r�x���g/'ӴX���yd�� _&��$a���Y?�_� �zX(ai��^b�#���r�?�J�D��v�ʛ��l�H�FV'�Cp6`�!�!�ۢ� �G��=�$�Q�v�h��Gr�'8�Y�������d�
�P���քo��7���($KD�_V�,�h� Hx�6�c�������}q�����n����
�>oMX����y�b��,����v���5_���D�L�@�u�~�LSaj.��3������F\E-Y>Qg#q"c��v�ob�
��ۙ����g�A��`��չ��ҖQa�b�,$ݧ�[������[Ա��d��P����q�QS�,	�ňe�ԩ�c�Of��C�I=���\�ųΥ,/EX6ClGh��:�N*��a�I�!F[�<0߻�8������~0�B2�0e`խH�dU�U@kI��s5��������+ �����ܯ��B;A�F��$Ha�q�Z����7�[�*�E��a�Ex�Qf���bPFU�2o]?�Y���		R��L���������������F�I�<����kl߀�O��b�Q�RS�5dȏ����Z��o����l;��?M/v5:�p��<�8\�%�����Bd���*���D��"T=$@ji�H�d��D�Y
�(�P�KA���z�y�>��X=_$^'+���B�57���q�$|��d*�E�Z��Y�L�c�[�g��㓋`���@�ݖ�_LQ-���x~N�E�զO�����ܲ�����d!��꠺�6��7�I[V@X@Q-Ȉ�a�?�<���]\7�*���=Ԫ�g����zs+AM���`�R��m��8��y���8�c)5]%m��x�x�D��@pц !�hʔ)�O��R5���P5@{ڮ@d>���h~��^�Df�q:2��o%�U�)�9�&�ZqTB��	Y�6g��Nթ��X��}^�@1���5,��yd8����V�~�19?:'wb�?�M�Ѱ�T$;�pR�54��gW�����/��1ad�����Y{-X�_c����y�Ơ�h��,5PV�"��N�a�56����_I1�U���dI��M�v5Ǩ6�(�8�1u�T�����DVbt�l���H=^ Lbj\T��M�b0������Xj�?4%{ ��Ն�_��S:�*"�F�^�Q�}����"Ը�ճW�(g`�������T� ݈�!����/�H�eɳcWW�ֈЉwZ2�E�1�C�S����8j��.��ԣN��'b�?j��-����'"N�&�PX���g`�M�1#;����{�Y������Q�����j�G�wc��������c���\q䖟��Ν{Q2����I��)�n�kh����d�Pc��/g��	��1F
4��Fûru1tvv3u��I�U�.W��ܳ��OR��~� X��	C�}��Ř(UDg�����K ��9N�r�*�Mc�4e�{����d�P��J9��uKtHԗ;�#�J���d�K�Ո�]]]۩nMC[T���ɢ���3}�)�E�qؖL�M�W";&��H��az�`,Ig�.|UG�s�r�?����"T��x8ń���T��4�L�>�[�����G,�1c�v�(��@k�"}'��1ޮ���Gf�aÆ}PM���K�ئfe7)��s���(�$D1��ڑ}�&ww(�E� ��M����ch_jUDO\Ɨ���7Ѭ�5k}�-�CX���X&�W][�q �-B��������DgԨQi�����G��Ͼe혫VT!�W�Ƞ��y�k��ה��R���ٳ� -7�n#G�L�[��m�0´d�a*V�Fd�%BjJ������.�Kh�G�{h��8�?�)7�<e�w����灲��5k�f渄 QjIկ7�1q=�x�Q\%@*���ٮ��?N��� @�"<-1џ*�s�|E�a\B���Ɯ��ٹ���Q+\�Ov=��y=�p��r�P�D�ArN�./���Dl�V߫�{v��[���z�BX��2�1:$�w�<�����{9��E'�b�Hۢ�R�9��l:��#F���)��^���1U��ފo]ˣ�oE���}����	V�>}�{�eV�PqL"@&ш��\�؂����$4 -��(SemL��1k���x�Kszi2�[Ru�;�A|_E�WԊ�6p}7q^��'S�PA���/��y�C4~�4�V�?�z��ItBlDv�U�
b���B:w�eT�u��F~/FW��UZ+���;�Ϊ��;�6a�E��rhx��$Q�.U�"w!��q��F`vG�&��ڢ_L����%!��?�Aמ�5�I1p3�dg�,�qQDT�����s���T-jiH��&�B�֪�o�䎋%���q�X�Det��`�h�cY��A<6ͭjr _+�I@$$��r�ȟs�)�/�`V�����7GK|�2���-��R���kܙ�C-r��.,¹�{M�g:�Y�eլ��А��J��*6��,�9+�/Ǔ,�zL�fg(��j�A1,,�9��b_*�Ǒ���*~�05+{���|�c�FL��/�s�;�Ly��:��H�Y���s�>Ǿ/UkT�޷?#�S��F��{ǵY�!���=��|�v����#G��ݛ�󼷫�K��%n�����?/����A��2�02�~�	r����?��Լ�%ֈ)jԃ7�|�}}�����j�#���ٲ ����r�;���:J�q�a�-Bv�3^EF��PT��6���,�M�^�>��=OxN���ke�,Q�ZjnE���{��D��b�7Dh%�ݑJ���|��o��E����B&?�����5�����9�|����Y�D�DX���C�o��by�峤Ooz��U^N�w�D_������v�Z�-���^䏼���V'?	��M���i#�Ѽ_����l�MF{�x��1 ��Ѓ�	!�j��g���ɓ?�hy%��3f��o��ƥ��޼�r�;���?EH#��䡫�fe֕C,�j��"}a?G�h����&��X5�]�$D��ɟR�*H%@[s���v	��~�/"�W����Go����?YF�u�Q��-h��uCUr��(��@��d����oGt�{�7-�~�s���]�'�\S&M��z��q�m<���x}d�ŋg������ROeh|�D��e����ya~Hg]e��v��Cc#f�b��;6�ڎ!C��z�d-z~��4eg]5+((W6N�=ߗ�{�{��>Z�t���X.1.d]����* �Y+r)��#�[��
����:«� �}�������q;S���:�E�엻�����r(�M%@���*r���n^��Y�E��D�hި!��������,�����k�8j����d1z�ךC&:�߭�:%���T����	]���n2�����<:�/QY�K>�k^L�O�V�gb�������L�1bĚS�L	�S��}�V�eq=x�k�L�7�c��-�H���>�ǻ�!��i9�/"Dd!�h��p���������1��d�.���"���Xw�@ϴ��c�m�7�߆4���2���1^,;ڊJ�ތ��GD@��k���F�<���J�.��y�%�7R�սK�����p���f���O��Rz)�n���2aK>Ӓ-̆k֮'|Oq��������Z���X�H,qQ��?�����~�զ�d;�/�ٻ����v^u�_?z��`˘w��� ���"�$�5'm�S;k��q%-"�1#�2�"b���l'H��;����u����G ;�W<Ԫ�
�'��!��k��JS��R�3#�E���>�������Q�]u�E���^�h����x��#�ҮW�x�@;>��"BS�NUѣ�#�_W �W�	��	/��K�Ҿ$K����<wX���z�&}��'�[�`_�+�8��^�ճ%%��Z�ukZ���E2�7�����<-�h��"�eBZ>ŲZ��;�[B�YB����n ��0ߧwl�gE巼�y��f[���8[��,DUi�s��*qS��u��?�:3���}�?Dh�1X���!^�ړ��5\���4�Ǘ*��zѵ��cR����z�<^��X��o��|*�uq�S��9�4ە�Nშ�(��*���&h\�ѭA³e�v�}�"��}�^���R�2o<��f�8khq��Ҿ��#�#��Ļq�7���u_.��>.�A��	�`'�r��ǟ�@Y}�^�0�뚞+�'�k�(Z�k��I����,�7k&	�Ϧ�G+/�2����)�*nZ�/������Ӳ&�s�G�OV�`\hs���|�rboNE�z�n1<%����E�gI�l˓z�	��V|���u���VeJ�����"��E݅�9'���1l�;�r��t�"v�آ@B������é�K�9[Xf��Nc��Bs-5��.e������Ձ1��?��?�B��1©<���d���ٜ��o�Ӳ��T��k�b�k��ݽ�8 ����L_��F�j��Q�]���UK��?fi-%Y;�܋���yd:�ng��9�����3~�;ᷩ�ⅼ���S�׾�Ғ!۰�N���DU%�::v�s�1�i��{�����|� �ePŪz8�݌�!���ZgRjxw����=�Qct���E��ԛ��ep��Ѥ��
��B\�Y����߅�5�������$T���(m	���ʴ��4{�x�D|�����K|�<�q�&Mz?˝S?�"�y����}/�fi�lp*�|�/�|0�zZ�*=`F��������԰jj|¼?�L��V��u	�����l�@�ETk�D؞pvi�5Q�v��pd�n��u���s�u�"�'��,� 58�<��xG��k�	[�G���}��}��T藊i�����r���m�E�o/��$�ЇROSs��%�f��^���r9~��K��+��E~VSW�<����� �͎�.�yF���P�ի�ZDmP}}Y]�p������^���G���E�^X\ѫb�M'�|����^yh��h��א[�A�'�C�$}�"܍9��sH�q۱ ����/��z���y�2�3���x�[�F�+S�#�=�=����ٌgv���Q�T��C�I|n�Y3O��[7�"�.V�<*j�7'��--�~ȾK{{Üs�h��� �ٝ���9�ۍ��S��#<#8^�po�3��25�m��ѣ@���a/��XO�%����2/�*9��f/��l7��e[_=7S����<��z�wD�U&�Eyi�ު̅���q<�M�-�4��h��<'��I��j̠��M��F������2���ėZs��K�U^4x:E�^�T@��U��<��ݺJ�����<�ߓ�����<�����r�����N��s k��Q>���D_��W��H��HYH`��V�R� �q�����d�,oO=3dT�a�T^��4�g8.O_=�*b�Z<�;ؿO�i����n)�k��H�5c��h:�� �b�!����>���G�Rt�Рa�Ϥ��ɓ'��Lb�;�d�p-�����l�թwr�Z��BIϊ2���a���@_���"���?�r�$OU!Yx(��dP�Ft�$�����l;�m*F�ú�����qٳ����<C����z���vWnQ]��=�-bu��3u���<���XYH��w/%E��-��P����?,�U�%���B�׫8+��}+�����,��ʗ���iӦ�N����gf�`K��C)����$�����d��5�N��*����X~�l��*�ݗ�%�{�tG��0e�\T�6�J��~/%.È��e�De�P������ů�]7�`~Ká^"�e�}����"��!;���K��ӈ�|���wS`*��x��<�M!3��*��Y6$��S�X�,�B\�c)�l�����i�e�Hl$@��$f�H��_i����s�^��ա�~�q�e��0u!h�y��"T}u�%�=�1Pa(s�lO=��(B!���U-q�
�Y;�aŠQ��n��8� q��R=Ӳ�3�-E��1��
{��'P1,B��>�7״<��Y_�<�^-I���b�b�݄��iX; *m�.b�t�~i[�\+�!���y�|K��t�%/�W��<Ѥz)V���X�
�%t+Bt�(|��H�m������oM�QS��X"8G�f{X��i�,"�`�����&�QO�e%
c�$&�����/�ŧ(�� @�!���z�r4���n�?+Ue����d9���>"�. �e��H�%��:e9\O�u�DHT7����,��X��#_�j�_/\���!�h߮��f�z42��8pd."-���A��H�?U��Ρ�!��6��Y8���;d��S���}o2ʍ�9��㾥a{��m��Q�=iN��3g~'�(V�Pc�G2ƭd�D/���V�ݚ��G����45�
�9^VP�K	H_�+��X����J3�����]���ނ��ԙ�Lo�noo�V��c�}x���L�!�5d�[X��g�p�/1�n,Nd]�FUl�/�~bt�5T'@�o�"n�5z*n}��n���gmc�i"�K�YR��x���b������YLJ��X��p�5����XnT7��֛k��iӦ��s�D�/���L��w������W�c-@�E���_e���_�u"�c�l��Of��tZ'�˝_�&t�����P�1��	�f7���<��c����dފ	��g�ϕ�HUL����t]2�E�!��b�����{�p�J��mpY�����TRm�c%@yN7�prB�����"Ԙ<"^d�3�e'f�D�FR��1�!�az�&��r5�:j���DP�Wt��L�ajL��4g#DXn��y����˭L%7n�O���gΚ5k��-�$�y����/%ӐX��yy�_�U�/{]?��'(n����4�Qk�&a<6�p;�AnaT�K��2{ɀ�"��<L�:���ZQqL�,�ȓَ����o��[�q�<	N�

?ҹ2Z�k�N�a�5>� >�"S� �J������.E��хi�(�œ49�������ȑ#kn:�`�k	_M���U ���X>����}����t%#v�!����¨�r֌���Ū�QŽ�b�|$@�q���b�ip,B�@E������׿6Gx�N-@Йr����Ss#+����h�*���2�il����
`����Fc/D�V��T�Or�2�QXkS4�G�f��՜A�]k�'>Se	�_�\���]���T�P5�1N��}'D�7�ѣ:�)ڍ�G��p샩9�f�^q���F14f����veߓ�T�P��O���p`yb�~��!�E�5X�!:�㾑�],�x�r6q���
�8��:��IDiO���jϤZ!,B�"2�F�O@�n�SF�|ﵺA�B�<��F�c��RuP�Rf�:�ͥ��6�	(��zd��\m���QP�Lb������OF�.���ڠ�E��\P�����%_��\v����b�A�N!�=S��Hb>�$@���m/��&SI,B�f��4K�U0jԨ���z����H�/������������mν~���gm���F]P�B��'�ǧ��T�P��H�SRO��K&O��NeV՗D3�2���iWD�N�$�d�k)�\�o/p��%@����P���b�W�zP�|jf��믬j"ś��<��V��%[.#���欛bYV�*,O �ű�s����ăC����	`,�!,�?y@?@�c[B�gKU\n��Ϥ��B�gm,B�'2��5��BT�c�����5eEV�Jd�<�D;a�hD�E2����V2�*��J�8�wtt��z�r�}��hm�!(�֛�%B�#�{�ߝ�%wI�}Y�� �P����z�ȼ��<�.k(��š��>U�a�{���O��i�osx����߫���\��� �V�Z���r�w��!���T��:_`��=*����=i]��u�".��J2M�E��1Rߠ�W��O'c��b��%��%@Q�-d�H ���,�U�sS��F�ʶ	�Xc���]0��9:��ƾU�M��""2Z�sJ�t.U��ꧢ�=H�=Iu<�����S������,�P�3xȢ�GM�h�g�<�kc�,��wɳ�F���P�h��fyu�<#������N�&tL�S�]��G�#	��1q��-�v\\����mrO�A��&�"40P����,Ւ�/��d��"�KLd�h]bT�,�y��J�N�rS��b�����#�c��%�Q�\�i�7�5�=�\�3`�,���&�If���m���RvB(�i0���N��:����]�_�"��џ'�$XQ��!b�/��W�흈�D���Smz2���E��?A~��������KDB�oC jC�%
!R��H˘RG��(���߅���uq�GRO��_�#L��f`b2Bn?~�@�<��LXkg,�w�]eWTgG�dt4��$b0�Q�fO�<Y��+��ˈ���{�}������.6Z��X���А���;c,�!8�XvR��4�#YoǺ���B�fp�,H��S�)X8�T^Tݎ�}�E�,�p�!5z5-0PT�/Q'V��
��Yv�a�+!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ,BƘ�X��1E�c�b2��"d�)�E�S��1�(!cLQ�o/�9��l�    IEND�B`�PK
     mdZ��/��  �  /   images/aacc0029-e57d-4614-a443-d9bee65b5175.png�PNG

   IHDR   d   `   �s�B   	pHYs  �  ��+  2IDATx���VU��~�� ;�Nk�}�N&hEa�i�1�)h6�#9���$��A����:�4JEѨ58c�|(��|-���l���yv�;��/��Cs�3�<�������s�sιoq�
�g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g8��ӧOR__�'---Ikkk���� ��/**zOysssr6�=!rj�~���Ǐ'���I����>����(D�s��}ًlA6A�nd�(-"=�-!���m�t�A�?e����}�����sU'g�:�TY-ׯ#[�^I�:|�ԩ)�Wb\RRR�455eH��%8��3��PΦ���+�&���Zҧ�s�F�c�3
=���ݏ~�B{���D�7�#D72�(~��c����F-�٫�8����7�n�!�*�7q�'H?��S�w444�KdX��w��A���_%���i7��觑#ANM;�&u�l�n;E�I/�}�{t�����Vz�3�^�x�;B��{�Z��p�
��"�G�y�3'�� G������$�嫹�QҚ�����/���!D��0�_���Ƞx������۷/�\����L�"��)�V�����;��@s���E<�0u+D�"8pA�E>8���b��8�1����ݛ�32r�z��>v예�B�7UO�-�6/�I�	1G�a������z$DU��=����?�⫑��]�s��F�[Y㔉8�#��$�bsFOA�4|���N��ȗ����~�rM��D^	�ի�mm�!"�!��zEEEbÕ�ȳ^�K��������O)��A�G��wԕWB̙8f�����/�#�V�!��	��q�ku��wg��dH]���)�"�9�Vg���䕐�#'�,�ְ��z��"�v�nCC�?R5٥{mu�@DJa�t�k��|�I�$$,��V��9RN��2W��R=6�}�~�F��5	ɉ!_�u�P�U�?�_G�+�%#U=�h}R������'J�{f�'N��zVB�6�����9L�z�g���}�s/�]H��2��lޡ�)�?�tϜ���k�q�C�gI��p�u;��O� �	�Q�%�ڙ�S��Z��{�o�7����,k�����'ON�n��`��FZ녆�R]6�=lB��8�/�7(>`=1s��N��Wx�ˡn?�h�s�ǒ^�5�I7v��H�n��γߡw�$]A� ��NsG�eCx��m���vmvG���_Y		��J��а�Q���~[���v״�k��ѡ� �7A����B�{�#2l�뉣��I�Z.�=��9��=)�q�����~Dccu(���Z���t���J;�B�o�g�ڌ��MB>Nن$��!�|�lS"�����+)��5��{��B���%l���9i~U�^�°����܅V�:��5���}�ey�g�˹�a�;��!�詶P=�w���VB��4���
�)ߢ!���		����љ�=0���gl/�QK[S��}y���
io�dǩ�kx�����9eʔk�-[��H�&}^|D�[����r���2k�TP�i.�1��{5���!���1�#ȿ@�v��l.
m隉�m�_-�C�!�V��i�P-z������?1�-4��W�W��/j!�L� ��`g�2�ql�K˗/�f¸��zY�4K�����N��6�!�H/��0`UMMM�,��ty �'����No�����c��
F��!�m��!aVc�y�+0|-eu�&��g��~�Ո��՝u��!�t������i����n�vtq�&��8|�NET3jkk��0 �)cN����QZ�,��?zmYJ;N���!���߮�m���{U{x�[d�cW�Kݱ��0�%UUU�I�H����㰫3}��D��,�l�1| 1���Bh�vz�+d��HjnKl���v�T�ra��<�	����Ӈ��/㐗4u���D|=/yw(T({Q���L�;80QO�n|0���鉕�>��y�:	a�J�u3ΚH~.����PYY��رc=��/`od8����y�@��#G�藫���0�<���1"ټys�/�[��%�)At��H[��)۷o��
}Uer�m�{!}��I�oЎ?��|�!�;�C4l��,$}/i�Z��a�9��q�-��y����{T���y?�JB-�)Sѣ�yJ�<�]�ΐ>?Q��SC��yR��7�Bи�]��HК���{�P�5b���Z�� }�'�ƞ@�	,6��/�moh��z#��-����VGo���U�]�����R�؞�攲��ǉ���-b����c�l~�m�l��?���/Y��	�|�h�.�q�x�8P����xq���e�Y��ZQ�~����	�4�� �d�i�X����lV�s�(��"ذș��u61����ׇ���}mXP&�^c���Շk/�j*6�#����t�g�p�r���n e%�uhmNC&Q���v�.�-h��hX[��\�\�}��a�DkA���~Dz����IpG�`�
:�ӗ!8�	�x���%7�<a=�vSAo�\I�R�&�ۑt��V�$�`�a��'?�S/��bm��� }�\��Q�ꬆ�:�ۀ�[�7;���kB���R�\d�i�������a;�-H(//�,���N��	i96,�2V/R緦��E�ꪫ���	g!B�M�����?��F7W����?#��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q�H�3DB�!��g��8C$�"!�	q���n*e��B    IEND�B`�PK
     mdZ�1��� �� /   images/1d90a712-93d7-4555-ae10-1782f839eba3.png�PNG

   IHDR  T  p   ৆  0�iCCPICC Profile  x��||eE���Vx�*�g\�$�{�R�f�IvC�]�%�lv7��l��U����E�4��)"ME��   �4AiR��=sg��E?����d�y�3��)�s$���_�`Ψj�̝�h�{���{�U�J2:�T�͒/�,\���Ց�'�~��ǒz}���J��~֝1�p I�W,��K���- �~��g?G?K�0��g9z�J�'�7q<�ݭ�S�d`���>Iƭ�?�ha��������sA/=a`ͻ����;c�I�*$�̚�x��ch̹���A��$c�\�?<+I���g�\�FЭ�m�Ϥ�%�����2���L�Ve)cͩlf���:�����y��C�4MR2M��4�1�5�kʴ\����Ӕغxx�ඝ�{Y��"��t%,I��ݒ*��,iƫĿ,1h�HZ�Ix�:��&��;�%�6I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m[��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����,��qA��m�b��(I�x0I־<�m��d���䶶H<os
?>Y/�*����������\�\�ܖ<�<���|аJ���a׆}�5��pm�C��Z}T6jڨCF]6�ѕ�;���ţ�����1��yb�cg��b�?��qG�{`�F����J��x��V�b���X�UN���ʌU��j�w�ֲ�-��կZc�5�Zs�5���'k��k/[g�:����7�׽�+����p�m�y�6Zg��7�k�1�\���6���͏��~1��m��~�u�J~��[l��V�m}�6�}y�/���EM��w��W{�+I�ͮc����r��[O7]v�v]_����w�񀝎���-�M����I��y��[���>���w���η�n�պ���K{��6a��ݯ�c�^S�q�7���侳�~c��N���L6����۸�����l��O����[,9���.?x�e�|w�CN>l��O=r���>z�1W�k�=z�~'�;�SZO}��#N��ߞ5����\r^������{~��ŏ_z��G^���Z��p�'�=u�/n��/�~�˭�ܾ�����;���{ο��yp���,�����ɦ�����y~ʋ�_������ޘ��No�w�����?���-�D�X���3�0
�]�ɇ�׍�`�a��='���W�4n�q7���Ru��W��r�*Ǯz�j��~��׼`��׾}����z����kn��F;l��&�7=u��o~����K_�дE˖Ӷ����m����^�ts�ǿ�B�f�o+�5�zzc��m�n�f�o���;v����>���']�v�ΏM~i�w�>v�M:d�nS�N=������~�w�i[M�e��{�����7��+�Zѷ��[�o�ϔ��s�<`�wf3��}/���9��}h޳��\���*7^Դx�%��ׁCK�t��g,��;7}��C�=���W9�z�8j���8z�1��=��?8�ǟw��?���kO���מrթ�/������'��s�g�z�~t��G�sȹ�w�����'����-��܋g^���/���h��+߿꣟���r�:�nv�6��׷��q��7��r�慿Zv�Q��x�Y�_t�տ��o����w>����z��w���������?���{���{��?�������?v��?|��?��§�yzڟ۟��/��m�����?���^�����m�+����߫�h~m�ק�1��ҷN��eo���s�~���><��?��֏�[1Ɲ��ɿvo�a�&������/��5�ͱ���t�����J�\���%��������k���kݼ�=�<���������������	�]���'��֗�M�p��-w�j��{o��ˇn{rӏ�^��+���gϱW���ߪA�7��5�[���o��rǖ��|��-�'�z��]��o'?������Z��b�W��N]�u�n�u���Ҵ1ӷ�}�{�y�^˿q�7��?}�����o�O6�6c�`�̡Y�g9tھ�w����>5����ko��-j[����t�qK�9誃o[��w���|�f��#ڎ�����;�裎9��s��q��	w����>鹓�?�S_]��io�����=�3�?�}x��|p��}t��?^q�xQr�'?}��]�Ko����O���+�ꨟ��S�>����~q�����ȍO���/_���z��nk��r�:���7[�6�s�ߵ��{���u���ܿ�s~?�����8��=鏧>���S�8�O��?=����L�ˮ���\�����~a������}������m�^������.~��7.y󊷮���8�����{o�k�k}8���Ώg|BH�#�Q�Zä�s>����G�ї�i�_{Ӹ�ƽ=�ܕ����ʯV~�ʕ���ڙ�����k^�ֵk߶���>����_��FS6^���Mo����/nո˗fN8|�s��q���~y���]�i�扵ݿ�o�,;���/W�[�=�Q���v�n?f�uv�b'�������:鲶_����o����&����;�N���[���ݳE�iӏ���=~��s{����ߒߞ�7k�C�O�犁�g<8��̧g�0�͡O�[mΦs���8�kA����p����r������J^{ل���~���C�v��q������Ǭ{���Z��<a��8���'|ʲS����ӎ��Q�}�1gsֱ?:���9����;��������p���s�~�����K{��.?��<��~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW��U�Y��U�w������s����`����������cW?~�����'�}j������g��������=��#^�ދǿt������W��ο?������k���[;����}�9����]��߿�?~��_�譏��ɇ+���,/n�$����]�b�No'�Ӯ<��wW�x���a��R���k�L�R�H`�k��$[�̱j�Ks����#u�l�)y`��������%�Z�Љs���־w�N}'���ڤ��������8-I�w/3������u]�N�������x�ۿ?���x�̞l�����񊜡�!�*n�Ff�����+x�O@����D���W���������M��Fo�����/�����o��*_��'���c��㎡�m�W��#g �N��޷S��a�! �~ ���C�B��9x�-��|K�_��	�v7����x��k>�b�|�x٘.;�LaaB���}�A�U�����߭+Aֱ4�m�'�lP���T�jK�$�����o��ȍ�7"����T>ukjA>����AYƀ[ǀ�	��ݴ��P7�N7W/z� ���!�)U���a��&��u~����X�~��,w�����\Ɠ˰i�
�>w%Mu2hQ�IԞ�m2�N�Q���c���\��ȌdD��q���C�&���Az���>$d����fh�Z�'���t|
�RY�,��b��O�!�/��Mg�5��d�!e�l4�W�1���,��6n������>��m>�b��;��bNV䝽�Z�V*��zZ�ۻz�vW[�g-�3���?gh���EC��U{��g.���^T�7s������2��}r����]g-\0<�?��������6���ӿ��ٿ��L5��I��d�:Ј�������v���T'��tu���X�i�2���oR{g_Oo[�$1��ή���m{m�sZGo{c���jc��}�Í�ޖ��m�}�Szz��u�M�6���=�h�:�U'a�s��v�o��Ο3�s���B3V����wϮ6��sw[�.��)S?�-=m}��o�X����jk��n�ȻuL�Ԧ`�X\_�NVm����̘�jmMp�XZ�R[˔��4V�L��l�h߫mR_�Ծ=��4�6����X��>�mj_Ǵ޾V0L�n�m�:��kjOO�Ď6�T�؆�����胈����Lo{*�K���Ϯ6��T�[���ՁP��U[q��gTZ4;H�Ty��l�W��ͨ�'���Se����͝8�����6eR�ܕ�{ں��A2˳>�4HqbGK��B;�G��6����o����l��Z�X٥��7��x��}_�Wml���tN�ڻ������]�z�v�ֆc�6N��m�{_8a��5u
��}��V�L���݇�����1�����'�����L��[�i���pJA�������u5ɾ=ܿ{��rB�{�=m�=�L�sT2�v����Z&4�#�dk�Sa%�Z�״jT-���U5�Së�ո0�����|��OV���g�"X�E�1+MZQUvSߏՌPR`M5��Q�)SVWtU���/c5�,SUY��pK�	&S!*&J��%3�GGX8��S��ظ��~R�D&9��(-m�*��J��t,�,u�gBXj��GF+�⺒�И�?v4�yVe�k�a�c��d#T��Q�Qe5w��"�i�0��2��T^�b���Yn���2)-��M���(;��1���"���L1[5�$�}d��������יѴ���(Q�T�1�����*V(3E��A�d��8F�4V�Ɍ�c��:�d��wj܎>K@����u^� �h���F,˔��g	�	�&B2�II)�
���DZF����f������D�љ�)��ĖZwdҰ����X��L�-�z6)T�Å[�)�Q��pH���� �ɌT�&d��Y-���:S#�z��!�&�f��c��3���VO` �rͱZ�o�Z�yjmN!�0jR�z�՘4�\b��6�*�ak�����$U�,�*+p��aF�jR��	N��\#�q� �V*���he���5�2)�r#`��=PY����	I�]O��X�m	��b�ؗ�}a	Ο�贄PX2�P9U#�ġk�R�
[�X6�hN;�#�feʉ�ڹcq�O>�s��#��I����N>'��N*h��,�B=��$�!�Ԓ|)�Nji��n�c&ͬ'���(�p�b�Y��*�5o�uDF��Wd��֑��d4#����� mWp�ďȝ
Rc��0h������ؘ�QW3�0PZ���P�
���{������V0v�c���P�GW�4��)X6l�,��.�9X��
�!�
�9�[G����9~��;l�(HѺ�f�S-S�e�)!x p�
6.!j�T����(��?����g�(�����"��U���6U�TBR�
�#�g�k�C�GX�)q�>@9�(^{^G�PEi���p��A3�6��[=� �i�������a��hH��K"�:�+���疤
5�)Ed@%@�f�0�Ԃ��@�pĄ�2�+8#�j�FZF`|!Nj{���6�8Z���7VuA��BpO%N�W�)��J���F��* M(��JI��p\���mf��RZ�@�H�X�V+1�_G��Y/!��R2L�,ڈ
,E���u�$G��¬�z8;�pxX�2�����$M#,�(nY�$����q1����% �T��qdX���i�F(%�:��f@V
SK:@& {��ZJG�CiZB?&9��ٚD�68����#��B���Bt *��U-
K�YOh�m�f�U'U�ۑ�`�F�wrHaL�>��@dX*2-�aF
VO�&a���dH�Ҍt�֎��0Π��a�a�{p+`W�ϑX=��4�גpp��wX�EE���!&: u�"$\�%,��(]�5D�����ı S�c� ��)����W2�>��E$geK2��[��4�I��L�ɠD�ӒL��H~�4�L
���<p0L�_�+Dֈdڥ~��5���e{���*e����8t�đ�U4���u�b2M^�B9%��W-�=:��Q��:H�'���j*��b�����H�#+ ��'C2���U}GA����#�t�^
�uI���(B�(��(��g��z�-�'�X*2�|]8aC���
$\챾#�#<�Qsʩ0�Ó|3b��%eq UC�AHڎ�,EŔ�q�9��!�������{8VSVȉ'�����J���LX*/Q�(.8C�����<�BF�E�!GqQ���cF�f$�.Z芑%E��! ]�<���QM��|ᨒ�#� �t��
�����[�*d�xc=�g >H�E���H�tMZ,Ք�1�����Fy�&B�V1��Y��%�֨\J���nIu'�i=��u D�����Uj5:f%�@�`�P=red.��paι���� eU�:p���:��d��/�� `d��i�@x6+�XZA��?F$Y\80��2b��T���9e��UB�����P=^���c\*��8xPޒY!]� �V��Ǒ
��"�{��b��2:S��& �!�:�hH�(�� V�-q�EGAZ�H�sN
7I�V�Ҳ�S4��"'g�z
"�U�Ҭ�g\,"��J���L��|�
I�GV�Z?�MK�F�\�5�r���K|kT�T��|�����@��%�5�pF�.��\��\GU����\�l8;CU$��'\zH�=���EO���\Ru&���qFs�U���%�=����� ST=�j�EONY���*ydEU ��1Z�-�:~��6p�)%��r�YL�d���b��e������9a�Գ��{6v������M���'+�& 08���34�=y��D	Q��a�������K(=E��B\Flir���irƥ�lG֔�{"IǏ�'�Hwa��o�T%�&@oq��q��ʼ8_M��%3�ۃ�b��V�9��&S�l*+�AظO��lJ�3��L=��9mI��R�|"	@LU"CY)���be
0@CN�ƔH��
��²��b�p����"�p�1V�5�e*` -�s��6N�SF5錕=��� ߗRM2/��:`=\`��g$�p<B9-U�Ud�J��%^3�SQ��rߔjT��D�r�J�f�d�v-�Ne�ڒ1]�5�JPq�lؐl54����֔@ˢ'U2*i#OE?
��dX����k�U02.:OH�Q�N%�IoyiS�l��xIFu[x�n�>H\�����)*�k*�"�PO%��J�Iт�)�r5Fኍ�)�`ٜ�)z!*N�*�@aX)=yL鑘(�&QBS�Pw���fS������ğ��fya3��ss"��<y�����%'8Nk�uC@���� Jz�����?���\����l6��T�'�/����^II��i��lѓ�}�]	XC@N���e./����?9˔�G:Lm1���\A�	T>���y�U�'�,�����9HZB`,�r)I��5	5԰�
���5��ꎰ.W��*�ɍ��e)|�I��)0r I=%�������V�5�
�R9^I��=� uTCr��X0C���2Ms��}Cڢ��R�l�}�O�Ӕ���27�M����C��
[�oG����U�YQ�Ӑ��e�5�Q��<5ݏ �q�!���[f%�6��R�EO�$=p��D��IVҳ �
�vT� �ߑP)�[�K�m�	T�b�S�`gy����S�[��(�
hKF�`��=�Td��~����]ʧI����Jz��39��T_�G����2Y��>i�,/=��J�?�GOS�ocO*`[Jv32q����0�Q��I�  F�ψ9=n��JCB�4u,.Уz"C��j��V�a�L�F����B�\3�S�+�g�%��
�8��È��`�);��)^��O{��y�f��H�4^�%D�J;��pY��H�M�,�a ��E*3����jUYRU�kK�\:w��9���.U�����n``�0���m��}���7R 0x�D����C�C_�!e�BX�	˥{% R���(��2Oغ� �]�/��'�YHH�С��p?Tc��VL*���0����H?�!��j#�I�:�r?�8!������TN�tY�4ܕ�'�7-J�1�r{� �	��T==�AX��7�DQAf�f�,.�U�&��݁�4�dh`�SWa{�/�_����{����IlXn��ɪ��ϭ6/r�a��q{�6ς��6�̈��-��Y�y �K�U���dPt1D4�;`����DO�讑�HXmރ��5{�������?wh��>&��x|�������}F^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� WuQ���   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    T  �    p  ��    x       ASCII   Screenshot(/��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1392</exif:PixelYDimension>
         <exif:PixelXDimension>340</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
����  ��IDATx�콉�۸�%�R.��֝������_��V���$�XND ���t��v�R���+6�0�����e-k��IkY�Zֲ�)+��e-kY��Pײ�����
�kY�Z��BeԵ�e-ky���Z�/����W�E*������+?�Wj������Z�^�#�� )��~�:��^T�#��J�_��m�P�B���kP�? �����S�מ���{������)��⽭����
�ky^9Ÿ�2��S����,�������.�[m-g����k��6�y?Q���������S"�)�h�;�/�����b�<&;���%�+U%�Y`��$��\䬲2������W����b�����m�.�z9Su���dEȿ\Yu-�+-�{�H�8E-�粒�K!���ŵ��.�:�{��r������31���Bos0]�YU�[9y�s�t:O�%��F�tc�����
�kyvy*�����<�g^N�W �"ߺ�9&���H�6z�~�iE��<W���oVV@]˓�S���cs%�/���ߜ�ܮ2V4�-3[P�>��\�g���M��nN�ƧQ���GY��
��
�k9Z�#���T欴����F�RZ]�S���k��Z5�Ci5����=��aHc�:���yb�y�o'x[�[x���UAG��&����*`e�߽���/O��S����#8T`Z�E@52Z�tx�~�����oT�qt�Y�K�}�3u�]� :����^=�����O�-�>}_O���x��Ȫaϫ��y�c^c+�����Zf���R����@[�1�$L�t,�E��@�X����2��~�����z){e0�ۇ�0�Ff�1���
38�
���
��Yg��L ����T����]�������9�+X�sw8Wf�� LNc9���РZ�9�]��-+���*?`���&s���1͆5���6=���"3@tz?iا��F���v>f,�r�d��M}S)���O����|���ӹg�I���#q� :A*P��AX�&m�f�]`�`���I�(�����^��ȼ}�?Rl&��n���m�й	��k%hg��4ь���F�'�"O�W�ݨ��+�~Ӳ�Z�� '�E12Zׅ0f��
	���0��DxگT0H�~�^��A�*��L�DPX�\�^�T����T�RJ}���cLZ���m�S���f#�&��lz=Q2F�c����$i _������jI]@������B���K�Q��u��YV@]���`Nk<b�:� I���4�Y2;$ #�y�,P�03�����o4 �R��@�JA�)	"�� ���=L�c�+(UlGPG�Z���>ȬC��.9 e~|�6�N�7�}N� u 8�#�8Y'��m���L����F�&��
@s�^k�>eԵp?˩f;P��=K�O��e"���l�>*�ƫ���HA� f|���}��q<Ui�����&p�
��z z�*!��&�a�ߎʂ�32��ޕҵ������'?��*e�T�N����Q�i�6�z�L����n {A�f�1|M�+���+�buV�}ղ�Z�D�(�Q��@�%,rd�0���Yԇai PԖ�����W},t��e�S4��#�c��Nu��Ã ��+Z����2Tk�&+Ƨ͸��ઈE5��TL'���v��m�y�z�}/`K���2�����q�ir �zXUf�[V�~�@�T|��h�򊨯ZV@������	L�k��a�zI��P�'�0T#���u>��d�5
��k�^�؞��C TX�s�h��v�J��O�}�ɋ>��Z�[ֻ�(�2c{���i؎Vo��(D�SV�V+�����J��*��ꔉq�;��AuQT~)S���w�%C�f:�6���^ky��Z�D�aQ0�����ab{�P	0Х&��� ��Ea0��jPu@Ы�1�99��~�*�J�g#���=Rd�������d@X�>L��^ݜ.JӺ]���ưN�h��Y��_��+�0S�t�D!��=�kݧ���U �R/��xq���b����
�߮���/e�;ܞL7�M��92 �u�Q�z�J��`��3�b�����	�*�=7�������H&�:�x>��9�>s<ʂ��o$P%�?�������~,�@�R��r�U{��܇�ɹz��E���aL�� �J��6$L,��>V������nY�g.�2B��?�^S�QHSv��#�� Jb=1у�U<UW	�����۲n#+�iw����Y+K݋�lT��t���!y��a��9�>�=��x1X��3�Q�80��MM�_���cF�mb�}�w�/b��c�.]�B�K�����jˬ[_=Id���|;�*��C]�u�
�?k�
�'���Y��Q4�(�򧴟���CuT_Tb�����h>
uU@1��W��(�H�%����>�u����p ���BDwڣ�R�^ҝZ}��:���� M`�ƻ� /��6,5�*'�[8j�PO��%K�e1١W�t"_��I`�%���.��#�����'�^A���
��r&S��	#�3Ճ���M����������\�9�ol|�&nT' �]�;+����'��A��8�ٿ�\��''꣆�	����F��M2��s�SWj&Y}�AY?���<	e� �~�Ć�"Ʋ���82H�w�����E��Sz�≡�9�N+��NY�g-O��njY�	"^N#�\���$�!�8�a0���
|2�Q��x*`nD��X�+e#����4�L�Y�2f���HH��[���Do�^ �aol�a���j ��L@8�> �q�4�Bn��ս�M��^���U�oj/u��Q�F1��'�8�'VWկ++���%?o�,�:̪���h��i�������Sa�c�cnY�k@M����(�@�O���vy������\
pe�:֬���f� FuIvy��0��Ԩ>�x����_[�]@F�B�R�-�/��P����>?���8��ꞥ�4!� �^���h�����n'F�}����hp��ak*���	�&�����>ki�
����Nr��_��}�1�k>�AY'{  >?	 r|� �-ؽ�xS	��p�,�	Os�5kz�4tp���r��r��Дx���*�j&S�&�l̐� ���ɋ�����v�s�S;h��D ��9j�*Wq����̵��j��Wb���21j�~��t?�S{���ty}�����U�fe٥ ��7���Ze��O*+�����c@��g��TFX����Y�`Qgq�#SQ7)=n���}����%"����	Q��X�$K�k�~�Y��3�k}�VZ�
�NPQ�;��X�W���دS3A���\�UJn���FV��%0����	�&�X/˾��`A�N�<�� 5�8�UY>����"�.��X5���f��r�bi����eԵ,���t|�j�q_�=����c��M���&X�ᜯ`ZԪn��z,�j��������+�Q�;��v{�W��>s����f�����q;	�b�g&��7��^�F���aC�6&=h E�̘|a!�w4�l����q������+��zӵ�\Yu-GXf�Q0����}���(!wib�(ْ(��%*�N��Pr��2�Ә��A�� �� �u$*�of�RJ�p�NQ� ��#�c��swY��H�/Ġ��TǤ���t��,s��vX�
��؍�t�R�6u�_��x�+׊�߶������@�O)\��yj��'}Cuf	v�Qu������O�Ы%^�7 V}7�X��w�^����t�=��"�3 �3v�5˾f����@8��~���$�_ �3���@�G5��<����(��Pw�i����n����35��y�q�y[xҘUN�VeԵ�,5���A�;��ߖ	z�h@J�Y������"�����>�q��a!��7��!u�f�,��f�Ϋ+�{Bl�<����p�&ɐO�ˆ�N:\� �����4w�����8Հ6�S\��Shg�6)���`[�ۘ#��0�@uk������Vl}��ZN���q��wџ�����0È�-,�A��PŵI���� 9�rT��.��T`�����ד�4�9���k�j�Pz�$������L�9��R���ަϟ?���/�V׵�TCӨ*�r��c�F-�K�Q�keF����H��c������>��
�C�E}[~�y�+��nYu-��`��>~���nM`c�6���{H���>]^\�w����Ǐ�N��ٌC�ܬ]j��V��U@�u��y9�+�z)Y�9I�Vr�v�(�7�v���.�����?�d`=��T�ڲn���;��(1���"�z&��v��d��&�3hCe MA0��$�	����X.̳ %j��VM���P���v���:�U0��&s��-�3�kj>�K��~�>M`����]@��;u�Z�0��KՔ ��VD,�jb��W��J7[] �Y��ڑ�܎(��/�>ML���*���wϠ��\�b��u��	#0�W���1�� �3��J�b��龓�`��A�c��X?�Z$⦝b�W)+����=*0����I�����9{K����s�!92�1?�?��/�����ҧ	��M ���]�%�ذ��{��kg~��f�A��EO�ܫ����sC�?����U����1��L��	`�'P%VJ@�ɬx��32r��ov�`-� ����D��Gne	� ����b1V�6JFO]�4�
�/ZV@]��3W�A-����F��]��K�5�U;�2}}9��O�" %y=����W���N@K�U��?쒪X�F���X�Պ�Pw���~�ji���1�ը�h��t�� ���2K=�������y��Z���b.]b�ww��N@�W4��^#�,�`VՉ~6^د�X��چ{_�R�^V@]˓J���6%�G0�@@��܌�j����?�g6�)���/����h:
K��Sā\�r��`ѺXڹ�<7���k@��� � @��(BE���r0%����;�����3�U���/_җ�M��QX!�Qb�UG�����7�@L��î���
�k��A�8rɦT��h0�G�cԳx22}x������0�n���-m���C Q�ya�ǳy�j���>�l�	��N�{�Q��='������g5P��E���,����������/�y;�#�z�Yu2�ʪ�D��P��q�Z�aq������������Z--;4�I��;Ď&������_>��������l�����?�;�B߫�ig,ѭ��k�����XfZ�����\c��xG+�X�����y$�|�.�M���[���gw��j�LSYWP:m|*�,�9�IV����
�kyva��A���g����=�ǿ���믿N`�^���Q@ S�z�{�������^������	rmS��a�t���_��c��� �[Rn�Nd��u�r�Ng��VV��eԵ<��(��f��Tt�M���@���w3��>L�)����`
 -&��7ʤr0�����0K ���l��5�p8C'�Y���+�(�7� ��{%�]�T�'uK�ٯbkU���Vd-/TV@]˳
'�`8ʒ�sԤΚI��x�����4��-�6b����"��1��_
�	a���ˉ��g��텄���L�3M��������s#O/˲�/+���YE��� n�zM�D�R�Zԭh��O��r�oލR}#g�3.����_KP�:����ID� 5�!�Ԧ�!Am�EuGPV]��)�Ϊ
���/��|}Yu-g��2��12��>��_\hb�1Sƭ��	'�3��^�z��^�%�Tƺ]�dݒ��MKA��TS�^\�bV���SUk��L��Z^�����g�����8y�c� ��E3�5�Mԗ�ʄ�9��o�N��>~�-����l��3��fw1�Q���3*�b�$�ww�@�Z��g�P������^ˋ�P��ҳ�~ga��E,ۙ�K���q�aj3�Yu�l9���MY82��*�Ю�9 ��VI@�ȗ���nnnd�BՍ"�ku������p���FYu-�*+���6 v�5[u���fqMa������0�#*� �c������^Q��H
���޽���?��$-Q̷����w��	<����lX�ox-�QV@]��:��R,�S����r��5>��Kiu��aJ���~�-���c��|d‵�U	��)k�9 �^� �D��ޞA\R�&0�lu�p����b�.6[[Rf՛�nYu-GJ͛\�T&4J^҃f��]ɡ�ܤ8����)�S��2|d���qx�s|}�L�U�.m��Q��=,�ਫo[^vE2s��4�J��Q�Xue;Lu�w/�W�/�$�'O	��������m?�7QV@�K����ϩ�Zg�w}(ńS�����d|!��t}}/ ��d�j��i�Z�I�\��o������ˀ����/]�pػ�D3E�骪��y�괝���P�O���Zib�K�vͱz�QH8j��1�w/+��e�1�OYP�|�P���.���3��$��G]ET+X��s�֗��&F����R�ѭ-���8�C�錴'N�M�d'@���~8p�n���jU�w��ny�� �U����2�OS�b�rnYu-M)�w�1%���e���ձR'ǧ7��@�]�G��W c��c�[���6[ ��v�J#�S
����EO4�w�
�!�
�k��`��H9nM��q��$�֤� �ܞ~����L2��`�	5�d,W=�Ǵ��_V@]��%lHݗcZ%�AX�D^j�z�%Jx_&*_ƛ�MN!��uԩOk��eԵ�J��z6����<=#�3P6Q� �#�ܲ��b�L���V�f�2ʮP��,��r>�͢']i��)+��EKT�	�*��ſZU����x6��j^���?cy���6�-=������b.Tk��)+���*�rѣ/�=^Ԭ����9�^��.2C�|���D)�>Z�oH;��5���t��Z��/+��%��O�������H�U\AU���y�ρ�W�8������ ��.��ujߢ~��<�N���*����Z�(=�R����{��T]�h����e��K���	e�49q>Y��U/#���QJZ�(+��%��^>�f~�) �g��-a?��	Q8R@@�T.���K���4�q�XF�Qu������7�0sn[!���P�R�*Yq�cb���MD~�������)(?���הe�_3��Q�/I�$$�'���1������Z�E������:�~�Ė�*'�;��,�G@5bK���U��^�J�q*�t���5IbiZ�g���bv�@\�;�+�u��5�
�kI� ��a�#X&Cj��=i��<ߗ�p�O�a��S7����}�"W����Ɇ*I
B٨�d)�W�>�U��k:e�#��e�!�g͉���8MH��?������1�QB�T8
�tӬ�%M�g��sr�1 m�tmVKky���ZB����V\�ޟqJ�&��ђǷ���ߥ���M[��:=H��O�E�+����4��Z�٧���;�.5&a���/��ۻ������U�h6F�҈ﯮ�����C.�Q_�����gЇI5FDl��$�Po��~��1a]O�H>=�E���5�r���?j1��X�Y�e	�����1j�~��'�����n� ^�Rٳ���<�D@�gs��T�Z[�S�mYu-�.4Xm	���j4!@�����/����{U$:�tq�d	 �蔱Q~O[�*�M����
Ƽ����)��a����s�׿����P�,�k�=by��M׫��h���ީ߶����g[;*�`@����"������-:�w,��c���
�?p���at�6̒��
1Qb��O�MH�7���6ݨ���#��3zc�wK���oRV@]˳�XĘ��:.��EJ�~�����	DiI����������΃LJ-kc=k�9
G�M���;1�>�Eh�م�'N�������ϟYM�T�� �IE�d�Pb��K�P[�������'ʏ<�����g�����72If�Q�SY��J�o�>�T*��I�puy�����XE�8�l��?��^�b��6��1�Ll������f$�qoT}2��8q��r;�<�* �Tz]T �!��u�
�kyV���TG��,H�DYұ�����ۋ-9}ާ�>�뉹r����?�طD�p��bL��"���p�`����g�����ݝ���(���RK�W���t�ky��S��$j<�^��X�d��2�n=I��w���~zu��yi�/7�׿��>}�ȫr^\\�Rǅ+z�L��
/���ӷ�[aϊ�N�vj��4��M��?������N��zg�0K�/�Y(G��&6Q�m/�ar���*��ɬU��疷4nj@�i�eU��������/�Nn@����@�6}��O1V]���֞�L��o%]k߉���.R���ŢɆ2�B{Nm�ۿ~K����͠J�I�
�)��e���
�9c9ѭ
�)c�����F;�^V@]�3����Q}(Ch*�N���n����N��ߥ/��ӻ�k��__]����һ����w�����ߜ���-�׹�OJ��� �������a�����F�|�)�3j�~��U0���/9'���=���Q�vY�(�!��7�����T;��YC�x�"�N�F��<"�&۲'{>�yx����<�F��0��IEa���Kf����˧O�Ç��g����Y 0>O��_��O.��0�(�e�:җ����������Lc�>�OV���,xMPȮ�ib�Su�>�����e4v*�W�.D���,��Hk,%m9�d�Y�;fy���7H�_PC��,����vé���J��Ի��W�4���}^���8*�'4u4���T���t�k㿙�N���O��*��mTv�Q>c}b��b�~����8[Rǋ��b_i7���~z�������K���[���;V���)��9�|�������Bg!�C�I�x�ډBI)�>1�/7_�����>�Ko���~��]Y;j��(י�c����v;MBW�ӧ_�I�C���ּ�F�V+Ћ=.�cT��O�鬛����q��p�:wdDپ!թ���2����縢̧�� ��K-������8��b��N<��I��R��|
u�C;��,��FBp�>�vNef�"�m!��Xr��˒pH	�Db��9��}7�GvP'������J/&�~��h���t��p�Ʃ.{�_�~��"� �Xv�xUR�j������S��:��g3��)g���9Kg�"���7�˗/���n(F���q:�����uY� �g6h��=�F	��tu}�>~���׿�=���_9���X?���(�?�����S{S��\jm������ ���I<߈�Wo���L��U��s�"4z@ ��@���ѷ��%z2+0����N-�^�L� p������U���j	��-1t��vKK��d#h���n�<Qo7%W�a�;?ed�8��PDI	C�$ȝ�[/.�	'f��/�;%q.A��'༘@�D���{v#���y�Olubg��_%�Y�5�]���6����g�C�"F>d���{I���w�N&֗�OߧɈ���ECmyr�	���[�]�V@�� 3�T����ԾW8�ي��|Y\��Ѯ=o���_�1JO-���޶ ���A'����tt��x���R;3���U����S�?�+�Y�+W,U��O��č8��7p��[u������7~|��A��l_+B��� ♁��1�K��4�qRp#�Q�ԩi@�tK �����Yw�NR�� �� ������_�6�����ω=�w�yֻjl:��(��2����.�劮7*S��>	"mN=�1��;;؟<0��N�Gq#@� �d�}�u/1��d�Ԏ���u�Id��&��Kn[ *M�^�~��ݥTCv/�F��h�:j:���������J�H����R�9����3ڱ�.�.��N:�N����i�^��I�"R$߹���
���Q��.�1�t
��p��\Y��%KY�@�t>�V�W�� ����X��Y��[�q�3�쳯���xQ{^L���I�><���
T	�4����	U ���}����T���|�T�	Ǡa�\{dT76Ą��! 3��ª9kTVJɶ%���x�R����$Hf����n�����.a)ӣk�$�6X+OgN E��3`�X;�>�'�R�5��Nz�<��Hi�OU����r�?, }`
#��_� o\��9��^�@���Iy@�Yf0P�b����yǏG�5y����+�\�s�\6@� V��ض��x�a}��:����H����ދF�q=���kre�28w?�'��4\��+�h��	H�w��Y����{)��wiV�:a�����[���Uyb�@霱)�I}j���&:]�$�����6��q���[GF�Sb@ꅹwj�g��`�k��K����9I��44�#�N�t�,5���#�DVZ�����5�=��c��GH���,���b"	���Ԍ�ţ�_��D���^j�e�Ҏ�]Y��ce^�q,�9�u��L�����BK�C- ��T�}����uD.N�E�E�TD��E�٨���Tuˤ&[}��<���o�W��30H��:+�'��'����5�p�T-ꐔ�{G�+Y\�Xt�2`O�l� ��f���ML V�3n&Pl��ܱ�	��TA�a�TW��j����̾�*9Y��ҡ��@����y�����̛(/���:�y���Cl`P @<�Ɖ�r:�3ƚW�.A�/~^bKK��F�_��T��C��zܑm%��}Yط�ޞa����8�|����/ׁ�Xerյ�a�c�c���E�/����R����a��R¬o��	<�Ȥ��}%��]ۑ\�R�)[;��ψA��V�� �*�^�7|��P__�'2�#1��r?ZÝOH�$b�lBxrc�|DG]���/X3�س���|V�ey1@E�!��l��'obW��h�o���#_�\�1�c�wv��>�T�m�`/2��Z��1��zC������&�����1�	�_��Q�5H`�ͺj�l���� �-"�Nܳ�����]���!���3��<�tA����F)���0#��1��I@R��z�M���1c�N�Af:�P�y����52Կ���;πG���1ql�G�.��%�J�q�nv��+�����/*�cq�)�d�ŵ.k���\���ŷ�*fb�.7<���Ͱ7E�D��k/t��G�d�'��稾�A�Vo�0�þ��ƄΗ'�z�%uGJ��O�*��{�p���۬KR�b�fpʝ�`(�����~�:�6���0Hv'����u{6��B�V���YH�卬��;{���S0~���z�����j��e��I���+��@=!��1�Wڥ0��������m�<໗�Tk
ի�c�0��Y�s��+߇q>�G�k]��":Μ��R����+��=��&�B��Ĕ\�D�-#������ ��u�ڛ���������Z<.2V����1W�x[(Ě���٩�� ��E�3V�pP=���v�T hT��*��k���%�/��\4+-H�P�Z�ɥa��d}z��:�Q:��"�9���u-#EI�3�d��c�?�y��Q���硄�v���K��Xz������P��j)�Qt�\R�(貦~��GQ	�dl�1t�J��Ԓf@cU�W;8��V�L1�DT',��D�Z��l�GJ��Ei�5���%2��銁�ٰT]mS��i�"J$�)̔\���W��&�7�0YCTY�J����@f�#IAَ�@���JT15�EW��*F"84"|d�&�4�(���ˋ>J�)4{��E���m�>�1�)�O�i����;j��RUÁ�I��f�=��>�0j+�����U��r��E�E�P�ndP1K�^siZg�
�480� �Ć�f����[�x���-͜y@��u,uL�f�#�w��B���o'�՜v�zv�MK:�xYc�%N�\a���6��^�:�QYc������'�ր*��%�'^�u.��Z���Z	�(�J?��L�}"����	�f<�O˽i?���`�� �uס\��6w�>@v�O�'*��� -��ȟZj#W8G�� �-�]��::��N���RyQ@��!sg$�|��"l����e�ΒC�l���f`��yE����g��<Х-%���,c?����q��!�tq��3�~��p��ejev\	2�rr7�VuPлFܿ�J����7~��:a����3�O��������[`�Z�3�d�H��v���I�~��x�ݜ�J���
�biu/�$$-������g�ɟ]Q@���K\
	��&����$E>�q�¾~�%lu���D%�8��*���%šw�A9[��QTꞻ��u��nd"��Ȝ�a$�cy��	b�h�V����-��Y��_�2X'���%t��� �4�`�i�$'M�G�[9ׇ1��e�5tXڿ�~�2�����Ъ����ĦP���xn�s� �ܕV�A��;7�`b��0$�Ʉc�*|+��+*=�J��� 5�~��C��&� �a,8OP�t�3�59�4fێt�v�sT�D��h��N��A�#�J�(k=l���97�U�@�,p�j��)���ⓗ�9C����c�	.�D�6(ĝa�ib��������#��>�B�:e�����*�ޔ��\���A;���E$K��6nu�K�qڧ k�qm�!��ӛ���<�euLa+�	�<��tT8��&b9d������D�B�J2v���ı�:d	X�&�>�?����Ʊ�-�OJu?��Z�v���l#kT���C?̼�(6;�/v6;U�^OX���T��{�E�!<}�|�:밦�1�9��3��0l9��Y$֝*(V���ƅ#EX��$�".��.���^���z�5�3�)Fu�ȥŪGJ��?c��,�Pf����������Y-f��ji���NU����.}�h��9��J% ,�I��R�L1&A����ڤ��z��Vf׋�`'��T��7UEu]�y�J�3�?� x��/��k���UW0NX�x�yS8fh�{�����Z&�(�QQY��M����=؃c�qx~{o���֓b��i���Qvvx�52:#�̐����U؈�z��Pq3�.�rn��.T̠��_�l��e�b@�װ��~z��r�9py#7�R�x-����@q
PS��L��@)�
�RԨ΀��d���`�hñ��ز��Ȯ#&f�h\����m[�K����:ɽE7��ڗz�v�c3~x������Ȧ0!`��Zo�7�5`ܭA/2��>��6�ЊU����aJ�]�[ĵI�����P��<tϷ�/��s�E��0�\���%)�����0�U$&i���Q\)�����2Z���" m-�fU��}cG�iZ ]pW,���\c��Ů��@��Nc�ǧ\u�Ȏ�D�ܴ�P& s�yjo.~�v"C�{�I��<�#,�0B���=W�F�n��ߍ�Z�
/��a�Uv*��U��Ǚ'�7Pm2�ve�����u�^|ib;��i��k%n��	�Ŗ&�F���O�F�ؚ�����CP���!b,ٖݡ��!� έ;@7J:�T{	|��:	��@4��aS�?3�A"�x�$l�b6�Z&���	�������R���9ӏ�"yj0��Sx֔a9'h-���!CՓ'i�z5��S�sZ:�ߓ3:��_��=8��h~ן���Tgt�{k�%�}�q�,J��4�/.@n$$ת�V����NA��݃�mۏ�D�HT��<U�r��~F<��y�7J81�g��Śq�MO�U�f�gL��y&����wl�G�����O�y���@:*�w˾r���f0�8����i����e�P�OI�1��N�I@G��ҩ�;y�����Yg�.���a�`T(VQZ�^���A�=OdKRe�L�x�e��n5�+�Y�k�t���Q�-� Z긕�"f=�gc��ߖ���a�S���`z���	O���8��x�����B��r)��5B8�ee��|YC�0�g_�7��%� L�xfG�<G۽�V2���.�ٺ��.S7¯��@�k��Z�4C8|�2\�E�pb�4!&�F�4��F��g��ߤ|5���):H0Ń�O$�ګC�����T������e�I�x���:( sS�$0�
���n�Y7��8�� zUѱM���Bu�z�,Z��~�����6"֢.t�U=���y��B���k����RW��p��"�*��6�>aǥW���+�v���~z�>3���@��>l�j�(2�@Ҥ1c�s�Y����:�����2Q�%�����CZ@�zKX�lq�ȈӼ}t��m�*w�S�j�>��������ƖT��R^\�g����.�G:jC��^40���K�I�IJ3�V���$'���_2}	K����������� ��ʒG���=G��ZGAbq���L߫m�t��3W��Nv��G�]�CտEXZ����G�/�r�8��B0J�>���>��U��L�;^�	҄��]ib�~â?9�[�Wq�S2Ј5ok�%ֳi��0���W��%��z��\���'c���. ���xȚOKU�l֯:~~�`�Kg��d�����<�*����A�s�{Z��+=&�1��ɹoI��xnէuj}�n�@��i���E�p#`BU#���I��(Ɵ��A�mJG���ޞ`_Ǻ����i�u;y
� �P1�y=�2" =��z�sPe����Iq�G$ 3��A ]C)����~�KP[��rw����`���Ae�Y�k�j�x+0�=h?�/_1�q�\��ЎK�ij��U}V���&|��J��_�������ұJ�X,�֚y1H��R��F|(�!�����o�T�H�����(������ˢ�=(��G~�"�[?W�BkŴR�����ٮ1(��Ϭ�H�����2K�|l�X9s_A�-9�PN�0�8x�}�2�>Z��+=�2������ o��-�@��sn]/9��V��&o�a�QZ��֮���c�0�s�i��*�������=[}XdWi3��H'�t,�p䙟�R��?�f[I6����C�_Gn��c]�r���G����.d��D�0�Uq�:X]�%O�J��Y���+���o���wؗg�yd�̗P � h�� ӂ�#��Ig>���EQ�~�$:�]�����M�����_��߶�6Z�8�Da�nd����E�WUf ^�!������CCsZ�w͘�\����+Ku�V�����H��W��u�z*�:�rݮ������b� ��$U�4���8�glمʏ�V�lr�2�o1|x6����pK0Yg,e�!|l�?Tq�������Íu�b�_5��=ZC�V0�0Ք�M�3�LXT9kNd<)L��#
��<�rՌ�ab���8����L��N��"�P��ZG~	�|�R�F�L)>��Z<9�=����(�(������+u���,`�5$�͹�d�P�ZJ�:�������"R�e�+��Ѵ�}@��:��K$A�am]"B�u� B=0�yN=_�-�1v�"��D�k��Ɩ��6�n/�;���E�h�Q^I�K��k�;H���t�]6 X�O���S�S���Xfl�c�H��n���=�����b�g^F&c�YMP� Q��yT���fnP:eU'-�;ة�.g�L�z���$,!-}[l2d��~L
�Ơ�B�x����:f즶w)�bT���n�y���yZ,����Dm�oZ�����E�N₇N��lܠ�j��4d�T�m�}���[�<8��A�z��q>k��js�|%�������� �4yb� ����+^����f��� ���N2�嶽rʆ$94��;�<zL|V,�&]>�����E�J�W���X�3�W}Xo�<�s��ļ�	B�'��
i`�����1	�����W��OGx0��,�nNf����˞���Lr+�F�L,���]dr�	���+�̉Z�P�& uum0D�! m�e����<g8�[~D�<�,�^Ȫ�)�x���2�^]_ْ��Z�����7Kf��:�(f�9�����[�Η}"_b�KZ�g�܌$om�:C��I?�?�߾�N�0r��ʸ���.�#C��ߵ��+��4�T�'ХY�"\
�u2#���]���M777lp��d�%��Xa�����ѻ����[k&x�)��"���"p�K�F�4|2�J��r�9?�������#/��/z������xz�p߽7���,���ޥ�������X��u;�wf�z�#,�:�\��%�k�}�K��	>�� �4�O���5-�Y���Mw��[/�����L&�ƫ���{(C�Y^P##�34�x�ۗ6���$GxxxH7�`���?T	 �}4Ηz�.�5�@t��@�Y�'��I/���R��>�0�g"ѷ ��QX�#\�V�~L)�a�/|�9�qӛ>���{�C�܏�ՖUn�1����hr��=z/��W+�s=��Z�/+I�,��#z.����s�@ ����5�|ʽǱ��g���x��BWP��4���2nDh� ��R�-�b9]P���/_���F�D~�q��~�u�N���D��3�a�P��D���k���m�����ׅ>��=P�ds�A���S�i5J1A�5@m%�;��I�!0ݫS�K�Kꉐ�E0�ܼ���'o�b���=E��Xl��eM��È��Aк�&S����r�ֶ����W�_-��1�tQL}�lح�oR���o5<wG�F�F��`��]g: ��I@J�h$���!��%�*��P�ak�k��a��#W���"�֚%$�tN�٠�_��Gˏ#�~���	 "[�Ҥzq)z��v���COYo���+H�-��W�s����o)��%��z� ������(sO�B�%��m�`��z�w�}�Ep0���}�]�o'̷^^P��a6G�X�H�4_��4�_י
�X'��I��1X��Aj�7i�b�E�����|��AZ�UK}�ӓ�3:ӷa�g�Ο�i�sp�gO����R�#�i��qTGF�HP���>�LsAy����=���m,���۹m��<b~�K
���ā�V۲��
+�\��Z&�׿������RS�)�7Z^	Pk񽠃B��E>�*Gꇅ�zU��N`J/b&P�\��W�6��uᅙ��o��=ٯ�&kR�cSƷЉ�=��%��>��K5·��D����H4M�S�h� ��/z�V�m�S�n�o�\	��KJ)?������)��d��v��]jGXѳ�v��(��\{;$�H��k��cSj}yQo���6|��Z�]g��>�h@㳦O���Ld��AA:2z���RI�'Cd��+;��-$��`�(�rhڃ͞��( ƙ�"�٘���V�z�{n9���^���j�Ƨ=3S]B9H;��X.p|�Ν��k���L�*�M���������9��9�'0�Zǚ0�*V�����G�63J�ȟ�1=;\̏#��˷u���kP$����;z1��;[e$Ѓ� ��pq�ۋ��$�$�H��<x
������gx��cS����+o&ϴI}�@)���1�_�������U���3����J=Ѿ9���F�9��9=
����]��R|z _4nW��U]��ŝ�R���G�[J����J�������O.��;���t����k򵋺`TBH����~N0M�dz���֙kY���0�	��K%�>u��hb���R�7O,���)3<�~��-�tT�N̔b�1!��G����T�篪�p3a=�C=�)���)�OX1�@�Dz�	W���U����}�3W���=�Q�+P1,��gi����і�3�ŒF#��egO.�/v^9<���z�}��M$���A�8?*Ysa�E.Ƹ�4= 
U%� ~��S	�GY�%��t�
@��}��;�Z�?>�� ��c��{Y�M<N���\���d�l�R��`|���y�`�BES\�CN=D�K���>�6�g''���dv��~-�urX��/��ҋ�/�S\�o���&?LqP��2��5|61g�G�6�~�D	����i�~_(`���0Tnw����Dz�%�:4z��>Z�T�(b�m:5�~V0X��S��F���@#Y�S�c����n���Ae��%'��9�?��4��D9bx���!1=6���H?A� R쁅�*�v�.�(����L�p��zۥ,���+i]�.�>�V�Y����!qK݄:�u}��@z�.n�r܈���= 42�ri3V�-��o�C}�R�r��ܿ����@�Y�F˘%� ���,a�~N m��&��_~/�ԏP^]/'�%��#%1�k�i�G۽������T0��@'���S#eأ�LL��  @�����}!��י��Nc��h��Z��,��R��*\����Bg�Ԓ�]}�5���B�n���l����_������������
�?��⓸55�FX�JN��?����Ӛ����F���gc��?I?b��g�_'�d}���Z�c �?����yY8ƪը�$w��l�G��.��J�����6b�QO�3��bے�������,�P��l�d�ʪ7���
L�/�.�}ʑ� Lt�)��X�1C@��t�K���@�'u�h�,�����[^���{L��%�窶�X���J���U3�㾩��1����:���
�E ����c������i4tp�k`��N5Xx����VE>�d�ҳ�r_Ͱ�e�(��-��HQ�*�G�	:� �w�5�fj��6 K^�no�^������1��*6VEA}ͣ:��?F0爥m�T����@����>>�ϒo�O���(/�P]��6cs�MӳX�gL��b27'������M,u�~����=e7�~S�R�dY`��}5��0�k$�5�����8�ˢܿ>��4>a��������Q{�#"?B�cݾ�,��0������+	�H���g����F�֡�W�������j ���J��e��RZO�BL�Б�l���$�/�������ʱ��O=�����
��翻�*;u��$)N	��Q��|�W��ȿ���Q����8��oE}�3�Ғm�g��S^PӞJy�d���g��K�G�a+��K�`U�p�ol�s&���ĵ���~n �~����=��A-3�����3 ���X��;��
9 X�P����V�:-��H�Ρ(��o����DQ��K��a���!����X��/�	���m50T���z'���� ��1�XT[�l�7;�w�z�~d����"3�`\h��|Yv�[�ZX.����V�z6�>Z�X��4��!�x�t4��2n+�,꣼�c4F5�)��#�\�~�R�M������5��f��&/�"�zf2���b"U+�G~\��^�0�����m��+�\�F�O־b���f&�/a���Y�yb�K��ۋ�U�������iN���͗�(�'����ﳨ�3IC�|�(��y�K����0�^Nb�ks�����$yȒ��꠫�R|>]�3d��~�T	�ru���Z+AKP��"�&�dm��z�B����'����'H��-�WQ��{X��O�\�'���z|����]ߚ���:��-4���j��n��8���j<[IFm���=ӳ���җ½�x;�3֣������לZ5��_�$=���&Ss�֐�f�Rr�lE\#3]f�U�ٱ����m��}X�8�������o�_L�/����K8[�}CF��:�
c�X�����{�Dҳ�~E2�K�j���.%/���fp�����qH�"�x.Id��C.XS5�юY@���Sr��yL�b �����#�j�-��$΄s���b	����+O�Fot�q'� �?귣e�.a�������I	�t{�uIU�������fle���^��Eqd���x�U�.�{X�A9�L,��AG8Ez�@�=	��P�M'�Ғ�wdB�;�S�[�t'��h�:[_�	��z�ԅa�[]���;:A�!����	�DD���96��y�d��<�^$�m���+zfo����C�X��8yHHH!�+�rWEX�vƜ��o�l9-ufOYO��%��ӘI,$p����+�"��̞��	:��v�r~GΚx�I��'�}Z��d�K�r�߳e��DPѶ��js���R����KEX���G� ���8� o�����Pbg�,�(��^�γ=�$��O&�φà˭'I�S�ֱX㩀��,�0wg�9��p����&����G&�����^`� ��C��=}Bѱ�,s �%N�l%���$��vL��M�� ���b���X��o�
��f�Q�I���z�L�~��'��:��̬��9L�9ko�#^;�-���� �۔-�o�77:S��� ���?vj�3]`�2O�I������Q�L��� �g���K�ԽUrX�Wj�)�c���Y�j��~.�;�9+0V����U0��F�y�A���|H�I �� ���6e��\:d������W$�^j)�lfnD��̸�˜�.z��{I><v�8 ҉��ن�X$�(g�8f�r X��6��J�P�bͶ:�U��)����G����0N0��w��J�oP/����K�5�?���m�e)ȡ����GYlG�V��XԩD����ʈ�!qE�ZA=�mu����&��L������̥��N=�
T��8}�����ꏭ�����-����I7���	�E�y(�u��!�:��@��ʬV��tK�R����c7:Wڥ��w���l�!tؔl���X���(fS�+�Ӑ���`I�� Ԩ�3���u��}ϊK�sp�~oI��v����`y���_[0)�� e�����������ig�9�xo�� M��2�ј��H�0�D�%�[��5N�xN�`��7��~�dʈ�<�đ��R,X�5�k����&�/����܈�GChZP�S
v}K��s�����˘QDU��Y�b�_;�f�'��=�$'�#�ǃ|&��W`���D9ee�c?��d�;�nܹH^t͡�l$�O��-���3�AA������td3��^��n︇�Qn�aĤ�8'�!�����p��9�,�z\��xZ�=�,|-���V2C
���оᜦ��dV\Uà]���I�AӫD`�?t�Rע�0J+#��AW��G&}�'w�k����ЖJ$��%���DD�\�X*ʹ^��'�:p��A�Z�KL5��QX����c��a�A'7՝��V`0�����+����� Q]���::��* .(�IE�biV���f3�~�j
8R�?Y)����ti�^\�Pe|��Ҷ!���\�^rg5�gm#�]��`�1��N�&�r,�y��0q��7�7U�ܐ]�?w�x\`�-s��9'$w���"��}��Ṅ�A%Zی�0�g'�
��X��j5��W��x�t�$v'��Qnhޱb�%<��4��e��ζ��#�Z|�F���)�Ⱦ��vVyq@��s��ݵA��G`�+��X0hM��V�}�}wq �8N����o�$��P�O�Y�H`�c����Nv�P�H�����N�R�y8���C�|~UW``��v���"0ڶ��]�q��i9��i���1o �� ��u�_�#\b��._w4i�J��4%kK��Qg^�֐]����D����ƨ<d8�>|�$<����cPQ��k��,X��������T�� ��������(�	���RO�j{n0V�H�g�e���Q?Vy}��ߘ��C_�lR��E��5R�R=����(��5xܨ��˦S-bl�ԧ~�E�Q�Ww����nzN���V_\�
�r��\�X'���z�:�( t�~d6�DM~�T�POf��� �%���6��v��d9�;�3�6Q/BI��Ɓ��W����X@M�u�i5�o���L0fE۩D�_Ä%��w4�C�n�v8�:���#Ť���G�:St�B*�X�����DǓ*�+k���]�Y�8@�$�4�J ͥ����Mn��1P�{�����~{��&O//�����J���W1���/�HU��L�י�t��iz
MX% � �xE����]�h`�a��FW��?-U�|N��j+Ǉ݃ �AfXQ ,@��������[ln�"k�C����B�L���to!���9��^�ʝ���p>Z��@ld�ո��*WRq�$Yjl>9ó�dI�;�����;�2Ք��=k�)�]:�9���
���>�����A7'������)�i��UQ��n7[/*�q����J�tp���B3��K26տby����80;7d�p�/�M��}�+wqzg��U>�<�9Fs[I֑��c�uT���q�T@��-1u��U@UTX�2^�U7+m�L3�y�)ݧ6NQ��Daj��躑Œ�b�Ds��k>Y�ze ����)+�.����������A�����a�𼸽;�B�*q �K���8%Lx��f�L���`��|����u��0�N��L���ܿ������zc�����<�2�d|��h�%Q?=��`�J:T�����
��R�o�`ا�EWh�dƦN}��	G@%v:5� o覊8�c�lƍ�	P0"0ݲHݱG�ݞ3���uPX]�C4d�=�}�LMA�L���I�X��t�Ӣ�qyq�{4��+nQ#^��ۗ���01�VWȤ �bt��`ME�{�Ԗ߉��<��ǼT�1��Z*2�/y��=:�}�$���tw�(t�`�Q��'�A�SX�}��uʌ�Z7V�h�%zI�!��QV�c���ȒY����h��vA�Q�O/ ߹�&*��Bфgb���� Ǜ+/�w�A�.f}c����i	�(l>uuP����W�d�zƤ��yk@�Cnl�/�T.0a�����:X\�A������	��.jBPG�W5Viup��`Ԩ}k��̪��k0��2A�=7�'fS����{խ��?��Km�e���Gz¹���I��J�R�T�TIG�%%O���Jm���X,fM^I����%zA�Mm��c�� �@T����-��)���XS���K�˳��z` E65�74��Y�dU����J��{�������ҍ�-��3�]�dKi�Z��=;�d��A���~H���r��$!�t��DQ2�!��7����e�pR6]PJXT8��lLQq���̌����. �>du|�.�%:$(�!�C�Δ�)��l�b��I�,T�ӕ��S2��:֤�υ���DDG� kXu�H��fu�zw	������ Y:�:�'��vP���<������J���Uc_./ޱ�:B�~�F���C���{)���f��(��bn�ܹ�����ý�"K1`��E��p��&�UuP_є�!)��f 8z���$��V����LGN�C�Az5F�z�z*�E̚�4����$�:\�lb@{��0���@�g�����)�\�b`���=��X��;���˽��}BO��-�0�%��2
�7'�r�Lm��v�# �ؒ��̠g_�'�e�ܛH���W�g��:��6�������aM��i�6 TFZ�XƪR?l/dI�i������G�[Ӆ�d��A-҇}�����խ/�"�2�}���A�͕ 6�qlE���oJ[��|Xw�[34���4�:��X��H��cm�?g�F��t��+C��ɕ@[��N����X��W�©/��db����vȀ?w�ۊaj�{�����OV\��uc �� ��Z*��S��,�{�*+>Y��)"��/�	P��X���4���`��#ú�D��YX�J��elā�-����pD=�m���Y8�� ��0T�s��A"�Lٖa��	 ���=K����PV��] [�BD$c��6���W�u�n&�,&&ºMgК����T��Rq�٭��~?��Ĥ�$̍���EϞ�:90Ҥ�e�Y��u���Iw�/�4�Vtj[�{����.\�,`@�#龻F7� �]Q߈E���RU3��(ZRl��F/�+���Ґ��W�jd��MP%p������p��p-US� �9x~�1�m���PAĊ'���(�=�Y)eq]2N ��	v �e��n5�#����$��$�1�J�X��F!�B	 e&����*�������5q�z�ሀ5x�!����t���_DՙVM�`�ES�mi��1��x�:U�cuw��X �>�%�S4|�� ����D�Jϐ�a�`�M��'Zu�c`T1�c󃻜L�{�������c�Z�B2�����'r�V���t=��"��
@���Fm//��O��&z:߀�d��lL��-����l���(PA�������S�}!�w����l��j7+�|L��#��(�SQ�=D~���8*3X��Š8ͶC�dz+Vpg�퓊��C�H_�|�@�΍D��\����X�R�n�G�8ۈ`���T431��]�"D͢�C�N~�u@b��:s&�1�ؾ�ќY�4�H�%F.�:	�'��@`Á��`��h+� �(��hYL|V_��
�~}^$��?�{�� �����oLO~���v
���P�_���wPo��zw�7v���M'0	�"�;TY-�����,�<iJH4�8..��|�V��t>�汸�*�n�R�B�KrۄD@(�j	l�"$k�L��óH�Т��T_n���S�3��d�@U��e0���3e��avfw��w=)��<�`� ��Mt�� 08�P@��`@Sp�`9
��@����l�R�A���P?F�\��+Wu�	�`��%�,�O�D�p䗊rp�A�eL<�2���@F@?�26��d�io��j���$��&؇�N�
|Ⱥ����QR���
 �)��S����;>��B���-b���Y<@F�Xu�zIdZ+I&f�H��Aԟ9�.Q��)�$����t5�'�F��;�O}v L���Fb�cɑ�B��d»��Xj���P�{3VZ��ox�~r�~�Z�/Y�t.a)Jy���`GN���cD��ˠ���͍��SGﴓ��Pr��Da;Ӎ�c}6���
�������r�tM*"ډyJ�*��K��~�
�b�ss�˔D/#�e�|4���>7��(�zU�A���� 
JZG�W���-Y&g�V �j�%\t��H )��ϋ����Jw�YL�^�0�����d:V�����n;����DB@I�;<bF�D�9Eܦ��l# �wʼ�J7�%�J��f�:��)}���[�<g�"׸`��5u�$X՗u��xŀ���% �&BZ� E ��T?IЫ����7-ߑ���������&�����n�����6H'����E��`���0.:����������0�}������A��-����bp��"��� �ҭxݜ�$vw�B�b�����D��M�f�;ҽ�9h��Fk7Ĭ/����K���|�1��1��%	��;*3*oQU]�	M�ӄ���hR��ѽ,M��5�{��a����u���K��ɑ\��y�O1���ܛ��PwXt#k�j݇�j�j&�2=�)�%"��jHOp]q�HV���t���>��˧���{���	,�b�!TŁgMҝD v�~��|�R����4>17��#G�~'@-�nQ`z��c.}̎�����6،��(8�� 4Y��흊nce�Ȇ�k"��i�-�٘/�f�.�%���-�.2t���	�݃���Z����t�U���3��p�uΖ���t�"�o���IPp�2�W�,��ى�4{�#TқT���*e�Z���Bi�=Sa��à>��S	�T�gD��)?��]���4!��9ݐޝ��C�1ۤ+IvR�ܾ�5Z�ɜ��\T�ߨ�J�e����U�'Vg�!��N��:�ߦ[c�t/>ާ��w��΃P�)�~��s-�&v�NH#y-^A?j�W��+Bt�T}������N}@̌�49�V��6O�^��f�l����YwV�H	1?�a·���)��F�,�����K�=l6˻���	���{'S�K�#�suy��$�_����6�I�򜲉���)TW�Th*fhto+t�������d9�zmL����:[������5�`{{�
�yD�{�RD<�H��˜�?�y>�܀�����_&0�¾��6z���M.%�O)�,� 5E��S�^�����A�Bo��쫨���%{@���@3�3��{�\��?}���%���O!	K�4P��Q�%	�.}W��%��X,�Mk}��˫jyl[`��>M�K��f�5�UAe7=|X<	L?�@�[�'!#t^��72` ���f/b.��v�řKR]�-��|f�kO�u��
N�2̂4``T�d��_��E�c����<��O���|﷢���A�>��ED����u!96R���j�3�7�W�8�:%؂�o��W���T��MY��{�%>�[��%`c�(6vgz��s&W*�R�a�"}�n���  ���	�=S�aU:I*�'P�ܥ�|��D�M�/?�i-�(��h�7]�/�tщ��	��n���d�OWWW���;��������1�C%d^ꂅ�h��PV7X����?��h,��U���YWbl5����苓e�Ec�\�^F,��$����]E�0ѝ�!À��� ����U!Y9#�w�;����V�L�8 ꢌ��h�Fź8��!o�e�/���tkC�	�7��Y�h�\]yj�K(W��ݻk�1�A�j
M� B#�樖澟긕��R�idU�͏�幰e��c欹� Rt�w{�s)�T�jA�oʢ����!���"��Y_��՘Wd0֕�ޛO(:�?�ްh���F��s�s�3�x�ߘ��DX:KXh�Ɂ	��e��u!�	Шm�y>��s��OO�}���[��K�8��f�>�$���n�G�T���G��S0�]9  8�S��ջ�,�� �P�_�i�L�ڇN}�s�1!���L�.�hˁ�IV!E��+5P�y�&=1�ۙ��b��Q��]B��"u\�����;��i"Xl7�`D�z����_��F�,1�+uwb�%��~��j jݫ�%��s�ԉ)1{�Xt����v�	f�{�����qT6L�A�WW���*�M��o��*�29���Z�{5(���~��*>ݖ��n�cƨ�,�_��q2(���D��+�Zn���R\�h��Ơ�	��F����&��ǟ|<;ū��������]��E����������'6J!l�:��
��'DQ��lE_NR��/����X�i�E��	�`��$-M��p��$�h�>�و����Fa���|�����1IMt��3�0�{z�U�/���!�g�۝�X��ؽJr�{�o��W�*_�ڸ6Ɗ	���M��D丠�Cm?1��-b�"�Z?g�^mk���ŵw3% ��*hRq���r*��;%B��<��uF�ل��4m� ����!Ys�E�f�-���o������{�_��#�a,֖#^�������W	���2�V�K���MfF�rP$���;�P������Fگg�:7n��]:�75)�I���S.g��j�g�|����% 5�� �ٻ��S�ygɐ(�樽�։�y�ό�>��?�g��b��/���>O��X)D}�\��o�^%��ͧsnU�b�ʔ}�gz�������L�B��K��8R�����8���ACW�86Ց���������\B�j���$(���A�]�`�W���V���؝�a0~��^)���;�uauUӳ.�_e���Y���-����e�a�� X���Rt��?$�E,��NU�wVZ�誸
�D�h�~��:r������@��ff���#�$�~�z4��x��R��g],tT�gm�
_>��_$w�.ʩ�������;.��+�ƅ2�}H��.Y]�Kc�(MƟG���oI�������!~��ݠ�M�P�,e�d+4X��|hl��'�"Y�0ܝ<� 	�������dH����D�������٦D_Nm��7�jh���BWt���2 U���NP1�Ө*�=�>��&b�f*��x��]� �w�w���܃��MmMR
Y��
R���ܪ�w���w�z�'O����B�lT�a�rޢ��HO[),y���x�jp��]k�.�&ˋj�ϰQĿ���n��c�4 �^C=�ɳݛ��tk�Q��V]��U��7�)1PIr3�6�@:Y����d�%��#r�M��P��)S2�l5���'[��N��T"q� �D�AAO�	Fv�N��".�d�� s̫Qr�)d�\nؗ��:T��,�	����3ǜg�O���:J��I��3�3J��U�Z)����(*��NnH�/
ҁ�{�=�K7�_����������'�	�(S�A��e2ݚ[���M�% #���2��U��QjR׃��ˌ�c�E�!�ԽK�&0%'}z�u�8���z�ޒ~w�����,�c  /�C(2�Q��{�n:��Lз�"�h=�_�_Ӌg�4��3��5[��今��q�Q���*:�����e�v�jd��������%������+�2��4PF���;h���^�FD�ܫ���z�^@��ڙ)����˗"�,�3Q�
��1i��U���ģ�-���AL��2��v��S���U�Ttu���ԉ�߅�
�I#���Y�{Sd�N̆���
D iY�\T�\��xœ�����E���������W�c���i�8�m������)��FA��)�D�����&'cz�mQ�sv_Y�a�4���/6�G��t�>~J_���������4�X�d�^!}�IX�
��/%3ը�|P7:���m'�/�J�4��rY���>�l�<�q.������bS������*�臚>�oϙm '㛇�3G�t�f(b��h�ׄ(�+�Gǐ�D>�IЫލ�'&CL�~���8HV"2!	�_��fы"��P��\���>�e�U_Ń��u�<�ۡ����D@���Y�'�&x+�M����B#h�������V���ʢ�vҮ;h�eo,�CV��O�7]:L�S�A�Q�"LU���Z��� �~��=�ʴ�C���-\�ڂ,����?��Dz��ӳ�B z��l��P!�$�1�;���D�/"����{5�D����B;�3�(d�4H;��&p'6�˧_������?uB�i�>TE� l8٤ϓ�A<UHj���;1�>��\D��yc5,6z����������d<4PU{��ިu���G��Io����2Ҹ�Б�F��5\ܛCs{*`"�V�®�x��9ZDf_X�hPYRh�}�XJ�14�����d��4�9���>}���]���4�T|��˨���{[�^�9�ʕq�ǽZtK�)�ؖ&�N<�H$�	����d�[q��������A\fh�^YQ�:� s���ɢ3�U�������N�>�e0�_���d�H0���
چC�b�ih0M<������I��c�@Y"��QRn5i���~���xn;������ƈ$'��0�':��%��/��p����G��\�������3%�J�:����I���*]7��D�'�&��'ѭ2�>��QU��0��������QX�C�L�pQ�F ����"8:}�����ޛ��m$I� 2��M����ε�ξ������RK)�ue&s7�dդ�R���J��@Dx�����U?�~1w�+��14LCe=&s�Ci8'C�.�"4�ԩ���pO>�D������B@x!w��5�	�f���k�z�j�mGo�+�£I1�j�����R~���45)f��czƖ,C�z�׫�vܱ�Em	��Ò�1	 R�(��2��К�:����P=�c�	�����Q^X��'z���X��3%
Q�3�_�}��x�m0k�#ن#���
x��캨�/�37�h7�*�b�$h���%E���CՇ�<��4�6�mU`��{��5����Źk9����=�Z��P�)����b~b�s��y���.�?K���f�5daJ�(ZU�g/���Μ�`�S)}v�'NJ�k.�:��gx�ue->�C-a��$�d�	(��0��z>�.�W>�̴��M���z�6>c�ׂp�8�.x{�x(�;�V�y��lrm��S7�Z�e+�N!��TjQ��ޑ�<wk��E�1���9�5r��p�B��v��z&X�Yt�`�!M=�ߔ����J5���0��h�mn2�8�l,Ww؏sm�W=EL���D�$g�����F�Ң�g?���>}:{�o���@g�p��lH�ObSR"&]������**�0�d��2���\�ʒCAT7Z���G?��n��E����5��K�,� ��M.��� ���,�?=}����콙���Y�T��a�u�8LZ	M�?s~�'��ĄJ1�3�󴧟���!7�����S;&60&�$�����S&�0���i��;�[;g��s/@r`^`��~FU��9�G(�cK���hG����	W�h�])�j˒H��B8�cT�,��>��3�G��Nc��`�|&�������ݍ.plXJ'[+��qmj�y�8��u�J���7o�ۻJ��A�������4�<2�O+%1:q�aG����L/=cO����~xf�)��'�eW �W
�zL1g)r����Z	w�{,�^��&��STIR�)�v�/]X�IF����u`�7jU\m/eQ�:[�k�9��}ǌ:�ʁ���V��xޏ�\�|��v�B�a�&��'Ǵ@�n�(��_٠:z�s���;�z2�E"*�p@�t^T+N���fˊ���:��|T9��o֌�l���ZU3�� ל�d��e�n;N�c��w�3��v++
 �:`G.Z��I�JL�!	6/`�'��kڱ���V�k1��F��t���������o�T��A�".�aR[�^�Xc8L���C�p)������]1��X�WՏ�8dt�����0$H�a�y��y���熛�9४q�&t ���k�GG�<����Ј����`���t�#y��|�G��J3��G@�c�'���T��2aA.;&U���gaޕ���\k>o�Ã��1šb�<:E�HG��ð�M��{���8T�@mf���?蟧��ǯgPe�~.���Hub��}��Co!���P ��P'�i��s)�����ߧ��L"�p����	���&��pI!��h���S^G�Ϊ���y�:��.��/�D�#|��v�+��S`��~����NՒla�^����<����//�"�ґy0�s�VS$�\���_;��&�g^�W0s�ѻP�

�3���_J�ն�.bx�vo<�8�d��||��4�:9���#F+B,��V�����2�<�Pѿ:Q���vo0g��v�y<�э5L����S�˰�VJ<��65j�n�*C�j5��9��Lg~��16����>Z�:8!SI$5�H�r��>K�������6�
�m���R���vj��	����Ԩ����������]��'�S�5�^�L��o1�'˥vcL)����ud��X���tޱQ2h;���v�ׯ^�gO�R��O���w��Ҍ!�ф�ď�;�=��0N�*[��ZX;%��O����R2��2�0䧧vM�=�Y��[�ؼ���}�~��>��|}n�i۪�J���l6��20e$xd� p>ƷǤ�*�(����sf���Qy�vdab����8a�R̈́�W��K���Rqo�g����{�4�[vBPb&tL/=�?e���g����{�em�Jx�ɜ��L�);eޕ��۰?�s�q��U|(�!OR��.T>���@m��&�`���j�T�� z����$��0D0�mc�R�!*�P�myS�t� �ٛ�>�����Ym��{�+���CJq/
�-ֻi$�b�ɸ�s�0N���NT".�>���Te��E��X�.b���=��ކ{<9<(	Z�g��*	;�Dv�͡W�L}N�\��0P+�c����+3��Ӈ��D�6�3�����M�!D��
2��.�U�ڢd�G<X��/�|�y���l���q�J�NI��|n��7z���������l�ۨ��`��.�K�u�E9)�]b��Ҕr�k1E���B�E\��r���Tjŏh;vdsvn8)6O�_�|i�5>�|����&���Q�*T؀�s���D1Ñ�By��ݠ�@�%���&e�yS��JZ0V�	
���j�h���.�o��������2i�������(�e��
wl�{�9��=�����<l�U����J�JY�!.1J�o�'��֦��p��Q}F��/Q)U�M0|���G���C�&��N��u��;����W���c��K�?i����;���'O���O���p24��o�æ��n�va<M�i�j8��S�B%�0pKer��K�ǂt���l��ؒ��-�J
GSBF��۷o�W��X���Ƶ%�!��z�JzL���2-X���H�x0E+aeN����J�a�ȣ3���雦�z�B4Y7�	������w�x�}r̔�C����eڠ�26������_�+���[���t�a�Dx���1q�J��,V|Q��!xIQQ�"O���@1��s���7�p����`����n�Q��,�n��\%N�~S�m_,�w~�V%`���O&<�6p�e'n��Y�Z�,��g��K���a��2k��wP�C����0�N�1J�4�DŢz=O:xf�Xp+#E�x,�5�f��9�F%
��o~�[��0�/��(�~0�����fg��+9ԫt3����j���"��̽���5q�]k��������zE�A���H��u�d2����]�����Ci�qt��������ϟ�b��a\����h��.��B�.]gN���G��K�Qa�L�N�U�I4����"�MY�@l�*�����%/�����_q�^B瘡W�mChw#+�rW�+��k(f��F
���Q��k�k�[�We�2l��S����d�o�b�r:������zmu��B�M��[$\�)�wGά8����[��OG��F[�͖p�+�IȈ����m������;n���>��c�m&!j�?��lp���A�D���&��%h�I�U$glB�U4x/�M@z ����ij?���{Ǯ�Ϸ;�,����G]@����6B��jM����G%,n1[��yG�O�Jÿ�O���)�0bZ��)x���і��SP������*o� ��؟���F�ڄ�1fK{��j�E{K���s�&���CaT������e��I��<6��[�8�mӳRb������:�M��Y�(P:O^�ѧ��C�iK�2�g~�%�/��!�pKwR8n}��h+���*FN��}f��y��?81<���h+�*>H8bnS-JE.��W8l$����qlJ�;�ލ���HZ2!z�J���d�1{�8��l����3�~�F�=~�,��%�~��خ��A5o�+���;��ޟ��f]�~�+������M��� ��������`4�!��QEk��1{6��"=����X;ULLnmY��C5�E����x�q�T
�l�55����]��J-jX�%	�K���#��"�x	�*�0��p㛰@�xC����\y�kM{Svjc=qq�g�`�?u�%��p%�Xت�""�"��wPd�}��w�{=[y�v�ÁGA�T��"�w4D0�+������w��і�y��o*8��=u��f�{.XC�h��'g0O-ܺ��-sN(I�j-L��N!�#<��!�ҷ�s7�}�7��ȿ:�A�Ӿ�3`m��4P	����$�k�޺ ����u3z՘��B	R̘�ߘ��EC~�s$G��g}��|S]P�XK����" �*�c��~�2ե� S��BL:x8�p���l�Q=�b6:���J��_�F�� g1�1V��%��</hK������<<�c�l11<_nH�IS%m�#췶+��>��{`��c!Y�*��Rk�3:x���y�'po؏������~g�fC\p�f_�d��Mr���.S?�h�
*a^���7e>�RN�B���X-��HoA�b1S��� c���ᓧL,}ʴfq?S�5qH�L��.=3�?�=��)���0 �ss����4h'�$��tol~��|����5�lS�獹k��yW���lH،޺�����l�����6y�ư��_��QJQ1���5������wy���ۑ_��eզ���߳��VȢ�hGl�S��{���f��K��F8���-F�p-*q�.�I}��<={�<}������{��/�L_~��e�Qr�J�2��<�`�S��״e���Zi[�`"<�H��x���:�J|Ԡ��Ʉ��LkNb�޿��b�=U�#'z����P�0{FJHذ��P�Ht�ʛ���'+���C��-��D��:����H�\F��lP��69v*�[u��!����X�H�7�_�`a�N�3kt*uM��U%L
g.�Q�!�8�:*��68.I��B��}w��Dr�Z���]�L�M߹u۸�[��Ċ?�Uw�v�9��s�9gs���d�@=�MUu'Q�a�@�MPR)�el���W�I�6)��2ԟ���j�3Y��3ӽN��-����g�����8g5y����Ώ�Lo^�v���T���C<�UKL��L�ڥ���|T��#��7�̆�^���~�5Р �?8!��S�Y8�Ņ�Ǹ�*����N]�P�3d�ǘQꐚc!�Ÿu}TSŚ��x�%f�w]`zx�%t1غ�Y����$����T�f�A�gIe�S���b~�<�~�,�#��%���Z�%�.���a$,ԦAp�whڄ8��C��rƲK@9#U���_�Oφi��'f��VE쓑����l��(CJ��Z�����9J�'�����Hs��,�A/+����w�]��/�79�N$l�M`M<�2$:6�˄n��g9;��\���75=��E#Մ�p��}h���1m���/����e���<�ﹰ3WEgN�mM��*����
��}/����[ń3��L�g4�a�-CV������]z���׶�pHn`�M"m��-�Co�zXm.���zZ��RqQMNI�@U?��"���F]w����<��C^�x��熐�Ȟ?>;N!�溼�N�Z�F���:V�Wn��<�iZ&��yP�藶2��.aOS
�⒝M�:�+}�+�g*�K���q3 oTmRDi��w,m�dXl�U��d�oʖ�)m	���w-��+kõrYW��"Px��f�^k��^og�w%HLob`9�m0j@y��뺦h���Oo���G�4���@�6�yc���
;w`��A��~��)�L�p�{�r�C���bx��6���
����j�GrA�#�'�ُ��U�B��d��sR�,	�����ca�`�.�aZ���7������E?��	a�d���t�e�~�16�Ǥ�K���/���-Po��T��x�v��Tl&�x��<~��޻g���a�ċ�XT�>,,���q//"���l�6�mL+�܍.�b�5�k=߫2�bQ��qSs���dֿ��ͨ7/�LK��q3H̐!�S<wHn��&j�4?$�c�~6,&[�3�
,��Cc:ۘ؏L�zҋ���a��4V#�E[x.k����16VQ'�~��si�I���j%����^��)a��i�{�f?��mO�{��L#z�j�[;c��F\Z�H�|�t�P��}���GJ�-�������3�5����n�����)��#`���dȌ	��M��$�]aAa'�2�b-�)��b��F\Na��ә'��8�x�lJ*���׾�*^G�Ս���d��)�J�FVJ�ŴS����ՄJ��Uo�U�/��=|�0}��ז8�P������p��O$��͆�hV|���I���e�+Fdk���
�_W�;?ӕ����ޣ��3-�Bz�08 ���ݺp�⽉����5��`�|d�������y���cNV7����o��8�}/��F���6)�A��BXH�>�<f�;�"�G��E0��Nߦs��e�hs���茆��,7������K�׳�X��В�ڰ��Δ$��Mq�~ʫZ�
��yQӿ?3q�g��~2��ɽH���յ#~z�=��0�²F�v� �����a�{�u���z�����I���H(�a)v�1��q�U�"m��~�!a�Dӥ����'���P�U�֬���	�ɫd��%�jEj�	�I�aP�8,��Ϻ����1<���khi�W����{@��̴�-L�d`	�F~c�w������}Ć��m�A��&��w��ϖ����K�{kT�ɛ��Glc��rs�0j�l<70�'�4Z� {zv���UA<%��F)�n��s�}�6&V �G�_�(��	��>#"0hf���86]�Y�?��rp�X%�kz�S��mx���Z�9.�a0�`�vPՅu��0�J_�ݧ�'&��Ffd�����}+,Fə��EV���s�a��K� lKZ:T5��|�O��ĠT&gGIQ�q*ȄOR��	|���&��<Ŝcbc�X�������nG7��9�>���?|�����H�{��f#��nY`dPSr�=lÚ�O�d�]k��Z���֚��ܽL��'�kQ~G��*�y8�_|a���B�?�sN,�6�5���.'n����;rG��)-��ŋ��ts�U!/�����^� `s���>H�MԜ�[;��QqS�@�Z����I�}L��v�Ț(�?:,�ș��%�E<���8�H�޼��r|cq}�ǄQ5��X۱�6��	Ɓ\Ri,�g�3#;FTP&����3�8��ͥ�F�H�lܑ����"�  ��H��~���ڌі�aщ���_�6S8#��bI��܇θ�x<���̛����;4F��KQ�UH�Q��6��a���EK�ԹQ�|P��Im^*D����|�	��n�[�]��L��Pw���<Y=��o��I<+�6�y�0�B���~��O�R���5��Z@;V�H�B�A�Ob�k�u�wo�y�0��b4�S�Dq��O�����We��8�^&R�s�DE�~��v�������F�F�9p^oq}a�<�DU�h��ydJE�� ��<Je�����������Ed�܌�������7L|J�}�I�mYW߳�'V�i���o��席m�U�)���,�]�q�M�;5�fS��׊�l������ʒ�^�aF#���[�vq�2��S&5I����Шs�M$b}�����>l��0��Z�,�LF��T�C`�a���٣=<0��`{������
!c^j��:��������&i>�qc��.�p��k�1yAʾv����h�!�Đ�Blǫ ;�5�I�%k������Z��0ʃ�����4*e��3���c=��D��%�D���r�'�eq��_A�PI-��r��R�\I��w+�fB�����db���L�I��r��f�>K|����%�Mj��Ϣ�	W�Ϗ��
��6ucݸ�[�����{�s�u�)�h�6�e2���S�H�HUg���DbIjRf4���c�0��8���� Ff�֫-j*6�s� ��n����ίt-���ZK���������u���!��`��6�f�/���<�� u��㨆�l�X���r���Ζ�+1�vM�SMTL�D=T%�ںcSB�|i���	"�ף�(��}��S�,�j�]Pث��F[sAS"��*{ڷ��ݴK�%��A���P,��p�R�t��;��2Z�h�->�35�n����o"|vA�:�G|��l����۸���fDL\(V�h4��I%�?���x�F���M����4d�;� �m��S�d��c����"G��d+W(Ai�27Ei���)�"kja�K��$(E׳kTeXI����;%�C�G�r�<P׿E��;��f.�Rg&x��
e1V����j}�Ɋ��|���Q1͎��~���_�9��N6�4�";��%���}���cgo�aLi�B��TOHX����S�	 �IjW�%	v��\pD������<7unդ�k-�k�e��'�E[�s���w�u��<`�HV�/������&pO�;N{Nɶ����V�'��^��?cM�I�l7��#�>�1��Nwb��[~��]�*�9���P�j�v�~[�������rx&Q�h�� �G�N���M�f�䖚;��	!���JY2�"�.�Ehp/P��b�ok 	����j��\�!�h��'�Ql�k�DC��jC��ŕ'���f�cP�W��c��p�.o��G��4��S�D�O^w�0��:f2����2�b"�}�I���.���6��:E�nx��}�Ml�����%"d�,�ua���Zz?�]x�,Aab+i{��X%^'z%��Z�v�`���ޟ�Y�!�Si�7[2cM0��p�"�o�ݭ��ǎ:S�r��s<�ݑ��"A"�Q����H�Dэډ8��O�ef&-lߍ�)g��I��1�x��تr�5�^ƕ6����x9p}�S)R�_F���߹z�b�`��\�*��J.���b΄O�1&�2	x����U\ۮ�M9l
�ﳤkߐ��ʏcPü4�T���	�[�ͷm��R����˙Y��3�j�`I��6��H���R�	V�(k�R�OSP���%.X��~�W��$���<�.f@�3�ro��ӥ�z���)3�{�N��f�0ɮ�cul�0[�����Z���^���k�̍��G�Fڢ�Hwcl�J~�\"�l%�F�ro��$�'�ؕt 6jb߽{���hW�{}���\��<U7�l���q�JM�d��L6�(����I�Y�ɦ��=5.\��+�V�^�����#)_��0̓W�f�ڐ���<�}X�nvU_A2�ߎ=�A��/q'/���!:�gK\5<��ʚ]���������	Ob"�1݄�o�gZrfU�P���M)�s�����4��w�)c$�ρy֢d`�vs��k�@!�Fb��pp1���ޫ���46�5�F�H�G'�{����)�{��#�Ɣ���LT<����f6��*�T���i�G#�p}0�ɍM�m7���ףO6��懇��/�W�m������R�Ri�Ί��9���a��I�vԝԻ�N�m#�x|�Rs��ʾ����YE�FV b~u5�Rm�=5�K\?�M7Ơ��)B��rR��
��[9��-U6ܤ׼T0j�ɛu([�6�IY��YO��/*OrO��ş�Bγ�c�O?]WE�,Y����Y���g���ΎBQ�iT��%��l�Zcb�&��p��%3���3r�wKZ��-ZDm�KP�*�QG�Gq���ӊ�js��x?0����;��'�F�unB'!U/k���vY�F��N񙰼S.��!L�Sl�F���l��rT�9A7�
�-�t��A�q+zc����Ax�8L g�^1>z
W�·�3�|ΎM�j��/�}�<�ԼD��M����fԼ�=p{VulU�pdG�<���ءOԣG�͓� RT���SR��Q����%&V�W��7Q+V":��ZS4����w�g�%��Y�Y}�̨;vO�*��$	a !�"������5,�w�qAn*�-���<FҥMX�9I֭� �"V�5O��%L���)��Ż�2�D��B$I;ϩ5Ƃt��O��
]�L .�
ɯn�U$'\y��x�tFYb�9"��uY�7b�v>�TE�G�F��yOET$!�h�^P��:������4���Xsp�rhGU�QI�ﶵ�L�����7à��$��B��0)��R`xKz��Sp���ɓ'f�`T0y\l�r�,�ML�)�dKD�ת�N	&�YK�4B�i
��p);�NI�LE�e^��9f�:~;�Ϫx6�������X�W�/�x�Q����V[n��U��3������rv)��J�E�Y3���d���6�E������~S���|zQ�y�;�S�!�ƶ^K}�{�{�,IF�&����u.�{�k�><)垟�z�~��V^f�>�)�.��ldQ�4�h?�_���_�S=d{�i�Q��sa�lr�`�n�k�X�*�]�R5�W��o�1U��nL�7�nZ���>�.���9%�uO�|bޝ)P�����Fm��H��hb�/��S�#�,�uAmqJM|��+�&�+��4U��Z��j�ro�O����g@!j��U��*�q�y�6�z�*�0����C�r�b�Z�g���I�W���3�v��R$��(��+Z��
��!�]���3�yoAj��k�P�JYxN�D����B=�&{���$�Kɮ���7�f}Jx����{7F��0���^24�m���9gZr�u��CJQi�Z�8U�b~��%c|kF0~��d6��X�sp(���cjf܅TV��0�p&��]w�
�PǸ�y���4������7��"h{q;q}��h'�Z� �?UAw�g?�e��^��s�%�;<������~&�+�{�q�M�������|Wx���^��bx�f
!��Y�08®�8�����l�'fS3�����	�RR͙����t�J*.D|�Ĉq �����5y��AQm�U���ĠSu�8��|q�cx@UC��Pc*�:���E�Ŭ���"w5M%�kz�<��|?��t�y��0�����7�f�����~{ZOa��P�H ��DsQT�L���h�����E��w9^{tvj��Y��������9�Z0�n�J8j�S�U_�]U��iLn��z��
��`�Eqvސ�m�W��U8����w�,�F��s�p.�b��6���GȀg>��Ԡ.���%�,[�t�+z��T<^�,I(�\��RX9�TmT��7�H�7=��G�P]�'��mR~4��q����v̹�L�HFq�$\ʒr���^�j�ɫ��W'�{��*|2����c�s>��6<���ɼ��Q'nڭv������Pog/�;�:.6�^�����6�E���2ڭx����7�_d��X�M6�<�����po��^�ҳ$s���ĈBި�+��7I������-[�%\f��觋p7`2�I��;�i��1NΦ�S���;��ݻ��j��?eg�E�':�0�{���ꈡVʗWw���:�/�$�D��#[�[���+�:��d�SYI�$�^�:hpb0ޗ�KpZ�-�&��m��Q�_|�=��/{Je�E��a����I��qcB��h�I;a�I�)�r�y�QUwl�J�B�y"�J�YA"$hQ��:�k�V[����Jδ�>�ݫ``V����c�B��D�q>֫�|>�n��uC��X�A��h��0Rx��P��>��;=�����7����sz��T^g���FŐ�,�-���>Ή!{�\�kܑ��]�A8�yŽ6�:O*��7ޚ��w�����a�� �FC��`�M��ʤ5�p���ߔ�:K���G~�e*��v��OE.��v,�M�W�aSI��k�`�\ֲJ��������ϊ=<:��>Q�*�B(������q3jb�Xj|R�����~,6�L� j�'�ư-�CY��LБ��2�l��5�5�)��O�]��'ɪ���?��\He�@JQ��o�,jw�-�����PKS�g�����}h6�n0���5�r<�J��vM
s镻�L5�rSj��������$d��2����\{BE)U����)�S%l`���׍�=B�h��驧��8��\���M/�����
N(SB1��:O@�x9Rɣ����vB`�)UQ��GO�~�����ѓ�셅<*�"W��!�����ۄ����n����hPe�����T�9-��$��Yh�I���_���ƵA�
�w�d0k���
[�bf얆Am	0��X�d�;z$��Ґz�0������wCyq���]`�B/���N�E���!Yq��40��y\���K�w�^�}�v�ꫯ"+�dS��T�`[�ɚoV[��2q��#���*��K���+GH�U���ͬo@U޲Ċ�]V��gR(q�r�,��w� �l9E�ט]�$�/7!0I:��5�Kżҗ/_Q��|!�g��Rz�}OvO�)Z�ob���g�R�������O(�sa�%�U�(_3��V/՝��m?*\��u��ٟ��Ų|<W�zc�aPn�@����i5ySR�jCĠ�L���Ճ�(J
�_�Ʈ��E!�H�6Iw��D�4[{����;I��D�̙-̵��q 78�	o�[OoM�c�'�i��H�����m�e��q�������8u�4+|BO)q)] �lǊ0kA<5UU̜�PØ���N0J���8zQK�p�����������8�2�\�J�HsD�x*u>��xa������~�"�4�9QЄ���}b������<���ׯ�����|``�V�<ЋoA}Я�s�Q��WlC��G~���#�ټ|��	 �G��ΰC?�=�V/���RƱ6��	��L�ub�U��~̸S�Q�)+w��o�8�3?n�Am��r#@�$������~� ��nnI�T��R���r�EYL�S�5��kz[�񬚄��G�s��q�|'���<�ub��/�=x���w[Fxjq5�������읜6�i�x޲���hV�&��V��*��r��"��m�W�U���
���m��Z�sq�e�ɬp�"�]G��lbyd��0�/��Z᯷�� �nB�[g�L�Y���Eo�Du��b>v���nb2�5&�#<5�N�?���g��s �-^�B}%�px���<b�l1��xC���}i�jT���W���j�#��1M�o����^>!>�F
�-m��M7�7Ƞr3�V�!�Dɂb!��aOE��\S
�P�ca���S��j�N�K�x�]#k�E�H$廇:S$���o�CE�N�~����$�U�(���z89	�!��q��4���+]ڽC�q6�[{�a�IMwd.lB����DR���'����D�]Y�w��3-�U-�m=G��楕 m>��	GkсpÚ�����&�=8�
�£�.��"\?�`0�� ��tR�~��Vx��
��q7��6�j�v�	��4�{:��(C}���o��b�Te��_�b�}7�F�{��������A���j�R�7��"�\D�K�qmJ �)ǘ$y�Y^OM�?�O���{� �Z�{�2�="a�k־��RC�-ED*�^I @��"�;��%x��"4��I�a�Q��t��4�\_�y��6�.�P��l����:�j0��5�õo'_4=S��E"�ײ�)1,ł���bl���a��R�ZO��*�RZJ�U��j����z_{�ٟ9d�jS9]�gm�/��~V}�FUa�̂�X��^%����h:��w�@�)��J~��w��4ajl�Ö��CR�~�Y����0�H"���{�"�)�w+]pBO-[��rj���/����\���䰎�:L$,]Ձm��
�w�k-7j�DqH��8��(�O>�?��~�Ǎ2�80	q�~\���x&�<׉�f���s��@l^g��y��Ք���e�)6W�4g#���'��O���2�-)�BJ*�!=7�����R�solV���P+�80���̸�vQ�o���7�� ;
p[ჩ�'&��<��ǆ��*�d$�`���ˆ]*�q�?�hi�}^Y�m/'Oԥ˺@ͫ������C�cf�!��{;�SƩJ�YT�
�R-UV�c)W�)B�\|�V�� ������"c���d�t\����^Q�ˍ�������N��L |��̉yx�JG�Am�G���+���;c/���d�Gl�P5��<Ø��g�7��Q����
�����ɍ�<��ۓZ5�-k���S�#���Z{�gۍK���`[y���̝�����Oz���Ԋ$Ƿ )'_`�āY_U�H��ϑu�&V2�U��W�^�&�70,���J�첉{b^:��ݰ�$�,/k�6�T�R�lO�����q���T38?N�'.8���Ԃ/r^�*]��`��6�BC�+<�k����z�Zo��1_��M��t��/
��Zvo��9W.������U�GPFDPr+s^�TOI^�n��#�`���X4��ꌋ����
W�f����������v�Ҟhܩ�n���b�Dz"�{��hj>����Ơ�$�k�;�����E�P��2�6�����4-�bM�NڥZ���)wH��HUkm��G���!�싁��?e�jng���^�6���8�g�g�}��r��0�Xd/^����B�l�7�9��s�}�����J7�����'�V$/<B�qe2v'FV��ȧ��<�����o�y�ni��?e�U� ҄�#biH��=te���ý��7N��3�>��c:���E1[���j��	��V.���yY�ʀ-�����x@�����y_���޽���7�C���G����9׆�T�[�dZ�$�����@���~b![9�"�+!�뷪�Ġ�6դ���Ę��p�NXxL�s0&%����>{o=�1��jo�������&�g(�c��J��l��� ޳�*�,�C&8J�h�ڍ]�*J�+o�b������������������*] ʘ��a6�yEA��qBx��ਧ;��сe�ONnY�6��0�K���	>��$XmSX.�{�̮�j¹U�Vм����:��5�E�J3���M{�N���l:6�N�iCԐ�lڵ�����%E������}Ud���Ko9��*�x;��;|���m�.�ZG
�v˚�)�Q�R�o��쪫�	���%���yH~���Qlw��V��v�^�6o��Ƞ5��R�sS҄���u��eA},~_u�x�ԁ�&WuS���A.����߇�u�ׂ��ίt|2��������@h�k�%��pG*�S�_���z4"�'!d�7�t��N���+[�3�;�����V�|�>v�}���kv�84,3ۤ<e�{�.#��zY.]O�������ac�g�!��u�ȕ���#���EB=�\R�����9|��m f�֨�>���������?�;�路o������[\kj[b��u��݆2��lx�p}�$�jӌ�Q��\q��I����G��4�!1�VK�r�{"��s��m�i�t��ـ�̞����u��ᣵ����vaK�~�Ѕ""����4�yd[޳�O��MK�i��'Y�<�=U����� Vu)$Eמ$J^m�1���v[��&X� ����Yb�aB�\��,$,M��6�m��w����6�(�x��v޲pV��Ȅ�i��m�\\���:�)���'އp-��1�Lh
}N�'5��/�z,�T���z�\�q��*�{���nU�M�c�v�x���A��]��8(K�v����M:mW�I�X�Ǌ�����$0�8L���P_f��Pkp䪜d���FU}�U�AG	�t�����6�tyv>���Hvdr��m�(��;��'_}�~����"{��-=�MԢ��ʰb�LP��ۗw1�U��l���^~����ٴq��ߋ�T�>�9��V�!��߷6����q��0��b���s��j�Բ՜����?��.��dU��]�䞎��&�j$\���Y�!�%�:�G�חe����*1E �d�Ol��d�	�Jf�N�yc�mjW��[۝C���ڿV�ō˜���U&�����JPO�G�o�ש���q�)�t1*\A�gfHu�Bj�F��}�'��L�,<׼�  x⻐����܋�Rnt�#C�	{vzf�Tޏyl�c+tX�Bd�&�R�d��ie�L4x��@�1&�*N,�J}Ҟ#5%�/'����n�T�K>M�^�J?��4�|��<Kx ��R������K����O���o,y�>TE^^Cm�qښg�t\��S#�Vz�*�<[DC����p�ɥ��!y-$�aPž�/�b��h4�c}P5i��m���F���"N��a���S�G>����-����Q7��2�*ڂ
x�yxC`��V�yj��>.I����ItR��zks`Ù�l=g�O(������{��Sp�������E��j��c��@�`��ڧ&�b���^R�����#�#��3�^']�gO�hp��$=�O.�=H�@H���㣋��]L{�����Ù�R��0�_���m�⦡�3{��/���fǚ\L���p�t�N�;�I!i�z{h�q�����a�mw�X�����w���w�������_��g�LFŴ?��LT�A	qc�Һ0lV�,$���Ђ:8���V�G�����6i�
L�0�g�b,^� �����QH����đ�/~�n�D+��W$�CD��d78M���|�Mu3�w)FDx��\�pA�JP�^��If���<��Uk¼dz��4G�5�\^����1l4�Ϣ��{^�z�D{�!�X��w.p=�ܜ��S���^��(�nj�qe~������M=~��8-]���P�)7�6O����������`5ޅ�^42�P�G�&�('�x�����nha���Yzj����̸�yK�W�"~Xވם��a(!�grl&�\��".L�n��L��z�g�0���wz��괰�3|��Q�߽uX �,����'>�C	�b��X�?4i�)U�!]O�emjF��d�W_��5+1}�Q2*1�]pQs�p��\"1��Bs��Е�z�z�,���n$�Wa���U�Β�ǚB�(M)�ISs�fPX0���NJ�M��Jx�/�-""�#i��-��:�\�R�SJ1��jGov���d�T��$t�/�:�cŽuQ�!�z�Fb��C�L�%6c�r�u5s"lD��}��ޠ�o4{!�<��˾�c�(���İ�XgZ�j�LL�a���`�Ō�;��9$���{�浽��l}kb��A�|"z�"ɣwk߶7��]c�o=��9�w������`ċl5GE�g`���M,<���򦀎��B��������������O�
���p97&U�>IJ����Y��[7����AIoN5���Ej�Z�k�"���"�V<�?��.g�0���K�Q`�)D�E_ʁ
Ґ�8
 �-�و��0sr#�4�J�ʣ��2�*a��Y��QE@V
J
�56tE�
-vP�1�Z��$����U��T7R�ĕ�j;KDn���0�a�����Q�ǰ]�Nt�OؼL�pI���]��-*T�.���-<ӛ���!�1M͍M^ͳ\2�5ljJ�v� �}ZaG��=������/_�1}6��w��0�n�~l���YW� |�}� ɂv8� L74�x���{lpWy��-*�#*&��F}VC�fN4��B�`�l0��JR�I�:�,nMa�U:�� �����>;;M��������OfP�{у�SqN~Z�	�Ө�_�k� �r@^�w?84�KJ���<���e�D2���F&�PW
<�2�B@��y�.���69?�v���$&>6!��qr��k���u3��,4SQwv�b/i���g�2������!�#����f�Sy�%I�jr�=uURt�M������U����z��;�pf��~���sAT��=:�τ�p@�G*�X���@����LM[���}��u�R�8�{��>�kR��\J
T5�v���h1��h�.l �wgI�?���ԫׯͻ�c!H̆x����VO'��w���ᙺ �g�k���h����֌�!'`%@wޞ����P�
�l��% r!����W�d��pC��E��w��� c�"�`���H�{��rE��'Ӽ���Ȩ2Mr��_q�Zi~ޡj�:�|uE>4�"���`�i޽wwތ^]L�!oJ���e�#�Y|�G�1�F�(�T���W�ԝu��ʼۊ��-�h��V�+~�q�κ�}�ٍ;��GAp�wlj��e�L� *��~O6��0_���&윛�#zhs�7��Ƙ���n%SGx^j�~��5XR�h���T'dZ#m�EO���7�BJ�~w�
�꺀��>�����
�-�B7��x/zWFJ��&ХI��
R�_��"�9'J����"�п��{˸������G��-�-�d�s㨢��4??��]wYdK~0#;M0�n�9��8���t/M�����Х*�l�4_�A�<RE	x����8w@)0�,��&ũ���I��}\�B3@j`�>�YUbS�A�y��(�*�a���̘z"o���4�f��$̢OXI�Z\��M��koP	�'+S�؍{�]٠v�(Ł��k�(���x��ݍ���k����<�B<��ܨJU�E��BA��KyB��q)|�e���K��T��B#�	���*!�揩�����W��U�����ͦ��Jl�/�7�s�%6������װ��5��uaaTG� N�g]�՘��Q����x���-@ ���� [�VM����V�������� o��}V�D�T��RPCE��J/ɹ��=�:�G�m�(�޹e�n5�ӎ�B��r��TE�'����&wG\e����Ŋ3�'��*����S�0��Wa����J���0 ����Ҽ��Z���q$������i��0p�&~��膠LD";����^  �T^�����c5�;9,�S���	cЧ��<�`/H*҄s4�F�_E�Hkz��<��6���ZkR1�ڄj����{�.h`� �������<�g��t�(R�j(o�q�c�y��Ġ��E"�,oV�������S��
[�)���JT�& &���{[\�m�Dx<�?�ǭiZ�t��cM9�Y{�J�w���31��Uv͂sNV���,��n-Q\K��HBGwS�v�H��9�:wR����΄5p�(`�|�����tMX ꫪ���:��U�at��8���4U3�P=��&�\����N..4U����c#�Ta�v^�
���U��hao$hJ���zA�B����X��i��a J	̓hs�<чDy�?��]ޅn�`��#A*8�E0ƫu�@ڲ,zK�nr%*��a�(�{��+����#�qqn���@J�M+m�6L�3'eƷ�0��{U�Ǫ���*�Q�%���6�
��__eoʁ���{R(�O�4X����`��S���{b"~��ߤ?�H�~��-�ќn6��ݷ	�C�Y�m�=z
2:����a�ob�
��E��%�+�!9�^B.,9����7��-w��kqm�^�
�Q0���0�)�ζWޣ=�{�ZbjGa���
��	h�	`�x�<A_D5�;h�����ϟ���kO5g�sohA��l�ý*�u��$�+x��Rq�:PU:w
�g�{c�H0����8�S�)T`�t�dŹXj�V,�7�ғ0ql:��C2������|�o-�K���8r��8IגZ�����o��h�6�aeЕ%Ji|�{�^�sP�����<�O���&]����h�fP�#9��Ul`�F"ܳ�o����㓉�h�RG��Z.���S��䕟Xa6a���SY_����.�<2������O��ܻ?=z�(=��K��ަ�O�7�s��]�֧���MS�RB�9Z%�DL��$8y
��`��6��S*/��e]�������2�OYk�Ja�mC�=lt�l50�imF����"���@q����l��C׃��
��6$,$����F�꺡����m՜�R`����o�ۻ�q��O�Q���|g��/�������o�3�N{�Gg��y�6L� 3U�T�I�HH@��3��ZK�ܴ��y���N	�u[y�Pn,xň�i�O�r�AŸY�r'9�Lu���z��դgޚ|�]��;�� �Ź9`@�oz_3~Sx���`H��j*7��YhU���Z��2RJ�qP�G4�?7��(�{�_����4��ӎ%a���k�T^�Ҭ�$�\���[]���3��<1i`���k�L�x�grc����u�I��(U�5�<0�id=�c�;O3���a}^N�IYڑF����Đ���j1c�>����ݹs;}��7V�䘠ӆ�0>�}U���v��P�C4���ra�/X��zw�	su�;oYR�ز�j�f!��u��`{�^LhlQzZ�<i[n����S^��j�։�L�B<Vc>{T8�����h��Թ����0��9+����,��c��i���e���R�=�(�L&Rӆ!GV\z����rVG�DS�bbO|�!	ѱV���í%ܐ�B��\8�!5z��;���X�L�9��*�fj���9�h���r��\��,)�p�%8N0Rn�˹{��U�r����_�A��J���r��
S9��y��v�}�:�x '�7�_�`��9�C�[&���@Qj�-[
]�T%�v}����4�Q��(k��\m���*G�l�m�IE¹ÐY�|�C�νN�c��V���a\Lggo�0�B�<!��<DE��D�����O���u���$$ �d��+M5Y��Ջ�'���r��{D��5쮬���p b�M�L:�� ��|;oB{��֣{|v��Y��Ng���ꍫ�Şj"�綢�.��./����#�DU�UL_{%�bٍqO��tow���:����b>�1e���b��}����+�t��}$����i���U�R���ׇ��L�o?��X>����6O��YӲ8y�x���w.�b{	N��a
B��O��	%����5����P/&/�:����$
�4����2:��%?A�5��{%7�?P���6[Ye��]�<cGS<����/~��� �u�XQs ���<��Q���� �	j�J���;�u��^G4�n�WQ�ޖt6��7Z�&��x�'%˕_��4��T�hYn
5�w���=zDZ
�31��4��������DZ�J	���M�*�)o8�i+;�#��sM^�ހ�Q\�^�	��R�21��D*�yҩ�V��IL/0��W)/7g�<=p�[H�ݚ���Z�}�)�CyL��v�?�gD�f��lg���9����Ժ�hL�����KE؏C���%bk��_�Uz��M������y��9������=KK_br(�3
��a1��^[)T"N���(��B�y�z��Ax��B���6����{5x�Ą����%��y��!�ٗ��'�WyA�U7JT�.�ӷo�ح�wݝ��Ի�A_�~�����$TӀ{���FUE�Ks�j�q��$��,t�a��7�G�2��F�6��ԥ�ئpI.2�s��HҸ;�"��,Ř��I��x���:�PKx����qbL�����&&�-����x^P�,jP?o0�-�q~^J��.����B<}W��6Mk���hH�Qɭ���5�!?<ҵ)M)����ս�Zm�1�����sZX�&�Q��0�!�����!�<�z�l'ˆ{r"yhNEvTI��w����o�����8zN(LT�(B�(8T���7��"&�š/RKt�N�|�T��ABO,}�J��FT��ƁV�b�[ے�U��b���yy�;[�R~�Ƃ2ʍ��&��ц��#�쭫�7���-��"e
M�$`Tjچ�a8�\��c��K�f���uS�A�A?��t�*M�Ŀ�{6_}��e�_�|e�dؐr�R����v���;�ǫ8?*�Zc��;��،0^<��	�xIH
ѓ�鄰H�A�B�(���<���y���&&=�a��aˣu|����?^e�k��YVF�yw��mD�ztˋQ`DYߏ��g:���b��m<����͛�0�z3*���2+̌`��;��&B�7]�?�۟<^�� Y�^��SV���~�B7k/ݹ��Ixqp�ݽ�~C��R��8~0H0T��Ȕ'#O$�4��I,pI��Ay�v�(���f�|��${�����0끥�loa��I�]��S	ݎ�P��eN�̭�QGfХZ��Lەq]�����G.���
X|������2�$$���G�����{�L��yX)�P?�0��?�ɩ
o�#���t|�B0i��m.���r��K����N�=I��zw�E�Bi��M�ɧТΚ�(% ��Ja^(��<�=G&0�w�9��CpO�F�"�*��B�a����E����E�6���b�j���cP�E+��v���i���!Й6����f����?��?X菶O�=��P`���g;f�#cE���+�����r�����5�|��D���L��<��(O��CJ-(�<X[��^n�G�����s����T( �e�7\�Olb#1��e�F
�1�/��#S3����_���4b�5�[�W�[���s��K�7�E��1.v��{u�D𘞟׽�0 G?;��hX���{~�s�_�✒ޮ,:�0 �pː��=]��0Fh?��jx������g��Ma��ig�;c�
��rCq��h��`^㊨��X����Ն��=����߽w�q�c�d��#�h��	�DTq��O���Ï���p�&Q�7Ƞ6�����7U'%s��Y���B�-I�T�A���B*	<��s(h*N��Eě�篫���\�	W`Kf��Ӷ�̆�i����9����yb!�w4�����'�[�{V,��*.T��HR"�ڽE3�ޤ�	�ͱx���y!�Px[[	�}�H�߻o��j���dH�Y�%�d�	w���k���^�]M��C@�CG�=3>�`� �6��m�x�������#]�;\��l�2e�`�,��6�bc�!�*J����kCD�g��Սd�|�9ᐧ�5W#s�R�}��G*����-з���&h���g�����D%lF0�Pg{�����1���N���~��}�qﵹ�Pׁ���F��h�P[���cP�(��0���O�WOEy�>�wL:L*,�[����o~k����oӟ��'�B֕t�Pm��6��R�J�KI��'u�D��sZ�-Џ���+�OQi5�ނ���P9�����z���{���_K�?)�0L4�4Q~@�+,��ņ�3��UfhF�8+�<�� B}��{���
DnT��$a�%�Jٚ1-���"������{5l6B��ɻ�.��8V�������1�ϛޫ/�2ʸ���U�J�MBq�;�����x1�K���Q8�ko4q��ub3�����D	i0A�E)/���Ό,6`�0����c�=A F�b+ ������̾(r������庪���0����6v%"�)���w��7�A��y�Ch�68�й�j���׳��!ɻ7o����~={�V�\��۷F�ί�?��"�>a�yڥSORY�(�
-�Ja�l�1Zs�{P�І��t)�%�f�l
)Qe�,�D(n�9]�лA���}�����бVSg�=9$K?yl�
��#)L���qa���(���b�_5������&��P�����o�И�RVc;~f�&~,���Ȩ5��y<���6��o�?�`����D�(�K�Ԉ%��#m���ͤ=Ǟ�t+�Ɇkp:�U��$��Q�tx8�I�L�Y8�d7F��a��n]H�\S��;������޳���Q�7υ���9B;8r�C�&����d88��qG����;���cP���M�M<U�Nޒ�0�/p�	�?��<-��������e�����n�S�f���e����Ј�V],6k%#ˊ�cb�0�H~]Z����j)������>���ԟ���[;Ef����]|e�][GOD��
;�Uv&I,[Ki��s����	0>����z��}�}*-U%�F`�'��Jm	S��z"�C��5ɬ+��%��wGl��2�����d7ěA�0�
9ȶ��S�x-����{��/���hRo��l
j��H<��xNO����&���KIʞ~��z�(���\�x�o�^�J
��}bn#Q��	e�p0���b���.��B�ɸZw�����+ɫ�0�����d�&��E�.�J�x�DIW֓�*װ�]r��7B����gT��:�?��-�׃Uz��A�> ���s��Wc:�t}Qd�o͞��0}԰�����jŅ�W������0��33p8�KXD#�i�X{� �*)��ێ
GH.@��ڭS	��=9�w ;��������[x����;�g�
͞	�*��j��JDu�?=�֫Z.�=��6ݵ#�	͸]Ysܨ�Ԫ'o��B>ٻ�=�Бq�j��#�k-)$����G�)�S����6�Q�7p������5I�	_Bo�c�65@�|D$+���Ӭ�{ؘ���{��m�v�;�w��+�l��� ��T�3]������Z��c{o��aH�x�ȼT�tQAj�p�;r�c J{�͘˖j�K���X��8����^�R����y�G+'�8�1�������}0Hv�rb���{������r$�/�ͪ�i�5UB)�P�_F�"%e�z����H�٘�C�
�9A��ݛt�ޝ�?����o��o�o�q\m6�6)� ��OG�|�훅���5�yo��;�6Æ�Of���	l4Q���T�Q�jҡU	� 4�3U��3��x�s.�DY6pS�:��� ��jVwe��.���(��n�����	�4"���s*CcڧS�����Ќ_���Ͱ�v����"�+n��?]MV�siy�$]S~k����� ģ��Z��O�����6Z����o����GG�4��"?T�U����0���M�p6�V������ĹےӜk�'���
��7ժ��+��9�D#��g���F��H�B���mJm���=�gt2���X=fщ�s��.s\��O�c�0ui߲i����֨�X��t��\C�����2McM�}��/x�"j����C��򸊞Ex�<R�Y8/Jr�6�1���,(.b�?d�Ł�bgK�������lg�}��'�(R�ԒOx�̀K�3�}��g�^C���g�k�����J��ޗԃ�e���Z���t�s.&c���	�⼛1������R8���gr�H,8���^WG%
����4&]��@1vp���?��fr(O�*�ئ��dq�h�������vO�o��(Q���i�����2ݭܢ��q��-�Et�%o�6�N�Mj���M�!B�_BBf�c��z�ZO����@�=���{�J��{	!n��Q�6� +�IHl(�˙¿B}�;jD�aj�]�O�Kc�Z#��Eڏ���ROe����6埀~���`��G`v��ZC��Ғ�ƅ��5����{���%�U02��?H_�����������_�5����_UF��j�k_�Lp�ը�j��Z� ����<#�W�joi2E�+)�����#tEk�٘
#�`\Sb��l�j�Z��ވQc=�$���>:\�[z%K39��	ߊp�����]q���c�_����kO�br?�Ǚ^�f&ּ�rC�����A P�u�������Eb�d)V���gڷl��U��@����%�i-ڶ�	�e�[8��)���_3���Wڕ$E�7f�<'
�絨�뢴�$Hz!�7����:����"��J]��ds5��ދ�Q��r@R��?u,x��>�X~F����h�hV��a��z�lf�U�X�(j�b1 �����H�߿����[}�^�����Gs8��P���b!Hl�(7[�����0ޓ�)A%(Z��b`I�I	�m�OZ�0RV�;�ί��k�s˳�_͛�Ĭ�DOL0X�'LR�һ4F݀..�]�J"�K��3սC�:r]R�>_��
c�q��T�A�;�O�4��e`�|���֖��K3�B��7��0ze���{�ڷ�y�P�}���~g�:���cM�p���fyiђ5�$S�
P�.k���X#*�f�
;/%>�N�ITCye]�C�Z;���ڹa��bc�n�[Um���M<n�Am=#���تވ��Z��X5O�]��a����*��7���	�>ThEc
#�	c�P����e,�9�R�O��o�$ͮ�9u�!��^ع�ih<�D꾰,>��g�:����$fO�����wFچ�P]�ѻ�ݠz�еi�L�*hj(1�������ܛ0o�~��`�Ô	�����r�TL �!s�B�yS�#x���C�y�����ӷ�|�I+_$��&}�w^��MN�a-�"��v�]0
�7�%���<��JAckr`�u�ƍ�H�x�r��~���5 �r��:�R�f�^P�x<:5�pY�3�b�M�Z�zŘ��������4��y���"y\���,$%e:
;�uǸF���~G���H����/�w�}�����K���7W�G� �5V$Kwo����ڕ���)|�Ih�j���*%�r�㛦�f�$Y�=0R����<��!�������IƣG_X������^S�7kH/���}K`�h �&����/mM���x�M��@Q�^^��x/���Ƅ�O��=�k�P	<|`����¨yҙ}'<�#J?b�R�ͻ�F�ÆLr׳��Qɨ��z��� F�'o�۫x��H!\���^�djǤ0��[�w�G
Cz�$���3U߄N�!��d8�ttγ���Vc��Ka����o���r�,�Z~��+��"��NO�V�Ԟ7��nX!>�CO��9�W�!ҟ���e�/X�hd��k��y�cҾ�ohH'����;U�o�ͅ�Ʉ)B!#KO��!5������޵K�#C�+N�=fh�C�L��1��e\)��]��:��5��r|������/F�n0u��]��G�@Uf�=�M��JN� q��L"��1	H4{|�N�f�?a߀[Vf�����6��R���j#;�"��݂��nj�+�����6�6��>�Wz˽ҁ���h3�f�ڀ��@r]��'��M�1MW�����<S�h����R�˶eK,��I��|%12�0U����9i^ = ���W�B(x�0Z����!P^�:��3�m�Д�\F!u�V	�����������*����dr)�۠a���]И���KW��\���I�v!ͽT�V�|�p�z�5�k� ~mƯ�*h�-�N����ռ�� �@WZ:���%�`Po����Z���x��ٰB������%[�����ʼAC�$-�d�e$�*_���MY���M���q�;�cd��-nQ����J�����ʓP�6a��=�7
%!���ަ�0����%cz�m�1��Y~�%�7/���2����d��0���8�&��
�*BD/,�3*��0��~5� �|�浵PA���.=}�Բ�;���>s���_o^���@�W=�̫�mnP2h79YI�U�t|h���*�wb��;s��PIBƙ�.5r3�j�{���w":�~�)�C)��g_W�mޢ��k&��R�cA�+&Jl�jAmUh[������I?���h~������+�T�	0,P����O����|�Ҍ�AJ�7�T�ӷ*��B�TF,Η�_֭�� ǶW1_�}V��h��œ��ֽ;�X�z�
-�g+m��uTS=%h����{ē��5ƴ�q��xjT���6�7Ƞ�kC�@:B�O�E�>�8(�lm���-���c�SX�h�p�N3���p�������`������i5H�\����
��)~b���;��(K�Փf#���ڥ�(�w����a!y��A���}�20��j.}zI�-˅�D�u���c��:�iP�0��T����!���8�� 3���V�'�8�``�%�O�������Y'譾����_\�~hM3��;����j.��{�g��ϱ�^�l��O�ܟ��.�F����(tk�F݅�ԩ.���	B�0�V#�)���isC�ƴV��V1��������Y�sZ��;�>�ZR��G�����(,�Pҧ~(2�^��,,��B������	���P`k����}9Vx1���y}�sM�FH��sϊ�Yc�8�p����͟S�;��T&Z��pXGL�\"$�,>k���_x�<D8�ƵR���n��es+w���"X9u�U(g��F��*����0�y�n�0t���W���w���'��7`VP�����A��7�ҳ�k}��Mzw�nQŤ(�V߱c���a�G2I8�ɉ37�8:�B��rܦ��r����վp�S�tߔ`j����t�j��c�C]x��]�u/)�W �����o��E����4�n�u�N2;�n�Bd?]�ɱL|��@%<��t|�R>~��� ���/���T[�'][��6��K;�(G7!��e(D�&y��0אmɷ���55,� �����sf��ɞ��̦v�Iy�'V��#<������k��:����BX�td��	?�F�FH��@�6P|������j҈�:1���a��䭍=恵�g�p�2�Α]���z��15l�z��)d$@����>�Wy�"�c�Q�pӈ�TE�"�������Ԏ�{� ��}���|��Ij���~+M|Ѐ�Y�E�`f�Ҋ��37��$"�'{��~r"Յ5�Dp�Vޑ���Ld��l(]�ךH���h4�ب�V;����ŝ;.\m�k;[��T�Ǩ��z!�'�j7J����������{&V�h�i|#{Oc9�/�S"����71�-�^rd._�����&>ޜ�;�5G��[\���]ӊE�%4I����1�|l,��}3F��_��lW�dj��<�ج�k�l�sr��w.�F� 1C���ѳ`@�"�S��QIϒW�-0�H8�3�׃�Z�
��S�s�x�I���[kw䚡�׍{d���uO��KY>Ӹ��ק����^W����d�(u�X|m&�[z���ͪ��r���[{\����rj�?�,��d1s}ng%�u�F���:��<��n$/^��h�Zbi��g/uϱ`2��/ɚs���x��ku���e����b�,-�-芘�~R�w1�"����]��W�����80�k�^�x]ȿ,����~�;��׿ɟ�5^�h����J��F�KMի��`�0�d���ܲآ�9!	�.#��0{�ݡy�uS�zQ��j��'L+���u|��������b�:Z,��fA}�Q+!������RA���WQ˃~H�A}\��??ZU�Y�J֚�*�s]���ObP+J���TOf��3���:��Liʑ�����[��k����M8��.�t�J���/<�qa���)<]��&GNi�K�ԉxJ��c�ghiOբ޼ky&�S����\]bl�,�V�Ҁ6#��}>����3$���:���L����-$��8���+�{�w׌g�E��z�u<<Y	5�����qW�NN��O�ʧx,�Ѿ����{�O�W��1�4K/���ㄟ��R�x~����>�[j<�^�^���9W	7���	����bQE��;͖�9�AW��+���'*�TM[C�+��D��j�R)1�fU��Tᕖx��A���^�A��{���٤�%����a��4J�`F��W��f�K�W��y�{b�횊�Y�'�S[Ds�5�J6��0�%6�=_��������'�Pm`��z �RǾW�>��Psd@��sb��)�$�-���RY}G�Vj�<�K��a���ޛ�7�3Y� )ٹT�=������t��k�tZ"qˉ��,*%�2KQ�Lq��XP�{�4 ��:������U]X>��;���(�K��^	��Qt`��ud�q@�߼��j��zl���ԟ\������)4�
��Qk:����e�-�-�]R����Smwܩ�&~ߞ#�.�Nj�r��uЄJAvJ���	a��_Y��{�8��z�8#�}q<��p,�!�~��,GY_���u���+�d���&����t|�\���:vrU�r*h�h[!EM%����E���O�Kd�͚Q��O/P��t!������}�I�9(�SK��]g�1����}�`u�1J�!vΨ�6�t� ��Ȥ�s��
����H�CV���Mg@3ߤF�>_�-��R��1�J���4(߰%���أ����}���U�P�p�d ��ԙɠ���2c���N��;��l"���J�$����@ 5�A]����{�紏���2@�.F�Gr�f�Uj���A�u�+��'ZB�qأ�;RJ���7;��c����̼֨�9y��X��RM����1q��pҥ����M5�66\���P�M�c��1���P_� ��>̑�|K��i�Ώ�9��65>�y��M\G9U�<~m2�[��g�R�ժ�Z��}����hTz�UU�p��ONW�F�Ix�N��S�c$jBvM0��m�AU�!�������18�lr�D��f���i�^:lL|��N;FtVOY��n�҂X�tK_�/KS�J��Rƅ'�4gt��Ih@=3c��ҹ;��r�0qD�Jn{
��(�&���r%n�oo`�`УOri��lg5k��[���Z�pPOA��%�ɭ���_a���� U&IY�d�Ԁze��*���И!�[#���޾�$٪�)3 ��؈�z���m�ASO���PK�NI"��C��N�A�pܴ4�~�cZ�EV����ڱ��j�A����T�crNH�E�WTA���R���`C���ou`&]J�:$v5Y8�0�d���:����Y�Ԭ�^;������ ��
�f�����xW��NT��}ä�԰��2�c�<���P�.4:���^���iXjJ�d-	xX��Q[��C�Z M^��Y�+1�媶�4�#��]*XG������e�r��!LX0��b�t���y��@�GJ@�@����ݠ��y�2i?$P��YU'��`M e�5����LvfU���z�H��͞4�N3q��X��v�����q���֜�~��Q�`�; kig�$ޣp��Z������O�4��$e�	���C��6^��̯���X��o���8+���LTt�P�s�6f6+����78T�C%���[��2Z��`��ȧ�ٖ^m4�ڈ5�+�6�V{s:���yx6)P1yV*DJ6�io��g5~9I�����Z�]��HF;.��!��c�۽�P6�d��Z�R ��e�Y@&��h(�Z�A� ��r%@mfqt;�T��&��o�#b�r��ג�������R�]f�.v|.I�ɕ�wp&�#JKz�+�
�Y2�n+M2s�'4Ęjc	6V�.3���uI��A2��@'�`Nx��yg���'>��%��Bo�R�2Յ��&H�!f��hS �:���P��t�� -	�ύE��],��T�ЇM��ߜ�*�@S�w�+,=kU{�����}��bs唣}�=�����&�r��<Y��C|n��1%�b�ި�x�Vtƙl P��5\_`Ș�WD[���OlB�ܒ��D����r��E ���������i�P���Y�h�Y��A�0[�l@n��͜&���|�KϨ���N�Rq�6�\_�׶0육Ί&\ܟ��>�Վꀚ��
m�P�IV�ɳ�R��"�	�-`]���5R�������v����p�2{�=��g���eC+���:��n	 �F+��p�	f���ن�F��;tUt��3�cϓ� ~ڈ���~��V��.��Pg�0��Hy���^9�������\���A[�~̡a���REx����9�C�9o k�0 o��F!�;T�G_��~ǿY(�����nܔ�(v���Z����fך�jq����)_�R �&�^H��:x��0a��+)����VC4�R��:�&#K�Q������r5/?~�!&*�&�h��*�+2��v���EJ2o��k�=�4k$�lZH�\1��=��Δ(�7�63� d@7���x�����,Ƚ�@�)���k���������OR��u(0�z����o}�7�b2,C�VՁzO����˰�[y�_I��"�@�]1��@y�2]�X�O�����,��ǓUQ0�g��ʞ�G6�,2�m�S���ơ�A�f�ژN��I�Y<�gO!�^OY�d����-��3�ڀ��5���{S���� ��tft�Ȕ걯�f���f�چ��3��}�R i�P����,)�������Z'4�7��c�Qz}*i�Y�^B�M1��A.�WΏ�7[9ڢD-��bFQ��9YJ�>Մ4����D��,���H\�	o���9�y�	!�k�c�����0����rOr��R-G���@�A%�a�M�)���χ���Ս�Aƅ��)��nk#���-i�I��uP����]�G�^٭J����X���[X����V�����5�����M�N(��"��h'^-s�|�(3�I$��$�zV��a,�loϰ�k4_��̲'�Pwk����@@d0�%;Z���/	�%����u��P��(m�����$��Kn���U�|�#M�����99C���4ci��n�e��
��)N��-8�)�u�a�03O�ɖ�2���-]�;+[��6��(��铣r����K���ͦ�yf��ɲП+�
#�w�8\?�;�n���#�\y笉R�`��!b]�JB�"*g�nC�8����Xs�fQ���뵣��a����4�2����Z��>�y	�U�ո��i<cW\լ8!�<҄Q:���	Z��@���P�o4N1D �% =���FJtvV��T``�gŁ�~�EX��;��:П-k�e�	CHh�p�� \Z���]ʊ��}��udt�l��?�r�_<@��u~��:a�x�g�t�Lk̸��!�`�O��D�0�,���m�Im莧����q�n/lY�嬢?b��,H����f���{#�u�-xe��=�2z��x��'��Gݓ��jaS�v������TN��{  �]�8��X�������gF�u��r�Qٛ��^��.��z�s�U2��*f	�}=�
�d*�>)tt��dlWM8��V�D�_& �XN��h��掅^9)���d�"�?]�@.���9����&gjuhﱌ�3�2׭;�L�_�� ��G�U����Q�㳶�Z5�j�
��c�6'��v��A���;`܃\_�̔�>KFs���c�`��`�?��ǐ"y�+m��h�4��3{1궦�La����w���S�������C�2:��`��3~�bڻ�����L�o��0S�@B�3`#�3Ń�Q)�#�����58Z7�6i��b�W�ٮn½b`���|���D�]Ut�X��7mA�fg��-��^[9騼aLE��`Z�Ԯa�5���� �Ŏ˘��hy4���ؽ�h�,=�j�o"�ӭlPi�ѷ��ƥ��-F�q3�K�U�>e�{��pGv��߳�$�X��-+ZF�w@�� �5�l3��*�ұz0G�_���`�6F�s���@��D�k�?'�iMܾ����0��MI�3j,[]wPSuL��<�v���:�W�}G}�Y�4c	�*���%�?G�l�h��M0)���ޘ~cǊ�.�㏔�0Tg�O���nܧ'u�p::b+�0�֗f�	{���Z5���L�9\�g����2�5�H{P�~�H�G����iF�y�\x�6��d�bL��5��Z������ϓm���PG[����⚓v��0㨞�����~��P�+�^k;}�	l~��a� J<��/���w��O��9�� ��>	L��k,`�?��2���tol6�8�4+;�~tO`Jr�-P��Tݧ�Ɲ2T� T3o�jN�yu�������	�� ���%`��NI�R�=�� ��U{����##@nԖ=���tOڭ�Z�Yc�^�����&��J�m��pd�9X߷~϶��@���ή�6��=����e�z�I � �߷e[�_|?HX ��O�)8֕GQ�:D7[.�8'rE��ZO�V�p��/����)'��/G�S��T-zNg{h�D�f�\PA�Q$"�cC3�U*�i��*��-&�0�����ys��\=��/����%e{(�Ja�{�q�e��Dſ����5��8�)d��Z�������	�����f�Ť8oKm��3�%u�����f�c��k ��e^��P�_����hj�	�q��8�;�2%�xJ5&��$p�q�%���Ձ��  :Y�9j!���όjC�:�a8��o�R���ru@��T,�E��4��d����f�Hi�����0#��1_hq���a֙Jd�K,b���=)�iJCzKZU�1�'6E9����6�>��(6�e����d:%f�� �5�R69�.y��O�!"?t*@�L�Z��� �����]��7����H;�� c�:�p8�F�Xѥ��Qo��i�6TMCU}0�jW��6�].�^����<̬��/@Fx�% Xf(x��b|��r�,q9�Ϋ�,Vk^8g��U�v9�.3����k7�K����9o:�O�y�f2�
��չVx��N  ��IDAT�2V4K� ּ�`|k�LhK�Xd5T_�-*@sc�{̷�&��!�G�k�z��Ƿ��Z�u�� ̆)Yy���x	�.������Ϋ�`�/����7߶Z��\���wMk �]�Tj���y�7#Q����K�.גM�抝:��j���Q��v����&<�A��Pc�tI'��=��Ep6*p�ar����Tk $rNU@�^�P�;�bw!��y�}�Sd��W�;����;�P��RY��9��.�z��*e�Y�}�^8?fǿA�)h�5�U ��,��| ��y�+�ރ�V	��R4��O:��=v���Yp�Mo�r��+V�1p����Jn�8:PF��y�y���(���T%X0�{���N�ۮt �7�!jC���}�.Ù�)�TU*\߰�%0ӱ{Uq�ɳEαG�%Ϫ�D�j�����b�X�M�%��T& ìPkYu�Tr������ʥ�]�X�;��<#Aݗ�!eaɫ�=�y����V�Y@jP?>��!sR�o�Q�K��!$ឍ�~����?M����XZV�ߒ5�?����Y)L������u�*��w�ܬt���@�<�c6�e;��痩,��i�@[V��-2�f���(�29��^w}H�u>H ����]�r���]��r[��Ku۪��=j��ڋ\��<�>���Q��7�>V�s$o%=;!-v:>�Y}.[��>���(����^b��U�x�R�*X��]�����a@�f���ʜs�)@u&��RG�u6.��n*V�å����&`��s��qyK�-��ψg��Kշ���\��.�gJ\��,7`Y��V�c��Bo��d�WnZ�u ϶�.�����	�m�)+�����p<��S���bm)S�qTM�	��
�����R�?O�F�i����X
 [�S�SY���$K�%7�J��<�,��K�?9Tj
��y�z1ub�9��<<��l��5Z�l� /�>�VfǪ�-�w#�e���kE�u�fW_�PK����99��h)�������N0g]��ʶrź��W�g8�yNہS����K�J����p�s�6�����+�{՛�0���]٭h�h\����Kn�t�u�����8�@�n��+l2�J=�kڙvɱ�r���l�A̏����2�w��I�չ��)��A��j:�oa��-��*F�W�R��/�I*1�g���R�>9���
*�S���yb��x����E��lц�٧�t�o�a�W�>��N��tA�X��O�m��&��4Ŝ;/ʶ��ԡ��eV�0{qΕ�=�`ۇ���/{Ƃ�j?M�m	�Y,A$?�G,a��3�_)\�~ ��$WK0mcS�_�㛎EV:�)��2�G�UI5��Tqm)D0� �15v$�������0v�\w�y��Pen;I�ۺ��!oSČ�Dӈ����Ԗ�Nl�u#�v�*�2�s�*;Wʂfp�H��㢰�q[��b�5IAhW��U�rS����n�J��+ ������<C�:7��b�G��=p׫����7�K��0'��8��Թ+�J�q����O{Hk�� �=
��}6�g�1ܧԷ=i����*'��/�8돨'���˛�|]P,��X�L+e���$N�[.� �~��t~ܔ�K��z$�9E^���n�1�n�k��L 8�&�`�	�������nԤ(���̗h����Ps�����`�2�v�UG����p��p�,3-����h�hí���|�ra�_�ܭ�w��|��K����{��x�c.�hK��&���,Lf�M<��-���K�u,�?�%�i�����N&�z�c���G3��7�c9�M��sD�F����k�k�y�C�@�(�1��-��V��r����<�!���P�<�J� �+�&���D���� ��ht�C�ϖ�~�<��!y��P�<�J� �+ȶM�~t`�C�[�P�<�J� ԇ<�!��� P�%i!�	VC #w���,��X�k!$�G�u�����[�I����W�q_����}���N{�{�������%�?��#��e��ҾVL�yO�݀jK����q�mX�ss]�.���K�<W	&���Y��{�S�|�+6?��x�y"��"Lw�Q�*n��{��P��5�w�O.��eк '��=d�k��(����0��*]�&��{�H�Kl�~�m��=�g�;�3�C�ƽ{�@yȝ�P�(K���|�CN�Py���e���h�X=�Z� ԇ����z�C~y �C�\I�z���O�5e<c�_Qݿ4ֵ<�sY��޹�'�$���Ӕ���\U���7�d�y����	1��>�!��5�����1-��L�T�\Ͼ&��� c�s�i]�C�K�6��E���Yڣ������s�}
���s���r5�
<�Y�jVc:���� �Xs����?b�yA��8�x2���,e�3~zKۺ+�{��Aq��d�3r��J��o5�8n$4�����x����x^:��wKeؘ�e�>klt�U��cy~J#�$>[���(������8贿uUΎr�qw�\_�`�Ӑg6�%�i�Wf���g���� �Ҟ߮*y�#�P_H�p�ڡ;�|�3������lM�}�2�7�/���ϸH;�xM�%KIl�������&����"��~��Y���=�� j9��9r
���5�=~�=0��~����_y�e��vƋGr����2��ru�����C���*��1ը���6n�	x�V��Mt�������Y�Te
fUϋ�t�|	4��ʧ��H����2��Z��۾-W��ǌ��oޝu��m��)r3����0s�T~@`���"�V��)�����)�3ݣ��#�G��R���=_���c�������6�$�m[�w�����G���ܞ��l�0���g���o�!w$��^�6�����bq���w=�!���aS偕y�C��re��Q])�x�㥜�(ݖ�bAr���_m��-�*����k�o�Kk�˝���cO�ܮ]}���K֒nw��ع_9���̀XF������{����U���w�,�<����8ӏ;�t5o��P���U��<���D'�1���f'��s;y|��k"��#�� ��aN�5��A���б5&�2����a�g;���h�Y��"̲K]7�T����>���w��Y��+*[f�_hD\�������x�k�����Z��;ƊG��<�!��ٽ�P�_E����H�}�v� ԇ<��G��+@}�ER�C��7y�㏗�>�!yȕ��y�Cr%y �C.�������� ԇ<�!��< �!y�C�$7 �K�����w�D��4�r��S�������s ���?��h����oGN�Q�ں6wLè�8II�F��R�n)��q��X�ۅ
ekZߺ ͪ��oE�?WEH�vh}߭�ڼ�O�Sk�+$�e�m2��I���,_�w&��$�������^�&(/��xj���ۿG��ߌ�LrӞv�ɂ!�TƑ���#GH�e[�p/S��jAV�N�;���5{�9K���\,�Nք	� %�}�(a�t"�=�4(�S}>�S��Mj;���9}�������8�b��k,ݿ�.{��O�M�W���˶�R�I/Ny�[��h��7jy\"���+�{����V��������ϝ�>�$��%��|7yHz8�n#�P���L���� �K�d�#e@���<䗓_Pgj���5V=��[ mX)�m?�!�5�T�[[��s�nlA�]A���C����{
�r�T5���mm
�ǿ{�y��C�(�.�fQ���1ru��_J�B�J��p(��EY����<�*��*�e�כ�&l�W��?�!�����w����
���>�!����W�����04>�!�4�>���;ö�xFJ���4s�ĕTe���/N�,�}��v"Iy�|=t0��צ����>���l�]����E�j��`7>k��8�,�s�=�B~�����j:Uh�5��-�dv
r�f����~&^ru@Żc�mj~��(+��tM?p*���{����w-f��~�:���x�k��jD��Yp���L̼����d (���d`�u<�4�ŒI�����D%mlp3��"o7���۽}M�w 7��|~����r�b˾�OT�/$�)!�E�0��&�A�����4�kݘi1?_�1��K�s��~�j��V�Wz:������?��/�{�Q�M��Zi[l���rZ��X��h �Hs�w	7���W;�.]�o;'ދ̆�Z�ĮQ]�HQk��U����rf�� ?��vL�W}�z�?C$[��k��%R �5��5�~������x�4��m9���(w%?��`�,���S���i�E/�mL��P˶>��r�7/��{���ٲ��3=���ju�2�D�ܻ��S~@Šf)�c��=���`*����q�Ƃⳟ1��r����5����A+;�gۭ�傦�ކ�ikN��y��ֽa�,!t��f�\
w�*�4��4�z�jW��샊����ܛ/���d誜���w]},�Ԏ�w,��K�]5g_o�Ս�T�|o}%L��:��K~7�2��O(?�.���SN���-�pwXP�f�n闯����J��޵L3��#{P�}���� U��b�������N�J���<[��E�J�V�����w(�m�2���`z�m�1�����J׎�_����pSIX���PL�pJ�UM���k���g�I�(z�٭T�{�Q�U?�f!jg�w� W4�7���c�i�F�?廫+L��	�䀪c>��A5��r�`J�j5u���8�pz}�7�J ��ٚ��n�֙8hb!6T�y��rY��@�~�hY钪�^6���zΖ�Pը^���y
~5�~��J��O5O}��PM��,��?� KN��?�\�å��IO�y �
.O�傭Hcl���/�9���N�7����v��y����/�^cqU[{� �w�<��`Yxhۅn�^-o���:������j���}+X��Q���}��ٞ�K	;*5�T6��)�x��mM׉�x�<��r�������T�����;�E�t�ö=�l�~d�95�W���X�=t92H���Sw3W��{�z�{�>�	8�8��������1ʺ~{N�N%��=��jSuȹ3FWOE���)Y��r�3�L=�6������r���n�T�5��h�ű��業�gK~�W�_�N�i���퇌��ߴ�ٿoo��w#����9���Z �a�`6-��%�I��OɆ+����*�m�=���S�^�@�R�L�Wm�ڵ*Y�{�Lr%�l���~�{�~������k��݌�V��%/�EPM5�"�]egs�Ƈl,ϥ�}eR8��Й��*מ2�_n�� �<��J���Z5�^�W���WC�U������&��4�KO�0e������ʄ����K(�..�Se_+���mnӠܫ9p������}��s;ǝՂJw�������=r�J�)7{NT��v_r��7:�����+S�!E�bu,��P�ZyT���Sh�T���x��kl�J4���O�ۜN{��S�
�惂�����２61�پ~q�;��/��n��ފ�T��<ԧ
�Lw9���=@��7�P7/cZ�<g�����o���9ЙyS�塤�Đx��?��Ë/���_O���%F�|s3�1Ը��|| ��{�s�~��x���:�t�sm-ljƀE&�r��Ln��HL*�;��V���g�3	j�rm��L}�
^�rA-�o�Y���܇�7ӹ�V�Tc�.5Խ��g������	o��L�����?�*�,)�A�n3)mg���7��.�C�A�\y�ʪ���#s�i�E�Y��~���ʿ�����0F]U�u���{k�bN�sg��N���\�{c���;�*�I~Ǌ� ��K���ݵ�mw�W�`�������5
����c��c6m�&�|����� ���v]���O�s-��~~���?s���J����X�Ȗ��s[�n��ݺ��+��D�-�K]�*����ru@5[M���s���6]2����5�4�4�o�q�3�/xӖT�sO�i��'�T��k޸G���{��|���7h������eH���k%m��U8n�E�uY��^��;ɠĘ�!3�[Q
1��V��)�9��#�b��p�
��A�͟�t�T�'�+�Z����t,#9T��l��;�U�ڛfq~�~�/|����O��7'�y�_���u]�]�Als��]�U��^�V���qB��w���ƥz�����7g#+��.[�MH�rtyZ���m3��A�Yy��f{^����`�����y�k5s�J��o��]��
�)�1"��_'�y%�z*C�$)�a`��s/�#C�A��
�� �b�̒�h�-��oe3R\�׀L��6�� ѻ/?��0�is��������� �~�z̨��z���+��-�Jkg�$����7Q!uA���	_;Hm����&���� ���V2�Sq�\M��-]1oŊ|�J)�%�0N�{J��:iuK�n��{ x�(�8����;��VY�nbC�3/ %�����N��=��6hf�T7؊�`i�0e��81@Fi�
���ܭ�bg��_b��uY�Oˆ�垅�o�9�i�X�7.����*�B����(a�6���0TE��~J20�l j����^�°����-N��="6DU?N$ݤ��Aj���������%W�%�)%Tf2�J�,W*T��6Nflt�b���K�$�^���E�^G,o�NP҄��cT�=� 3[g��nen���k1�L�@DY��U�ΗZ�y癉 '�M�3��lỶ�VE*.��
��؞�}��rm{��c{�	���v5��^��j_k����)����O�걵��__n��/�L,Յ*��f�ʪvX�k�ca��Wys�^�����V�Y�hQY�=�C|6ǹj��{��^�iqd��:&�0����ڽ�r�H�I6�3��^v�*g��n�%E�.!֔���)N��*���5�h[�������iE�~Z����3��h4*S�+��|	�s�}�ِ����&���bZ�5���F{�h��L�4��.1@����u�Ճ%��U���{�d�*�vkW��V��0��pk�yejm���1P|�[y��-iv%���s����$>f]φ�2�z�fbZ ��%ҫTc�rj;z�]ƾ><st��L����p�X�l��$F�&���>���$�U�@6�
NmJ0-�U�qC��C�zU�]N��JPn%?lO)�Ե��>#��rj�^��ޙS�j[ j1>�cX�sg��Ċ�V&��f��7��|mӛ_u�w1Z��j
_�7 x���Vj���{+��1�/S����x�����p򲭮~���"��d�'���ˢ�r�*�EB�4\:�YT����j?�ڟK�Jhu?�����u����62J,��,��N�U��`���=�(+ξ��i�1���Y)��BS�p�2G#�X!�Y1����e�聵�ߜ���B�����#���g�Y�5H_�C_��±��Kb�S�'��ݓS��Zcv�L��?j�QJ:1e{�ʦ����ab��p��ޥ�l�E�)��{W�M3�c	���8���f �90�h"�SN�������P 68R�Ylp�%�J#����y,�VY���XI.�鉧6f[rj��Ti?,�J����-Q�#��rQ^;z�Mp�n���[��vM$���o_S�{ͣ/`��M���]���/���g{W=��Q��x�	d���w��nEċ��p0�v
�儺��.k����)�� ��_"&�`��Μ��E)9�l�Rņw���G�ٙ���g�yߵx���x����uK�mb�=lr�_�x^�TZ;�-��:&��S��[��'��P;�������S1x�z^�@�u�H���i�ur�>�Mq�6&���Ѣ"��E[���nǓ3Q�����?�<�����9����K�k����U� 6���:O�d��-$��8T���X��f����"�:�"�bEFw���R��u���6A�k뛭��D���.Y�3��� h�k�s�k
��;ܥ�ί�1��;=��ťo�wu�,	H��F��mQ�K�N�%����Z(���Ѷ��������m��{��s���1j�����_6�o�/�8�����Yè*-�:N�O7��]|D�ޑ�^5�Y:zR@��~f�8)Y��ɒ���:�����}��i��P1��[��K�\�Nۋ6杣�a"�B�9g��Ǥ��C�������TZ38��Z��jn��>�t�Lא�kT�m�l��-����gX��N>�%�?W2X��W+��v�y�n��j�HbYY��;6U.�$�#��1T��(/�XR�XL�����̀]}�6�{^�ާ~�O����'���L��d�����zw"h|a��/��R�x�=s����ԝ^x7U�@@9�ӉڤWv��1��������V'@mXf��B���|�e7��Ap��"�S;#3����`��`1Cu���n���P;�(sRc}j�gi��"����Ń��M�>i��;Q���n϶�.7��`�!c���q��*�����͹��IT�K���Pն��#B�SP���tZ����S����LM�����mS��q=~h9|;�KI[t�2Ɍ`�2��T���K����1i�d�|������;)|i�]��"��1m�Xa���<��X����'Vie��i5T�I?`|�ygV��K��,=�Nޛ�7݃LG��H�u�ÿ�������{p{Ѹ"��B#!����2�A��PL�Ts�Y�+���Q��n����:�Q=��~]0M��B��D*p�Fji�l�,��K�L�6�����9�S����� �ǯp���E����2j����_�<t�;k鳙.�A�!'Vf�=���6C/��3Ry@M���Ax,���pH����<���?M*և�~��k-�:��՛����|��gf#2���t�U�N��E@�\��(b@�op�&� !4���N�B;I�If�dv��A;+�ȀO
�]W-��9Z?��T�שnILt"����8��͌1=��]b��I�=�x8�o�]�zu �VS[�v����L��0��e�l��	y�M���m}m��J�:N����G��S9���Qzn'�<�c?����^�uT.[�uR�<G" G���t��:���S����'~gN�B}�j��˞x���Y)�)�� G�1�b0����+)��b`cJUV�` ��͠��uʰ@r�H��Ri���)�ԧ;�����ej*����UL�v��,�P/*{9@�ޣ��uߘA�1.f��'<�b
�=U�9+Ux/���e��S��G�O�I�f ����Ϊ��ۉ<%c:�����>f�F��ji*K���O	<x��	{=l���KW�X_����<P��!&'3-tV��S�5�G��/��'�s��Ͽ�fh'e���S��NI_�~�"fJ��p����k�=�_�u1� �O��Dm�VHE��po��V;!s�"����Ƒ�`_H����x�U��1��J�FuL����K��:���/L$Q�����H�8��i������<�i�' e�����њ����:N)�1uff��bM�H�zrVg��'�y�,3� ����H�WE�d���-�:MFS�"�-ZJ>���t�'�1)��1�'d�,�s:�O�ϣ�˘,!ʪ� �����}�ԌтiT��A!�6T�We���Z6�Z������~N���29�<��ʷR�ɂefe�V�C��`E�l�W+�����ږ�� 2_uu�:CF7���`=BA���MM|�=]��[ީs3Cv`5���� ���jh�L ���@�nd5���4���L�Y���;��Od�e%*.ݏ@��@�ߑ��̠*�4��YY���:Qa��q)�G�{�Y�B_Y`�Ӏߏ�%�Jϳ\T�T�S=9�t�Dՙ�i7�3�ɩ�r�����Ď�IK��YU;�J�_�r@T-Ț����Tv�=��n���D@���lIr�M?�1Tv���gö�"����{�.��!m� �5��1)CS���J:���{1϶=ل;�Q]�*�ݙ�cp<{a�P��FV�T�Wd�v�>h�+q�]��*��~���h�$�D�}�
f
餍Q�Ŗ�f��1O�����\_��gQGɼ���=L,���Kzy�:ϑ���z�	+�M ��I�'@=���j����>R�m��I5��t������LD<�j�S^������kQE�%Q}RY_մBB��k�@�&-�y@���X�bb�>��ebv���'}{�����B������N>||�q�晃Nt��_4*a�)�&��?O��c� ��4Oi&_�|M���O.׷o����ʦ���}�u�O?�?p{�S��z��������v�I��ǍS���B�;5wd��H�r�7���Or��)��3�4w��l����_�Ec݅��Ħ�msb>��j�i�tl�Y՗��S��&�Fx��t��F�_���� >jP`K��QmP,P����V�Z������hvP��g옹�`Š��Zj$���e��zF���#��U�Q���:*�G��C���<=?M�{XT�d{a`�ze�%�Fd��%'���~�2Ӭ�@������۽h�����g�������N@��:u����q�?�s��gg8��8�8�������ӧOʢv��V�u�6���|�NNj�V~}R36���2�:V��f�O?�u����`O�����"�3Y�e�w�Ug�B�Ea���LJ|�h\p�����
���]����4A�
�����}��y�ݙ�Wڷ$����	��yO��J���4�rL*� h�N�Q� �Q3Nň�-�:6�P�E�v�����������1�:��0�����g�I��Κd���6GU�z���%yMpF��Ҁ�Y�U�]=$����Hਃ#�MU�eeO>(O�;L�Qfΐ� ��1.ϩ��C^�S�XToA!�qfk�NK8z�p����qޫ��P �X�_�-vou����;�8¶:�T�^@�8�>�
b䤙�)�;�}w�^�?h�Щi�h�X�T�Ԩ���I
�x�S�$}�[�:��cG�ij?b��v�z�`a��q��#���%}��=awO��5�oFSOe�oB�|�TqbudW5�e/m���$u��{�eA��j�0�؏�l�����R�%Em	�WR��i�=O�[8Tx�5��P�$���4���y0rz��Nl�$=Ox��������noe����x}�����_�k�M�Kjw��`T����L���s�r�2�i�P�ډ���<u��(`��FG�z���胛%�����*�&�kϝ򩲋yG�ꜚS��<�<`z3�[8�(�@�~؆��B��B�"ḻxN��0!���+����PE�g�~J�@5|	6e��̩}'�aI*�� �46�^�1o��D�w�"�n|����7V/���������f90�]B6�����R��zB�A�T��Q���=��v�Ws�*���b(�l|j]!�S�% ���.WOѯ�7��p��`�D.\�?���(�P6��w�Ol���6ޤ�(i_�-�Ɲ{c��7܆\��ã��hl�ɖKQ?�L@0_�3��Ii�:��?�d@�?;zu�a3Mӽ�S�Q�xK���Nm4|U#�Z7���5(��C藩2���5}�T�#��ԉP�]P4(F`���
I<�I]�?O��3ٓ�RJ9d�C���P9;���es����y�f��.�Q8�0��2�3��tQ�^r���GMn���F�]�	/X�@� �j�Ҹ�81�f�KB� �:�~-u��Hz]C���X71e3TfR�	��}.�O*1]���A��5���6&;���߮s�;�y|�������۱�!]p�I;~8#��,��(8�]�Y�HT�[����4�G�w%i�[�r�����o
;���R��������I���B+tv*�כ�A�<Yy�nEՂ�'=��\�کN��ݑME9'�b�~�	��&9����B �g���A��F��ҏ�⓲*�!ZHW�+��ڱ���J�N��_S�~�@��ǺIE@-���D�	T����C�܈�'	����
�}p�� �8K��]�E����F��+�s�pF��L-@¦Fc3�>�D�a����!�8ry;�n'e	��4g{���Z`]8^�
&�$��f����NT&V��"K� =��?��ZtrBQ`?n�����v�Ѽ���d�����$�LU�md> '��K�~����y��o� NF8���q,>�4���Nb��\WM��K8�2t���N ���*&(�'" ���;�U���^dBRG�j�`�R��ۙ�	��ݢl��Z�o��x�a��#$��cRME�����>z����n԰K�9�ǍE@<B�x���m}�Rؔ�J��ԡ� Mqe_H5���T��沍Lla�����$e��$��p�����U�;zJ��d�NW�P��h,�'��Bm&�A�ଢ଼w�ٳz���Ǔ�z>1�$1�B�S�1�'g�)���_��Y�������r����}�Z'�N2�9$L�xՊօ��Q�B�+qr-�āU�F�k߄w+�k�������1����T`��~bL9�}����~(;�Y��J-:�Ϋ�X\������������D�������LB�ѵG5x�)Έ���D1ƨ,W�≏�▟�����+#"�)=��P��|���Sb�-�N��L�d������C����u��ȶ��//LȄX��C`J[�&���XB�LJ;�s>�_C���?��"�� �5�K�#�59�eJg5lT1�\�~�X>]����1}4�I-eUK-{v���A��=5��WЈ��;�46���y�zBh>#x��Q�a�b��̋����S�/G,~]��Le�I�z0�� L`��=d8L��0�0p#�r[�"b���Q�'?�ϻ#F��=�J,�ep���Ӱ�4�M !���������r=����D�Ղ�|�@��W'�5p�Af�X��t��m<���<q�P��e� ���1���LE�<�qx��{��a!z���]�]�y�V��~�@�� +CF����A��L><�4(Y-F�&i��M ͓ �hv����X�c{{a�x����{�m�r��RhD|�ٷd��X8:�u�Yl���t��$od���|�x��	\�b��Y��*5ƿ�5���\�"�_fG�֎Wݨ��\_�.k�����vi����RI������BdERg*?�(L	c*!�y��z�S���:f������ ������ޖ\���&L�m���c,�Dk4xr�<Tj*Xu�:7��x��۱y��18sR��T�g��6�~�N�D[;�g�\���u37���E�V׫��Y
�[���u�.��f7�����󈉲x��1E��;�������������lYl�c�T����9����������[���JH�=��2�~}c����;!i�8�h�}��,A�s.M㒢?^_���`�QS�z�az#P����7�@NC!9C�0�Q�����חW��']VO�th^�1�����q,�+{�ɾ��l��-jtz(��;���*+�tR��S�O��������ET�v:��' zzڥ��ӧ�n)�頁�$��Bx^���M+gN��ꎲ�آYمih%����f���<�����V]#����<u�8���-��� aG�L8^���݃�I�H�|�_)��Յ�U����&��uv�FeF`�sZ����F`�wV�L�,;gaﯔ��K+����V^Z��U��9���/�6��&u���;%VH�[J�8aρ���	y(T�?������E������~�������P�ΰQ�tq�����ǀà�|�c��s�ؠ��s��I��v/BZ�����������6)�t?
��������ҤD�A��HW��%�C���F��>���9mac3{�Q�Ti��C+b���*���7aIA��:�o/~���$�Y��q�'P�z����K� *�E;]~8L�D+Lv�=>���Uc4��9�|'K��C�4��̣jS~�T6@��e`�qq���dC�KZh������1i����f��lp7l�7�� ;vf� a��ⵍ�ƛՀ@�e���:��r}�w�L�񹣩4L}	ͺ�Ԟ�:�����f��ó-����c����%5����?�$}�򒎼
p�+�TC�'���k�l���<ǔRj��ɲ�5Z'N<1%��K1�P� "(+!�2���f#��bap2��-���6�*WM��3T�0C�Xh�����HHu'`$O�d�dE�(��3/)���F)��=�K���yH&���;��n)��auU�Ӭ��+���J���1;�(,ZL�a�L�L��Yųc�� �dUX���u����j�)I��J�]��2:��f�UX�g��N�i;������i��iq�����+:ۙy$禓C��4���@k�US��W��f�:AT�6f��ZXC��"� �rEY�f��,��33/�ռ61�2~e0# ��>=}H�U�{�S��qJ��ŋU�$��b1��Tl�b��i?�Z%9�"�]2��$Y�^���%e;/�����%���ԧ[�U�@�����и���ҥ��-b�]�f�2��I���.Y�����M������E��(��l����A��hI*����	�MlH����=�j,�d�#;��ç�y�,��}�'�����N�]�<ˉQf��`���
h¹歯e[:�=t�O[n@�A �8XF�� �O�y�,'|�&�e�\aW�S(o��L�DĲvh����Ѱ~��xU`'v�As���BTlR��<�����?�O�P���d�c׽��X쒎Y�?}d߃���;O�(��0�{��l�D���zه�Ê/�e�H�Lk��o�
t]�.CM�� �/f�!�Xz�ه�	��N��_!;LR��g���"�=edE�4��̈yſ�=i�y-nOgHT$���{QN�����Q�>J��ab�̲�Z� TJ�֌���?Jy*v���nBY8��Ճ?�@� ��3�ce�u�c|�+��m�P�U٢-1���m��8�Xj��J�ID@u�c�}_��R����X�� �c޾+�Wz�kH�Z������U�y�~ر�]��k�Umh���sJ�+�
��K�-�Ė��r�� Zp�?娙��M��_����n'�*�^�+�2]�#K#B�˘�6�\�o�U�@���=|���h'�D%��B9Α���2�Ny8N�fT�Ȝ�������f�AV�dK7��9Vn�	�������C�d�;&d�P��cO�x�%��G�3�*�uV/�8���L�+�-��jZB�\/�=�����: W�h*Ŗ��|���s�ņ��i��*�/QM��(C-�K�h�Y/��'LT������5�deͤ�چK�[3�l�� �����V���?�W�C��!¦d�� �Iw��QrHR9���rHKH*:�Q1.����1S$��n��,	̞�����?d�kZI*]������{"G�d������"-rߋI�������Hn�x]�
��?�:H6�2J��0�,�վBd���W	u�@d
@g;�4�d�Jd/�hd >~��wz)�
3(��=!Ϣ��W��z��1/����oNt�{��l�%�2���CY��f���~T�MNr-³��zk������ߕ���}*Y]J��F;ހȀV=n���<�4�}*��GV��RW̜�ڡ�Q�9:�͙�	Ydƭ4�ZT=yv�l�s�'�쑗��E���^L�Qw����] L#QF���?��o�E�J��Z��3PG���||�\��~�𤌷�c����������ͱ 1˄#O�<1�>,mpBʶ���r@�ؿ�[EԌn��N�jlʑ��_�R��Ybx5ϑ��R��xm򷗯��GYCNy���L6��PC̙�������� ���*	���i��r�^��eJ�3�c�r���<��`��1+-���'����ȹbSs��njNX]ֿo��n�kN j�ٽ4���j��-�����>1E�����<{]{�X���3��)���\��m����-�ޚy'] �Ʀ8���>��{\�AU�#���S1ڸ�R|�#vi2��tO��ƚ`�����c�9�u
s����C<ÁA5w�C.�`K�D��������0g��^�����e�53	k���ƑArL/���?�Ⱙ���^�D�|�SE�9���?=�/_'�:(y��A�s���b5el�������t�US�qPzv�y�-�3 Ld� �Q�dE�LĞiq �R�N�Z ����Ύ9,��y�Z<>W�k��[�jO��Ug�$�޵3�s�"��}/)��ݒ=�=�-P���T楺��+�B�W&�Ef�P�ZV��.	�w5an��P&7�{��L�� �=�"�H��~�ʌ��D_��L ����C���z0�j;�"'cb8����O���%$G`;]L��9CG�3̑�+&�����0Fc����u 5g�}	�U{���Nͳ�Af+�A���h�%NP9G�X���ub�d�κ�VNH�BL�bP�؍,�j
�EXY��Z�ʺvJ���=�)︣,�����ꨡ�d��dEPQ5�%�y!��b�CF����amB�Ll<�-s)k ����f���|����P`�h�Ԃ�'a��|*we[��}�Gv� ��4���s��b�Q�+��^���k��~�,��%@p��2n&Nh����7�W�܏����r0&J ��$��$�~���=�a+��Ϣ6�$�U�Q�&��-m�:t/��v)�&[t2�iOU���L�S~��t�Y=.�����z�m�IP6��T����>/���{��Q���0Ԣj�4�M
�Z^��1�m5��U��$"��yV�Fq�X@�+V|Q-F%��:����-܎g�QRڨ���e�ɂ�1��d��d(ҐO���2�{����k�:k�PK)��%�o�ɏ���A�©Jd��	�Cd$�-8.���5\fn�I���l�i��&	 X�����ʯ�h��u�6x���L�J�׾���cx�ɫOI��4���J���D'Yl���*f8�I�X�)9�R[���5�f��H�-	��d�G��������������q��)�v���0��`Wc�8�M�1�H�t<D��G���:��/E5"�]�%c?�%4jH�����S~����0m��1l�F�2�Bɣ�`|?�v!�ؙ���=za�e\T�|js}���(���
LW�+0m���P��G��:Q��*�7ٷ�O��B�3��f�R�AN�
�f�3�
]�p~}���*����c~�ۄ�k�JyG��Jc�������_�E�mDZ���:dl�-�u%;���yl� G_�&y�1���+eՏ"99twhpIQv���?��H�M" N�RƴOHш|��L��u-R�:��K�rо�^iO)���v�ݎ+�¤${=E�8��|�3Z%w��WU#�!:^�tx-�Uf��h6��A>�Ƽ�t�e��FX�G9�*�|���3����#�2`�����>C�~ݥ#X�fґ���L39eБ-M�4Ц0���ٌ=��go������f��{T��%�v��V'宿�91؟3oU(���y/,i�����"�E�{�ؿP>gD5.���@O9� Dx��)��	j���՟���Ǚ%"-��;"Q����{�]��=gc#����Q����0&�k�I"^F�L�m� �F�ħ�T�����xԭҳ%��q��'��V?������y����W
�z���5�����(U2�Z1�X��Q�+r���q��S�#R1�!���z%/?�������a�9NQ����{��}���]l���Ӑ�����G�v�K<Ӟm:� E��Q{I8D�{>|Jm7J�5(5�]��D⅗����NA��AT��gSw�~�����_�}Sv�M��W��u�<�}��YL���ߧ�*G1��Tt�R<�s���4z�Z���sLr��XT%�������KO��~~�Ry���
o��x�)!�Ų"�6���q�kS���jտ�4��mGJ!R?"������6����Ӿߩ�*r7���l�:!�5{�b۸	�	�kHN�2&X�2��o?����ǟ�bO�[��!l ;p�M�4%8_�#�Tt��t�2v�0��]�aR��������b��h?���i��ˁ�9�4�@v� ���(eӐG�A�S�o�GX���2x��j���>��\I�^�l1O���T���Hѽcl��!M���WD��=��;�����ʤ���$l�#cy�К��X�T��jw��R� ������vL-76��� Y�'eC�d7��Ē1�9u|�M��׿����)�U%������#wB�Aܶ�)0���s�u������fV�'׸��^�g���U��,)��A���d��\=�)�����]"�9���`dLpi=�Rd�:Ɠ�KdB �"�=*�3 䜁9 �����$5Ř�qAGv��be�F�.��J���ݣ���ҿ��21T��堲C1�esH�1a90���=6a���7���X��c���c��ɎH�X4�G^8n�#�Q�1���D�4������¡^�!ݵ��� {*�C.�b(�;�e�ǥ��Tr:b[^�Y�u϶Pn̲�F�uf�x9����A�f�B��}P�TU������f��*�X��[�3!ލ:mu,�� ���1zEwH=u�v�";X� |����1-2Ј�Us�t���� �WU6Y*3�=	�Y��N8.- |��Lxp*s�3X����0�'u�qv������%�"3�����.N홓�p��Ž�8���`*�D������ ����{Y=8�����M";$��my�0��9�ٷ�A��+`��6��c���cN�Q�m	��F#j�6(	Υ��@����PS5��E`�Yr������y����B�bQ��8��.1�#�s�~�َt`�t+߂�3:eGR�}ll哂�y�qy7FݤZ~eC��<0b�'P�z�:��9,[N�!^V�Px�0���Ub�<�skj��<�m_9l�K׿��D���l���:d�P��F��	{���aV�PΊ��ok�c�R�4&&/%�2O������$l����U*оʶ��v�sF$��,? J��\좴8�?�H������P��Ǐ�x�a�4�o�M�:�Ԍ	���JY��o��k)1�q��j���w`��飏O۱�F�O,}ͥk�������f�qi�-��9�So��&Yg����@��{1\K��vE4��ԳNl��d���f~d;%peU�*�z�aH�ҍ�%5�K��}�Gt�ʃw�=�G�%@�������>}���}�N����w=eu[��Z��5y�G�L2���7���� ��K�S@��b�i�}L��$
�ın|����8�V2 a[��"Ȱ��lvϢk��?�i-^�H�ubˋ{|��4��Z��9����_릕�pt�{�?�:��A�m�MKF�}���M������_��O�N�me��#�n��0d.x�I���=�V�X����TM<�����ۛ���Q+�MAEw΀]��.��_ƪ��"U\=�vh�+W
��PTW�FY�R�b�ˁ������1Ҋ������; ڣdω��� ����d�|L�@Z�V�`UsZ����8zEPyċ�M=���w������Ug뜥�y��qH����_���� fڬ�u�������2%�<� (_|B�U8a�P�*�RtɡP�	��M�O��R�Ez��2�.�$YT�=a��*���EU9.�u��Z�S��t��՟å����4�-N�+ 4A�T�Q�9�)����?m#����	�ߔE�8Ȼ
s��N�t5hQ$u%"nl+�$`�	l�7��<��D~̄���73@�����l�U�'GW�\G�DŦ�cY����\5*: ���,5&��E��.*� w��W��j<^:ZTm�?����P��P�0M(v~l��v�l��S{݁����c��o��9[��>�K�/�E��R,��o���e����lqvl���1��
%�@����vn3�q����M�s���FP�R�_�}s`��AcO&78��jf,3gۿ�z�]�$��=��	��e\dt<�qOo)�����I'W:�����,��z���X]$Ri#&�"��k����/ {9L�����*�����:iy-Jr��H�"%7G,�Ge��<T�������ڒ�)!g�_�6Uy����������P�[��	c�� �*���I�\�j`Q�}T�ql����QJ���u��K�c�]�N9�󇷴/{ߑ�x�$�������li�(�����Y�!g��J��(���c�v�%�	n#���]H؆Γn˒4	���P��=x$�`g�.4|�	a)α�U�<����Y�4��;�Z������L�l��~���P�1UfsF5abՀп;���m@$s`�	�j_=�J����,����̡�|5O��˸0�hQݟ�ڒ٦T�'?���I��N ��,=��z]�P�����_e3L�,����y���M����y�xl�L�&:6s�=ۨ釖i3c����j1DRm�v�P/�_��e�d7oDR��*�߂�lP��t�|��$ 0+���1���{�&R� �S��>:�S�VR��j.[B���$�����i�b�G������f,5��LptE$<�̜G1�8�d�!�e����?���v4�ȋ:'F[�Uǝj�ڠ�Э���B��q�50�fe���Z}�qo ��R�,�(;��qc�nF��0��{v�ו5T��&�F�#�b��QRF/������9�!C���R����*޴��"P�iU;ٍ�h)4%	��N<�K�-���
p{��&�8/F��x=�"��
S-ԓ�y�ԯ�U�Ϛ{�ۗ���y�>N���[,��b�n�yE�t�	��8��gב,�j�����q�R>T,+��S�T@�>}|N�������((��������%�$����7ǘ�E�L��2�^�.��}�����s,vpT�Em`I�Bglɖ%��4�C��2y�&�컇Fo&¥^yC�Qٮ0�A���3�)ոU�f�+c[#��;�;�j�\4}���,���ֹ�ktC�<��H`<:SA��Rd ��T㱣��=�rr6#'��呂�RN��J��oU�B 	�;lT�/��lҲ�[��7h�O�jB���/)�ʩ�~ߛ66z���?c��!�4��bs���L!)U��8�(%ff��+WҸ���)�NX���[s�a����{��T�����1%���=n���Z�u�1� |Щu�#&ApN(�,^�c�t[�N~���'�?�`��;� �a�W�`�࠲�N���R���`�Ps	�$���( �@Y!�j�@��8�8CV2�uE}��]k��w�z�ꍗ��s��E���I�g;����k�x@�N20I�Х��F� ����j�]3�ǔ�u�2N�-�*%c�E�(��N0������K��Ǥ��\}7���똳~�E3j����VS�DE@�͡_Y�A�����%�hҝA�3����ޝ��u
pq�A&u7�ѳ��Z�5���f�� ��,��64��1G�CA�EYZ?y�f�2.6�<�!�R�W 5��mt;�\��y�I81^�;
���d�������������o/_$�>'ya�AR��X���3�0���_���!�zZ��6{
T�$��q��sA������s������9SU�ζ�.�0l�v��QY ��R���)	��|���f�ޛ�=�qR�2��2d�D*��9IW>�_e a`��b�8%��0U���j�27u$B�N:@��KamA�8��� t����ΣI��Q�33m��q����Ef�&�,�n71Tsfg�ΐ�TS�� 3���}�WLJ�2��ƚT;8j⑤m�K��z?Y6ʝ��&0T��q_�[+�ـW�]���I��8Σ&_э�ƜC;��l�)��Nѣ�s���՜RF
���C�(�� /_�������~�"u����矶�N���=H���t?b������f��=f�����#y'[���x#UB@>���:�}`j)��z��+,ԅ�}g��A3p!*w��;Z|���'�Q�R���b��� 9[�,d,o5���d�0#UK��{#|�w%M�� ����w��A`�Ksp`rR����ź�&� V�	qF8>d�c~r��Y�����)ۤh F�[B�z�4	s�H�����|�&i#�g��5�.b=����a��+�T;+�~g
}���*�,�V�t��rOp{�w	ˣ=
������Wh-2�Kj���/ʀV�y�;ԏ�^ڝsb(��f�Pb�2¯$�`4�����k7ה�{�ͳ������AC7(	m1+k���KJ�N,�ö϶v���d
�͂�}�/T�&�B<�/��Q}P�1�����)���4�ai�S�p��Y�6�B����NR r��,f��A�7VU�V�%�X�.xyXǦ+G���b�z� �;{v��y�yx�Zʉct{��d3�/'��&F�YV8JF�:��j�33Q��<I�mu;�nj�w��5�8`�hQr(�A��=]o1��4]V[�r�ɻX�M&����7���.���m�x'������P6;j+Ʀ����A��J)Y��k�h�!y^o���H���Q��0'ڗh���!ܯ��f?��,��$ ~�����k�����1T��vu�*��U�-���,�-��
��\Z��J�s���j���F����N���t�\�|��l[՜�#�&[dB�K&��t�ۅ�~�% �A6�T���	�k�w�B�l�NV�F � }��z[�"���V*9u�^ى66kK<��vz�2�֑m�;�n����W��1!@��N��h��1GD�h��H���ʾ4���Xof�\�M<
!hsxxȘ0��)�F�/b�|��xZ��i�i��q0�ds:*Sۅ�d�4A{6��y�d`@�]Vf&$d&�&���S*�bdA��ٽ�E�1�H9���x0ٱiL��\��W�)0=`,�*���e˦���&��J㤭L4)%�ޮLEs��L����CM)����N���~$�yg�Z������"k���B���U�QUS�R����N���Y���^�`e��\�]ڕ����7���Ւ:�����bL&t�R�d�xL�(��9��M�������ó՛�<����҄��r��ng�s������?���Q\R�{����*��h�U�l ˙�leö��cl}�����p؛m0��\�$�݇�w�B_�@��2��_`��EPUe]{�������$�b:hRO�3Ϯ��]!���u�
N�X,�i	al��JE�w�I_�F������qp��ɪ!@�X9e5�V�_-X��~c6f��l-� �u�*yP{(���)�}�Cm�ooY�Ý������1�7��Ī%\_�y-�f��-F4TV�h��K\wb��A@��t9��z���A�u|���~�CπÁl���*����o�W������z;��$�(��&�'�� ���������:��(�`!�<��j�x�M�O|���MP�RRU���	�'�,�a�i����.:����̪ሔs��V���Ȓ��v��M��r��qe�	�~ gL�0	`���NV8�E��s����Q���R�o�����#��q����@\��*L�1������y4��h�1��ץ%����&X�6V�G��0�4�\E�6�Paf*O��`3`BJ�Q7��9{�\#*�1��:x�Cfs��B�^N���JܸL�ZJ�܏������������O�>3���tK���?뻒�8:�M����k5mڠ^tN�ۃ��w n8�}'՝��S*�>�頵�i�C5��BFNu�$ӝ�ERf2PN[�=,��L�ň� P��I�(w��*�J�#{�]�L*`�����n ��������͓�R����We����NMtoPǉy����n����+p�j?@tIo���OO��?�i�/`��C�f�xW��puZ���Rߝ�C��O�>�q��J���!��cB����>�c"����R4�u��H��dc�ը��(7�@$�e�q"�ŉ��
��^4 02�+��j ��E�]��"��WU{Դ~�(����u�.� 2cr	��^㬔�s���^VI�B*���GY��C��� `o*����ͬA� c�8U�.}����ExG�����{�,;�(��� �/1<����1�D��$�0����nW�e�w��F�3Q�;�:�d�+x!Ѩ�3*�|����JVJ�ڊx�Mu���\�Q��w�wN����[�yX���V��'c1��OV�$Tw{]���hx�/}yǎD������J╖�9��Avr`mb�z'8j+���yO�j�f�Q�.bvJ��.q����<��.h��v�m�)�=��%Y ?L�����7�6���9i<�F0T؝6x����\�����eae!���[�U������,A�R�A�����<�I�$��=옝`�)�S���!@��!{�NS�A�#֙[��9�i���Фo�X�\���&�0��<�e����SPM�:��!�%�'XL�̳X���eo�;o�B�w�4j�\!���*?�{�!h�yb�"Il���f�p�Mw����'c�X�@B��:Fٳ���b��	K�x�M�z�s�5LLm���d�c�2�@N��������Z&��Xm����4�������c&��4�A���S;ӷWJ���T'�S�~���~�>�L׉������;�.v�	x>bZ&�`z�p�^C���{4��9�3��%l��tJ>	h�G��-���P!2T�5ɋX�p,:����q�˟����ܻU��Tb&��aVʁ���-�غ��}n�܆u-�o&|N�Pe����_�:L�*
�0u5y2ah%���YR3CHꗝ�0iu��k���Z�������NUttDs\(�����Q���Gw>)��tŠ�P�ua�"7�����n<R��pLX����H���!�v{zy2���ާg���v�1/0�\��1,�����>'Th�+X}��rzi'\���%@�G���ᅳ�w�ٙ��M7Y&��F��!L*�Q���E�x��%��1sb�����o�ٳ/��+��1���w
	�2v�'�bS	�L?��_$��Q�O|{��&"[�\0�gj��mD؆6��@u[$�:��*U_��>�C0~�0+���d ��ql�c�] z��(h�[�����p��Zfz.K*ȗ�E�o)���kc�̓*`u�^TF�a=�m)(�0v{�m5�����X^�i��\r�X��Pl��5z�FR�(͚��a�e�4�D
�X�u&�*[OcQEvw���R���*�Wʫmu8*�p5Yx\ՅU4������j7E��,\f�m�����8�`we����*o��	ɇG�+S�e�ϲ�A��;[8���#�<�l��}WTYgB%���ʮ��ۇ���E��S��Xꓪ��d�$����H$.[��LrŲ�1�Cx'yg6�M��<������Eˑ�M�Ꝟsz����LuUe�K�	\��F�Kr)2�&�顗��ˋ�6T:hA��,v�i���l�W�V�!`Es��բ>�>��U��q��~x)I\~�^�����W���$���������(`�!*0��t_z�F���P��*v<ƚt���ύ�Qj�\j�U�V�E���r
&Et`��A�ׯ�w_D�� �����]���V[k&����׶S��W3�����C����b �, |���&hӻ�JE$��D�.n��á���^�Mۢ�{_}߮�,o]$>��\���XFO�$N���;��T�5P���!K%�w,�}����.E�T�Q7�-��0�	0���(�cˬ��ܫ�� �{�۽����-�Y��(ʊ[^��?��u����z[��d��o�?�����xK?
�1�f�͞���3��t��s��:Y�SË�bK�I̅�omѦ�OLC�g��@��G���*�Z��
�$��ׂ��\�ye�n���8cz]z�Q*���oZi�m��b�VX��hv�B���G!���8�*+kP�*mԊm���>�9;k�Cǘ�r<S�2Qy��Dy�����Ō�n��f���[��|���f�ySd.).� �]�Iy�n��V��:�Vs좛n�h�;�:�U��1�2� �2ෳ�4r������W��s��������_�>�/M"��F8�YQ�}��D.�A��yI.B��L�DO�����/��e�ì�
$oj�kƘ��ݷs��7 k��C�Y�5�k���������{<���}L������1���H=Η{�`����^�溄@�I�ԞS���'趿���_��}ۀ�`�Zl�Svc�"�{������'.p�N�������?{0�w�C�]0���TU�WXkD�oi)��Di������l���p ��A5\��Ď*'_�8����-l��� kd�W3_�Ѿ���]M�t/�� х@�#U����;D��-���תbaԠjE4�_-��ڤ�Z(���I��Q7κi�_s{WV�����!ت�4�ݒZMao�сB����dn_o�5�ec@G�X*���W~�!���¤�b0)�E� �c��-�E��-bBT�;�zO��ئxZ|1�I}ׁmᴅG�N}g܁�1��R#�h�֬�}=D�9ۥ�r���Ȧ3��-��r��>�>Nh�|g϶Tc���7�3=�Ǐww����곩�>m��Ǉ�Kw�i}��/��C���-X�������8��|Dt��.bg5D6��0�a������j �C�5*|�U�hư��@ǯC/?A1�NVו�l�۸��@�	��v@o�>���z�#�h؟;�X��<n�R4¦��\�4zE6�X`wONO�C-�T�.����+[Kn�葀���a. �?.+r;�£M��s�6?�7��?���2y�8�h�PN�����~��;���5��o=����$zvK]4<cV����܍	�����ݣ��7��؊?׏;�T�<�+O�H_���P�m�t�����G�4��y�O�hL'��}���ؤj�g���� �j�������o�0��K+E��()��\J�l�z'buv�&��%;9��P�|w�~�
�gX�kO9bc���&$Tؘ �3`G.��Y����{E�]�r����(�nUjA�EN�����l��xV�Ab�ڱ�؜ D�9��.���hgĩ>aq�,��n�h��"$fWU�i,��i�����v�����LSE�25I�IiP�9�Ѿ��cXy�~P�LW[�����U#��Y0�-o����I��M��9u�Rwq���Aqtz�S���^���~�t� �f�����o�âA��/A,��@ X������[�O�#ߋ^h���!JPY|�u��I�p��v��w=D�P�Sam0S��:��� tV���c�a����y*[�]�Wz�x�k7	��,bݺN{`O(��w{�8�CL�0��đ���'	���F���Ί���� f@��8���b�����E��ܙ6��(��I�;��� <�A��`#��ۍk�����E�P�׹����`/���cJ�YHe�,q��[�� �S�H�C/.�믺�y�ަ!]��'1�'���?����V=H��(@͕E������Kwo��XY���������X��PW�׮;$W��m��k�p�rk��L�<�n��V�J��%On[ӻ+
���9�U>��&�����\fڤ��?�r��co���-�����
\�U 8�;X�_Ƒ��a��x�W� �6�Mp�y=(N3}��@��7᪤ u��n����0��@�:>��g��i�����`�6Z���;U��`L>�Y���f��>���;;՘`��!���$dE\�!�F�
5��y��{{`|%�']��є {�v������~��q«�dz�3$Q#&|����h!�>�R3x9	�^��������-�EÇ�B��~��?��H���DTl��*��֏�z}�}�_��v�=`.�Tw�J�������f���TYK��b �Il�Y� ��D������"S!v�Y-qZjx��cA�������+y6	q�@���<��J���� ��L��o� 7��ǪC�E�;�}������Ǉ�?p]V�4Lr� F����>�%^oX�=�O�b.A��%�����*����	�>��>���TVK �	`H+���ߋ�ḿv�b�(���`���1"E�EcC��WI͌�`�k��>�$�%WS�U;7N��m1�n�����|i��UC�#��"�P�T���'�P!��+�}���\�P�ӛ��4B]�a�|
u/���~wG�Գt��n7vɍ��vV�}�j��9;���H���V���`��;\Õ�>k�E"fc�X����s�Pȳ0���S_xZ�ب�q/�m�I҃+Wl/.�Zݡ�'����I�l�����w���C|ףE�B��RL��[�h�X�B%��j|�u���I�Ll[L��5Q�M�a'՜s������~��AAsMU��<S�;�o'	k�TY-���8����G����`�Y���[��y��d�T�*ޞ����}�86�o
��oO�J�%��և���e��S�1�b��|���e@e�Wb��ȹ[_�p�����зF�hfb�G�]�13������Of�<�y��p������x����H����Gq�"��`����!�ɂɪ�d;� ����6��Jk��x��^�J�ar#h���ޞ����:�ሢ�5X q3�3̓V˅N/�W[���! 5T-���3�f��y�������Y?̪�P	d�K��_��C(��
�y�2F�i|��V�]�� ��Q�v���$7 ZhqO��a�G�Xz�h��VWp���U�dK�V	�����/�PID[��\-a�{�P�������ZK�1���>}/���H> ��{'l����8���齎�QE d�\ݍ
b:�;3�m�GE���lZ������!+�Ws�)�x���� ����Z=_��7)� غ>�ʈC�����>��:��ipUgdX�Eub�i� �l2$�%�?"���I��D7�����F}]��U��AG
�dwrU*/�Ok*���O��"0>;����%��C�Z��8_�;�VooR	�L����YK��e`���u�R�#\G�4�$�֧L(��V4T�����o1�r0K?��M��ڇ�����k_�j�\��j���6xK�+���Rxϓ���k�#i���zݎ��8D�/���D �㮂]�hG<#���vu �>���>km�6'n��օ`�3��.��� <���t�.���̂��ֶ(�
_t����n�Y�����G;D����+�����.R\ꓕ��!
C�Nn��X���;C���.C���J 1H�.�T�!�B�%��/D��#���S֎�!�5ư������G����6ͅ�G*�JuE����yV�3�lL���yتGP�7â2 k���p�_�.8���q�E�DMy�F���������I�hر7E��C !H���#������JFB= ���#tǙ�3) 6����)��+1Q�* ��룉���}.�������\0��3�DVWD#�("��g�@��Ǥl~�R����}�޾k����U~{�X�烖�Er�	�b̩?>����걌�ǌe.Ĩj���]�.rb ������`uCS��l����]���,Us����?Ę�
� ��p�	[�ĺ�����=^d�����H�v)�$��g,���bn8KvTgUE���B���T�%"��V��6-�����`�n4��`���������~ś"�V�B 1��ƢZ��~��լ�(��8�����u;�o�h��zt��;�a�B;��	c���^���]۽}��:�7�ɶ����b����������\|�������S�SϔB	]�h"sQ��V������)��U��af��14��V����zF�djup?��Ǎ��}�A�T��F��c�����o��8��ߏ�q�\+��c��8�Tlw�i���-
̠H���Hݒ����P[/��5��ky�y�k��`�`Ǉp.�F�f��Ik�笈�f� -?�:q�Q�4�	�z�������)� �5	�p�d>������Z
����oؘ"��.�s�['�:h�>�;�Hp�5u0�0�-(�tW�+I��k��V#���`@���%�����OR��Xq�H�y��,��k���m	�Gx�4V�����G��ߡ��|l�EW��a��X�3�l^k/4~^���Խ����}�P�j���"g��9U}��±��7�^�)�����z�v�x@]�|����&�9D7%�ے��.~�Ŋ�K".j��վq�Qe�zy�\1��$�J��QMITNP½�(��}����9Vw ������/�E23��r��}�)��' &xx����˖0O�0%�:]Pt�V�0�j��<�6��U7 �N�Y�vfr�v��=��w��/�׌m�Ϲ/{�1A*�%\W7�3�N}�������� 3�������s*{�m�=�~�M���ރ`��2�!����f���{����
6�:��W��Y�K�lE<jw�*��d�˥f��m�/:��s��`<C_��'4�x0��r=Q13b(FlNZu��l�e�G	��%�Yd|ݥ����T!��o�
� R�a�nea;�������}]�ܚqRu`���MNr�0oK
�A$�q�;���q�vҧW�	�k�o�?O��9����}�@��S��?��+�a��iy��2���mLF�h��:�l��d�̭�]�Tzn,V]�o���.&� �1N�?h�J@���R�O腗7�]����'�-���0Ԧ��mˋ3Fkao�PYT$$OH��g�u	�Q��z��t���<��=��<zp���Ax����",��V~,$1Y���䖡4�܍#8���/:�ɬPɀXÌ5�S�{g��;J�k�P~8ɻ�i�}�7���+�tk�#,�o{l������f�µPa@tW�V�=Z��������>O(ގ;nę0@b�*��J��J!0�����U_l�d�Q�ЇE���F�<.T��l�O$
�-�>�0	�,�S�: �x��|ϙ�K,�p�y⏢� �[	�25���3�w����Ў\��:�A$K`���ӭ��ĪC (vP߮۶.U��T��]��ZCʩ�5�(3�Y�Ҷ1�|���o��փ|X�W�zQ��	b�N���m�3��%���Ok��vY\ų�	�hz.���"�* 
�`L��i����ܛ&�#�Y�*$��!�B<+.��{18���@��+��0�l�@�T�Q��V����E<X��ַ�A����T��%�qh���4�Ԡ� �I�|-��"4�+IC�!'R~��1P9A֏}.�F��<�D�ѼP}��ΰX�����Ņ��x*\:�E��.�7퓾ǘPi,38�� d`���� ՚�Gu`gx�\�0{1^�ġ���5Z|�Ƿ�b��;��}łG�!�E)q���Q��m�^#)2F��A��D)汪���D�����i)����6�p�q�٠�t?�B֬�	���5;��5����J�-���h~�,����aA�8�R��X�� �� �{יZ$��rġ��G'j��8d�$��N�-X	Vt{ �'O��4`.
I9�t��`5�'�08�|)C�@�#���Y�5�8>&f�j��M���{dt�v{=���᫕�� �"G�q�ya�sKn�`����й� [��]H�j�U��>V���O�,{�-�?�Z����2'�"���y�}d**3zAE�-�8"��ٺJ�L+�z߷����j����I�����?��s�S��ęB�ZEk�5�����K�����"	�����$ʹ�AG�`b��vN; ې$�� T��>�u���n��GA��cwn~�#6�@�6�����c�fL�$}J�ݧ1H�%��?#��3�h��Ǧ�.ś2��}�4b+��	��L>b	ΰ�w% "�+~�nY=��xc��Bg�5������}A�F?pm�z$�H�*�V; ��7���X<�`�c�:��̀��8h�|Z]Gݞۂ��z?��>M]cio1����7� ޑ�`h����z���������	������Wz;�%�ϵ7M4AD"՝J��gⲅA31�`
�s!���*��h�I]?�s%��n�����	1&`6��������OAU�� '����>l�4���7��F�;�b6C�$�/��XUa5
��nA.؄U�M��M��{u��}i w�p�*�W�Mf�����x,�NF[�j��/H�J��blr���c�W�r�lA^`H,I��;����g�`@�6�=x8��%�����?hއ�ю��[�A~���ނ�g8�+��<6��1�}��ڽR�zWZ@v|�/Hϋ�����h�����@�{w�z�ɫ�"�b��}nZ4R\40�X�[��� ��Ĺal��t�o@�"���|�(��￙��w*���n�(O.���&d��E۾:0g�K-������o ����ʶj�g��	�W` ��{�VP/�)����k�@'��6��͠��ݵ�2�.ݰ�sF���ĤЗi,I�����^��	�]��D���\�����0CB�5�>t������������w�����P[jQ�~t��U����HX9���5��O�U��ܫj!R�m���_���Y�A�}�#$�_{vz��o�铵h���[�s'b�3s�@�+�r H����F�x��a4_�f&R_� �$��eI]�N����gu���Q �;�[t�ys�Q����m��UX� cj �bn7�l�N`�\i�;�	�?k��	AY�a�'Fu6��$���U�,�{t��7Z�3��C�z�Σ����MG�E�W���!uIwG�%�=���3�&��8����,� � Q;������_�%ʚa�D!%�+�����K�#��y��;R%��Jǘ,i�p�P��c3۩����4���:ܚ�t�&�Y*�Y�D�����_U�).^AI�IƤ ,6�t��4p�m���s2�7�!�z����:�%��^צ�׈�łI�B�j�����A��O���Ҋ,9/Tp�P���۠$0�B�� MN�9�=�P�� �x��E��_ �D��~��]����u`o��4- 6QK��
�o*l�;��@oOuPJ~�AH��\δ%@��T0��^.�W�?�[�k�]p*��8�磇d�I�)[�gv�ʅ{�/i69�8(����53X��%�f����G�ʂ�>"|)=ű�w�+�6�ۅ�_�Eu�Q��]^HU��+T�0p"���&U�y���ǡ�q=��-P9h, S�X9ҹN�X��hQb_v�	�'���8�ؿ�����+B$*���7���@}#���>�uq@ų���%�]ז]2oO�e�b�P�]H��@��
���e��l�bS~�h�V�D_��$�������6�zl[�]�#��#�S�1��ƛ��{��Y�П�T�?�},��$	��D���3Jބ���� H��9!Pe)a�S_c����U�� ?�%9�������L��z̃��"qR�7�� ����ų~��[k�;�7�$L�5�_�>�ˡ΃T���ثN�~��܎�]J�˂8��v�� H��?��}�-o���	P��3�ˑe�
H�+���b`�D���UN#�EC��!H�u7�i��CeH�S(Sv�Ie_{��.��DT8ދ����a�V���5���j�ij^���t�K�P*�Yy�Zf#�P�U+_��^�J������Q~1&��G�+"��q�9Viq0MD����"�)1X�(�_�w��R_M�U�p����G1eh)���EP�(߮�X)�� ����k����"X��w{69�қ���� TI�Z�����LBWh�#��[	�W|[a_I��"�r\-�m\6����s�c�⣘�$3D��ϓ��l�e&Џ��bt��:�J�I`�b� �$Rs�� �]:Ԡ���h'n3Jc�c��T>a-� �j���?���X�.��J���QH��*����)��2/e�.z�zҧ;SĽ�v*Y�,�hHW*�)aH���4�a��#e�Un3�K���H<��l\��7�X��RWou<�5�&=�ʯ�8:Xㅶ��蓣�v�¢�c���د��:�/ ���_.�����^[�.���H�����)��E@]T��8���U�/VP����-�H����{nT�E��#����X��87'V]R�@�\5Q��EӋ���.-BVMu�q��t�"Ĝ�xi�>
|�K����/�^� J�|�J�?�K�\��:b������m�V�^�0X��]��O9���Z��������[  C	c�=�Y���Xd�G���D�:���`�m�i�)���/ޏ>N�=[�Ꮛv�;��%-~ǒ�KS~��A�ϗ#� 5Z�t6�ăl�/�06M^��O�C]ݛ�Q$�|8.�ǭ%��p���~��߿}����x ۶翉�o���?4pt�k�8��M��s�h�]f�E�Eu]��/�5�����)O��k��c/?�������j�҂�T>"��>{a�|�:0�!��|oL�>X������a��7��5�耶�i�#��POtvO��� Ф{+�A�=�(�t���ڣn���m���#�k�\�8��ڮ$�NB+�H+��E���mQ���ΔR�J�;��w����}�N��k\�(��f������%vi��Tw�|g�Xf 5*�@��� ŉ�K�qn�Sn���D�m!�9��	p��Ѥ�零�@CU���i}���)��Z�e	&�
}���Smt��}RP��\�f�G��o�Ӣ:����������-��������K������aˢHi�j�D%��o����h;=�crK���¹��w�bʢ��Zg������k��nVk�^��:�`h�/EWu��^Q���gU%]���I�+~���&'�H/��	��@Ww@���V�O
)�b=F�S��=HЗ��l �-�2B׌^��b�ZeuF�$���`l/���3�+x��i�X��&jEY�bۚ�3:�Nxa�}K���A�2�;��b����y�J���ZZ�!<���g�*ķk�'���.��W�<n�V���x4×���F[l��p ��t�GڱU���}��{�]��o?�������-`��q�����v²���_I�s��+�� ��+#�c�6�~o~o��Z�~��3��R;�u���oyk����~���wN���D;�mK-gLg���|���uu�9��²'n�eS��+�)�uJ-b�y����F�A7�k�?�U@&B�zা�O$��#�Rl�.`:�F�?��R�n��W�� A�*�b,9(���l�[rc|�4����,z����Hb�h,�z�E\+�b2�S�s�X��mYT��ߦ~�0��
�<�Yz3bd�_8 ݩ:P_g?-ݕ	Ǚ��;���n_�������۷��Y�{8Ϳtv|�f�&�z_��{W��~zE}�.
'ł�=��寉
}�p���6��e��R=��ǇdP�7�H��	WJ�8�.����3�%"�KLxl�[��-B��u��d���b 
�()��m��E����0��/p��8A��v��).GL������d�E�����n@�NU �!��U:`[�.��X�q��y�O�~/4v��?�o�r�;�R�[?�,�Qɤ�E�Ƀ�|b�q��s4$��V DǢ9l�����i�mE���������?�*����� W���<�) B�-�����m�<���.m��B��]<F��ȃ�3�nI��W��*09�1����ZW����5&��70$��{�'0�:�2_���mP������wka! ��y�R�Ws��?��#@�i�)�>zsLTepY����c���P)����DF�+w� �H��B�������x�Lԧ/�o�L�M�u[��u����%ܕ�~$��b]}k�o�F�.��q��޽>���ɵ��/i7��xU,^_�UcwԼU�I�_�r�3�MY� ��.䤺E��6����R"~�����31�mzV��\Yg� �,����0��7�,Vg��E%0M�0|�Lv Tχ�1On����B�3�c�S�|��~x�3\m�f�����?�1�eX���Y�ci�ɠ�мP�πu�s����f�b�D��1b���Y�Q�F�rP����(?m߄���-X�o.ry���bb�8� ���TØ��� u�x� W�~���/�P�ԃ��Uw�!��t�b�8���`��]�C��H4m�+@l��t%B}�L�'�[[a����Vl�Q�gF"08�9e���6��/&�����;Y�oMi���G�8*S�ig�:��d����`��%K�Mi>{	bjy=q�ŇA} �Gq����d �1��Ԕߔ�G~5VJ߃�IM���	��;�S��>=br�&m��*�D_�۰ÑG���9W;�OF�9�,�_P���:�=���ʋM�Â�VG���-�E��R�Ɇ|�c�{��yW��~!=�[/�;V���x������#���Џʅ?��wt��J��z�э3����'��/���l�u��u%�=$1����������,j��$XӹV���}�Tk�_䏒�t�q�l�.���d��Œ�����g�_�Om�{��F.(�"Hw�2��C��HS�	-��� W�1 ��ʈ�/����C�Db�Ī� cL�#s�؉�%5�I* �?�u��/�d9�v4�L,Ę(�#��Kw�  �3��w��f���S�*{�	uU7&j̹PE�n�j^9��S1�P�i�gg�ߪ��#�P'���r`�Yj��n��۬%]��d\�ga.T�=#j^p�9=��}u�b�iL-�w�)�MU�-������Q3<w�Zb�B����"�]]~�0�FI��{��$��b'y�~�r��C=���@�,2b`X�1�R�6%��P]�6�<�apls��.iE�j���mn�����Ǿ���<Q��ҐUf���rK ��59C�q,N&'�]�%�]<�)�M6��@��3������0#�����(j��TV>3
Z�p�]�`9�!_�X��NO5D�*��I�,��H�Jeem+/!х����h�
܍(�����N�p%��ׯ�䤻���z���!^��&�@�*�AZE�҇II��Vol�m�μ�G�bu��v��MD=�^���ֱ�l�Lrη%��h�c�F���ӱ��An����z��~��8�f>��d�0&�6UI3���"�]�nKeLj��3m媥��M�'dv�����2bu���M������-�jӈ�ZH,���O����V��C���J�����~ʰt�\���wL5�n6���h�2����ܦ�����?x��"{��q�l[��oM����c9�L�K��R�~��q]�*
E<�.C�fe`R�;g^��>HaͿ?-���=R	mVF���tcƨ0��W����z�޸L:AM^�����8l��m[�:f���2��Է�����?.�5�+Z���#`<1�З��~�4Z��j�L���T�N}(y��3�<�+y tݩ�~Js]J�Sy��+�s*ړ�+>Wd@Ex0X�\�SU�o�����C�U�P4��Y��E]5�"��^ީD�Ds6k^���n��*��������I\B��l:�<c���d:A%X�O%ʧ����������y��5ʤ������:i�k	��a9A�ExQ��M���&ou�TmT2,�� u�NE�A��W�F�.n0�q�q���ږ���}���BE;���Ib(�b8�d�*cTf��A����ju VЯw��{���@b��mG�r�3�2-�N�� Zt_�3����l��8������'�
+l�����ʸ����|�#q�0f�j�ʀ`�>�I���������lt���5��|FK�,1�3�#M����GW?�c�u�(!�b�q��\�O��7�. �|��`m�(-��m2uu��&֒��d�ݦ]��x�[�r���!�d� 5���+H(����!G�o�������=z܁掫��=�J��S;�3.���� �k �D�v�@�M�Ѣ���\?Tɦ�n�P��y�(�hNH��EP�\ޭ�Z%��ս��|nN�y�;��]+3�F�������y<��կN>m�lHe���^�[�w��f�5���2�_�^�O�m~�ɽ?���w� =0��e� ��F�"�=���ޒ���?�"��=.5��3����"3LG6�°�\֪��sI��%	���B�}c���Ķ	H�@b�j�'a㙃&���g�@�į�RU�ʋ��c�Zz�c?\�w)�&�9m���,�QJRxO`D����bEj��1��~7�X���59X�WD�������um�˃ߴ^�獍?�/�(A�\��e�����4Q��b�������:�">Wù�o��Z�$K?���R���T@U1J;�96c���%v��8���<!@X�N�*���
��j��X����d�@"�����, u}��6)�)FÛx{ܒ�Z�?ӿj�j�R���ሹ����b0}�&e�B|�<�9l���m�zY*�J�`+U���I��) c�V�`wp% 
��qa+�,!�b��A!.B�:I(W�w;[⤚�x�����J�5�	���O���f}<�,��� ���_;��H��������0�	B��l�̬��PUԍ����" �Lz����*��F'}�<�H����	F�`�Xj.Hܚ�M�U��LavR������DD�F���KQ��J?aT��_h_��ק�y�ݣ�;�<Q�<�$�G�G�����\�]5ɏ�ކ�Bw�d�D�����J^�Jz��/�N]�$�K��i�.)ew2���O��f]���zQ�Ѵ�%��Z������nk\�7�R=�tw��P���$=�F&�'���E��~���!	��d(K�yn%'Iv�d��5>�DV�y�_��������WzSTqDW�*�d���s��8&:V7^���aq<=3P�uE%�LX�q���ș�f�|?�6��nL�n5C��?�\{�s���cy ��0i�C8!x�_/D�H������d�D�����G�0�`�"��8���	���q���:��.�L�)>Y�J�#�B��9��}9�;.�<aL�׏�GP�N���U�J����\$?�}�-����/%�#�r���F�¯!!�My(�a���Na׌��bދ��>3w�	��/���C��R9LJ���}B�G�rx�f���D�i*.�0��k��W"E�Lڞٓ�j]���� �xz����+���l&J%0��A[�{Ĺ�
�^�o<1TV�er��P~�$U��Y���i��YD��F��x{�}z?�<�����*.̾À�s�H�$wmGo�9�PU@u�Ҋ�QA���$��g���֕TN��l���ܓD\JùP��(@��#�g�3��ecI�W���h���Hٵ&D;�]���1v�D�&�T�d�s[hU=�r�����r\]�6N�:9������SPn���3}%݃D�ӡGzɃ�|�/�yT�e�<N!m!%��EL���jX�Š�6���<,�v?3.���S��	���Wz��䭧��ӺY�
~��{��G��5�:�Z��bu�o�Z&�:�H��������H��~���@r /��eEk�0/H���T7�s�6�b�4W�|%="��l6�O��I&z���ޙ��+�ߴ�N3�Oyo���-�����%HN�x8��a!�3�S>A,��zتm�3��u����8-�b%-q�@ ��x؂-�%�eT�>��B"���_Ԓ^�l�Z�骂U
��=&�����΄����󩟘z|��y��P+LAd��n�c%=�����0���g��W�������mK3�T�7���M�=����B;neh�MNCK�e��__�����b�5����6u�qe��t����`��j���@n3>��[�~\�������w��խ�f�iQ��|������`�*%�4b�^f�Y쫓�-9=U�`'�;�8J����I5U���_�Y��7�����Ens�t��K9�� ��6��w�'m����L+;�&���K�ܣ�W?����P��mX�:��է����q<�90�LF�Z�1)��%���smw����Rb���s�;�BP7����T'70��-��i��c���`Љ_��*��� ��_��MJ��1>�X��ۅKW)�p F��@8�@Z�%��V�7�ޗ'7fW��U�U�/ u����NC%�:k�g���J�Y�%uLYG]��ab��/�]qp��� (%2��O�P~WĻ.�B�����*�����Zۏo�R���w��$�\+&Tb,���W&1��>�]-{m�d+ 2<���5��s��N/�۪�p��JƁe�Ku��*L�	e��g��b�U��j��A�6�@���H�'��;�O�&�+�i^=�7�nRF��ܰY��z���mK�g���9�z*#����+�S��]�]uW�<{�W��\٬^�w�n��P�R��T��<qJ�2�yy��B!�ƦP,�� �y�����kl��׆?_�bF+UK,�q\n0����C�u㳩��zF����t��|s� �o�{�R_ ��Tc@x `�}(�_L?��;�(e���2���d�=ꊣ��;(AW�����84��+��_�/c� �.��$�L��*��D�v�t-q����v$���E�U�j���	��&+�@�a� �;�He��A��?s��E���if4�~} ��f[���$4�C��I�z3>-�2ރT�Zbw�$�2wtp�`����W�~Q5�*���:���J�:��ŴםWp�yv�	:T�d��`�
�'�Q8�D�.	<]0�a�� (�C>)�ŵ~[�g��#nK��g�_	\�p(��ԩ�����/`wx~�4�H:���]O{�Ӳ�<�u)��8a���L"3�ug]��r�`����-���o繸D��Bd�G���K܋���u�i���'�fAz�`�\����_�x_h�$���۲�(m���
_���7��U;��d� Z+}Q��A�~a�߄j>�\�s�=�B
)G�l%��I�e*�(-�Ew�r�l����f�:#o���g-�tNP	��j2�����������
������W�Oa���e�5���AwC�yRv�T�[�ѥ�a[����-�H��&Hu(S�{-'��谵���_�U��5���$����t�^���WJ��rw[��e�.���n�a�<�^N ������B.��ns�9c�Fu�6W��JRFT�Ol>�|(�8;�O(kh�}�Ɓ�?+�P��f���#������Wb��M,��]�"ex��������*ݒ�S�>D�a6�(���4{�H�Y����Ϛn���}ˋ�P�+���ϐ������Y�g,ʩ; IJL��{���X�]�s3����a�*�n����WD���p�M���vT����R@�O�L���c�O�ߚ���L�f��o�xe���� P>�	�k��a޻���B��\/�_���K2���4���թ~���pe՘�� JN�0��_T<^��L��8��y�Y�2'.|���UZ�jZ`�� �E��4@�w^Mo"��h +���c��G���u�0���N�qE����Zc ��e;�N�`
���3���t{��-6�|h2��]��� 0�5�=���h���;�1�U�|/�i��5l"wԣ�H-�!΀��W��jӿ���(���&��IN�j� i�7����W$Ҁ�|��Y����V�X�F������[o���\��p:��j�ù�V��ӘK�����	�����!WP�a��Ӆ��+���*��,�>V������������9C�23�$��󀾲͛�L_ڞ�ů��N}^6�����AZ ���ywc�2��n9�|�E�=n�z���,����י����������Y>Z�f\����[���%@�E���4���l������;TP�RO��h��u���i�� )���k%:,O� ξ�cQ�	U�_�~�po=���X�vq��{�ޓ�v�{��k)�i�~Fԭ<�Kͷ<��~�dZA	�Qe���zl����v�̘�_��� 'X���E7���#��)̌4����:�� H+�f��^��bt�J����h�\7c4���e=���IS��U0�Tzma�Z��.�mAX���XP�°i;��t�O��?�m
�pN݉:�2�%^9��;b �����כ�in���?��v�����o���&��T����� �Ou* Q���� ���4\ԢR50g)���y7�\�<����C�6f�� ��$������RU�)������Bp��b����5����L�L��A���6�ی�_"m�K��V�#�?!0=���k�n;����l��[�/e��əbfxPz!��4b��٘��
l$�Q���]�2��%�j������R�=��I�z~2c�p�{�ٕ���c�e������מ�����Z`�i.�n�Pg��H�\�>0��������ｶ�1�Cv7<��T�������rõ��Qu�B��sA���6U��ߌ�f�3���>p>��?i�|&��)����Yf�vP	����t�*-p� P1WD~1P�DTK)�wRYh)�b��="�J�6!��s��S^v���X�|��Яtw��-��X5w)����T��5�J<>-���<�IZH�a�Z���e�Qw�ǁ�V������i;���<���p�@mH��7��p�쯅�=��JH4�/����I�0oJ�C�P�q�&��x}�!\.�9QԾ���Ay��:n���h���Ö����C�_O�	b�H��n���{��;�L�%�WJ���{6������2��mꓭXc��*sc�� �b��=�@�H�o��O�o�j�W������o� n���t� >��T�d�<L�u�o;��J���PMi�W��Aq�V�A�h��V"w�r�_�Ÿ��+v�����*ӠD�<Ǚx��Y��;ѯ��4���S�n?�����_(�~.,��w|u��y	�UIa��8���)����m�n��<��79�.��씁��r#�(��xWu�N����]]A�M�����E�����ݕ���e�تG^�����(���J�O:�|������@`b�"1�Veo&�=%;}�˲�{�0����0Vjz�kr�듞��^̀�c��_���m;H�?�.K1`X5K�1�i�%��W7A�J�IצI���� �����R#��;�XT��4�[�ti��7���;/LE��D�:`�l���Le�{� Ư?3Ų�k���iA2��Wl��jBe�\�.����o�t��a0k̢{�n��6]ڽ�� ���"���o��լ��-��ڮ��_72ݟ��O�-��i'z�"9 �y\�EUP{�c�n7u�:�xS�gt���ߑ��n?)�Z�_K�ߦ�k��cE�l���H~��O?d ����`e�.g�g��~����J~� k�][�B mj�jL�wTQ���_����ޓ�}��}�r�Q�+�L�*%B�Sfz4,�>�F�V,������ߙ����%���r�1ޫvu��CA�꾒�����"�#:���	�oqTb�9ջ��9���|������7v�~~d��zO�^>�C�X�K��X�b�Yh(MN�`���>R%Xg�w3�83�
�:�����q���uw�?���X�v~���a>I?k�'!�s����9ѓ�]tKηo�D>�����4����|�s�� mn���HZ�m}�؉�Pշ��m�TlV�I�L̸�������P�*B��t1������L�O��3��q>V��9���-11І��O�ه,Yl"��5 � <aT��ڵ��i�<x��w0��2SH�t}Mq��8����{3�=w\kA;�W��,ӾX���B�٨/�zW�q]��/7x�8&usq��m�",�Rf&Bx�z� ��h�c�xP~��
{ɢ1�/_}��!��|��������`�n�`.%�у���Kc�ti����-�����@�l��~�g:~���{?���D��%2 +%`)�w��O��k?SAf����Iw�q����5@5e\zn.�VS0�a��,	<�������0��p�>c](��*�r�<E����`g�$�８�҂�!c��s��B��z�2�R�+ ��%�0 ]��ĸ�Y�ǀ95 ��-��뷈*؁�Ѽ�:�������?_�j�>�Y�P�y�r�
��AK���)=P;��Q_N���I{o�RmKY�����C�l= ���$�_��_� &Z�ep/�Ҍ���{Yk�� �-��8D��ec���I�{ߕ͏��G�J�Tę-T� z2, ��n�C�O
\2�yQ�w~���-�+�	k��� �����B]�S�k���a��Z �-�զ�{m����Ѐ��v��� �<E�
�]ʺ`��K'�u�?�(�&�+E+���(��.��A�ݝ�t<���.�B���d(�5���V�\]�(����xt���^����x整qs�.;,��>�BZ�'1��K�_��NF�)�ﵝ��<��y*�2�.ͻ��3B>+UjØ6�k�5�!>KMR���`o���H�0���)���4��w-�x�A���������P��8r�����ϋ�_E�m�ڭt߿�va�<=�h�G�8��%��V|��#oD� �9S���H�@���(l|�%��?c����<� �����U�zz�}���ճ@��J�fYT�%��]�"e���f�=��3���#P������>MZ$�L��͒�U#ܮ��p�ss�IE!������4�j���3��y3ϵ\�2���S����M��׿6�^�.@��������� �)���<.\�wF�y�=���Rr���'������芒����5�T)x���Ź���ٞ۠j�h
�kU�Ϧ	˪�b>To�-�-1��0@�IWRV3��\�{'	��ٳ���7'g�$����ג�ۏS�.-�`�j�j�<�H�
��89���
�G)�5��,�����~�nUX� � l;J$w�K����27TJ�`pxֵ�5&�+~׻N��k���$r1��7��W��E���5\5#�T��iܷy���.i$�������l_�ԋ"��Km�>�4G�qnHh��R��\�1T��i���)��zT���@�l�py��V����)ȋ��x�a������	����P�"K���G�R� ϭ��y��f��|M:\��${L3T�������zz`í%3T��c+�Q��b��=��]�5M曪����� W���?h})�T ��5�70��,���{Zֻ���z���n<�t�hb}��Ԅ#�ȏ���f�i@��WUݳ��z�8�N�Ut�gJ�������������t�S��l�H����
�XIw9�<b�������0��)�����:���[D\t� Tb�aҼV7*�>KW�J�'�o�c`�&?�{��-���y��#��9����y��=~�N�&���Y�\r�EvxV��2��e�5Vۛv`_I�StL�-�,�*�m��� w�ߖ����p�d����ǩ>V۳�5�5�\��J��`�#��r׺�:d)	(zI�l���n䕞��YmY<��s��ސ�]�g>��y�^�zפy��ή簎�t�Z���{LyOEIy������M>;)�,�Y�)�L��N�� ���T����fv
v�V��b~)Tr� ��O3��n{$=����>ر�ͱ�����ゴG׍�C���9zQ������+�@S���"J�wi�b;;j�����Ca��s'�љ0W�=������lT8ÿ5i�o����E���^��˦{��f ��~D�"/sI�E�y���k
�r�'�]-��P���
�Xx�Uc�~�j]��aWw��9钦i�m�|!=P�o�N��y��荰:(���� � V���Yƛ��S�a_�n+"����6�� �]�pp-��?��,~ �Ɋ�:�[Ym�@#���2����]\[�|��� U����~�����0�>жj�B���P�P+T�y�o+�����]���� �i`���}��1��I������j��k+����}{�X�W@�����I�D	�ŷ��-Ƴـ�>v9eqܹ�x��p�\��y�Ϸ�!z8��]M���|-Q��+:�j�C1���u>a��s���-kj�4�����+-T�� �H#��N��T��U찜�+��Ws<�k���-۬��㢝��R�m�f%ͣ.�]�8�n�\�_lϼ�X��k�ˆ��}^|���oL��{��\V�?�zO�jYI]'�V�����woJy�ؐRE�y�N�i�H�?�)�}$՛�
�}��WXvJw�g~pK�N[	�ҪB��ub�� %"J2uv Ԏh�������clq���x<����ӇmY]�.I$C�5��}h���q�$r��zGߔP�'����0�ۨ����M?ס�`��*��ü5A<�/����Hq`�դ�/2 �����Ƕ��60��E�����j��`�A����#��
�W-d��՘.0��Y�TǼ둈RA,���M�&����C������|��<o�'�iKO0��-bn9Ww�x�5�X�"�}ͫ�6�ڀ	/�(U~ݖ��2�;�m�~Z��C��c��;��oE�{.����ݴ,����R?3�NcpoƷ��M�bH�#�(��1�=��8Oη�S6�H���c1r�M�ύ�76���%vS��QH�i55 �l+�4g�gy�+nM��C�IZM��;�V�;k�T��z�ch��:������Ü�����ߏ��N��Of8ٔ�ʼ���*���m��w+��w�j��
T�-��5ס3��i�{��Pi��Q'Lt7�q�xvz�](��f�k��Z6�cf �Q����<��h��[O�Eo��y=]�_,T��(���_UU�Ƙ��vf������~jpӃ� Ug��e�E�jƟ<��e|����u2�����-t�nc�M^�1	�C�&d�� s�(.>����j��'����u[��+���@�5�"-��7?O�1�{nz��JWPiw���z[g��O���0��n���8�B2�ew��gu5��BIMu�F��V�F�j4Wq��f$XQ�W����W�s��5z��HB��j� �J����Y4*�u��f]��� 6��J��P�����ߏ���:��u�:�M�"�3Ԧԯ��������z��Cw"�s�����+,�y�7����R��Q�:����	�$`�Xf:�� ��\��xJ5�T�9�m*���AHE്2�u��!�Hz�d�ߜ�I~N ����v�5V�I=&+:o2�]�:fOF�z$9��d��N��a�z�j,Be���=�>���#�F�fn�
���1�՘g�U��n�y������gX�l?Խ�BDR�vǳ74jK���&7�W6������_I^+�`��BC/ k~�)"
Xl��Ŏ=r�)?
:H�pF�m����O������g��c��Q_�SB��u���:�?{�T�R�k�1�w��(��S0�=�"���6�Ľ��g�A���-HJ����qW�Rڧ�~�=i���T��u3o���T�^ ��KNT�2E�1�+H���{��i��a��M۶�A��@e��>~W�S=�F��k����{�9G����[!=M0T�(��-)'4��`�kl;SW�2BV�4�I�I�}m���N@��~�]���,=&=֘�3^���� �-��{��#ž�!>ˈ5�2^�|b�]p>]�ǎ�T��I�mA��1��t�B�@��{] *����@�Q�LNR���8h�,��M%�ց)]�z����9"��DXiJtr�sS>-���:���Sa����Wl�)vK����~�5s�["�:����j�~C�Y���i��J��*ƪϿ�T��2#_���~�_^���[E^�C�LWE�y��}�oO�+����2D�B�Ű�?L@u|H�`�t��1���8.�%�	ѿĘc��n�>>ǆz��6�K~ƀ}C�V?M����0�_j��+N�@?�[\]���,,�֨1�'��H�JV�_��Qj���D�gQ��V�y��x���-(L��$�+�宺�i�N6���������O50`7�x����TI#�ɒ��P!����_u�Th�t�[��yC�c�6%��zX�����!~���`���OM�s�"F��r���������0v�������A����LW�-�|\�z�=����fb��W�(>=���BI��ef�i��E�"�ܞ��WB�M]�I�=��Qb`p�^��w��)s�*�9DpNn�Jnp�}�C5��Ŷ���Wm�%�� �X�P��� n�R�</8��Ѱ�T���J�b��b��V�w��Ѩ��4��ɶg�a�*�l�0��S(���u���DG���B�ҫ��b��`�4�>�[�����i�(��ٳ���.�x��W�[�~�O�z����G���usC�j�u�m�t��^*`_u�CZ��ϯ�4�Wȝ
��$w��f�t�G|���{����+S�b����yLu��bزj��q�87葦էu%���߫M���e@��vA�O݁��ձ#Ot�hA�����~<��W�w@���~�<e�%&��F"L��w�c(9����K���� oE?���u�*v\�������V��*D�Q�U�9��.i�<���Jm|m9-mC�Yҁ������&�����G?�CL+6�1[�&Zl�*��a�=@�����m��'~��-��������ȑ�Yf�.�~��؄���e��V�15`:W��m�����]̷���PC��,Ă!n��u-6�C��\`�����8"��o�=�[ۛ���t�`˩?��!�éS���-�RY����7����r��ۡ����q��َ�?��!��+ғj�������+��hx�X ؑH���9�*[_tJ��ōW9���k��`HJ�;�f��p�p-i����o-��v�"U
��#��(φ��h-R��{�b�G�p��Q�t�T�z�ZɌ�ו�ꈚ����es��R�k���%�B��G�]w ��UʃV��GL�q�S� ��m��Z�d���Q�D�du�o^	�D��3�,�����k�\D1�:�)F��4�0|E<ʛ�ԇ��KI�)K=��5"ʅ8�D}���+�F���ϰ�GW���tZ16��_y��:�p�ȷ�t��l	��6\>�A���N�7M�}��߇�I��kB<��Sw�6&�a��Yx��N��b��X�(�I}�ni�7����^�e�o3��. 7<Y�sy�`V{B*����ӡ@�$�y����'9��:��,m]M�o����yĞ�
��2�=��*�~���~��� �880:9,��>���@50��P�:�ql^����~~߭����!�d{)�K�u�p�i?9AH�\yj�/�\�AQLr�U*��1xO<�L�e��BcҾw���t�����bQ��<4�S�y5^� 	�@�q�K��������}-9����t]x ��L:O̽����Xa��_B���E\w�X���;-�V�ė�?�'`:���e��_SڸƳ��d1��9q��`���;�6�L��0�.��+vk����;U�.�p������?ޟ3��ՈM*	HG#^ʽ�ͦ�� 5e�Ӷ��F��$m��CFx��1��l��7�'��҄�����b?p,�U���~��$N��wZ#��_o�-v13pO�D7 ��&�Ӈ��^ӱ��T�~�|?�սb�:�Ѻ+�Ua��g�������q���;*�L�7���Ȱx��# 7*��J�s���w4���Wѩ��$���)�l"g�D�@���S`������Z��0H,�����)�����5��DC���/"E�:J�<'�y���ߨ�2ߑ�q��
`'�EF�2P�4�]��>�f��w��{_K�=�E�m(>ѓJ���$�`0ݶ�=e�/�^^�Ʌq��?P���49g�jW�H��$Ų����c��u�p�%�5J� a����m�y��e�K�͔��]"���-�eZ���h��;�K	O���jw�w+�b��Y?2\i�)ѬX�F�~�L
M�IQe;���;�s�1����4i�`	?�`���[�90*����EwB��+9܃6���"p��W�cC�G�q�Gw��Z���ƻIh�Usb�2�>��fH��N���A N`��AJn�2�:�,W���2<'��6kL���m,Z,׭?�S�HJ�ס�^4t�aXҟcU%b�bV �f���D
]��x�t?Vס��a!�ME�h�'�3���(<Y�Oj��dR��q4DmSy�k�����$d�-�V$Ll��#S�};� ���]��M���T=Y4~�5B��C�z� W����m)��?�����ޯ Z\�0g��K[�7�{�:TL����p��\1������F��84L����Kb�Ҕ�i���ş��X(�v��+����&�?�,*�%��D
x�0��B�mwCzd�H"�4�*[ro�)�Wnd�ۦ���\B�yf�yc��8{�����y߯���'��;ݜ�P�Jk���u�uWF�)����r)?�<C���祧���n ��_�QX�s$V�l���������
�yI�ޏ��L˟��̆����瞘3��a ���V��S{,Ϩn`��t��J����g��$��������:���㩋/�a��i���y�[�Dqq�� uH����s�J��s��i>v��-$52��M_��I��yG���(�l��Vʶn±ߝ����2kL��ȟj�N�[����E�UگV�"Z��="�Ĥ���>��D��<g�٣�gk� 0R�������2�|4���7�_ w��Bw�_�&�~�b󸩸�����D�<㥩�������g��gG�[�B�u��I�=.�Ӫ)��g�	 E�S���j��V՟�6T>2!�q��#~�F�WD��Ţ���W�2w�O����b�-���*a�	�~�_Ďvu� V4���%��1���Eq=��Y�D[L��ۈ��O����G�ia��h��s[1�ȑ�O�T�r���D&��y\�� �#K�ERd�w��*��o��i�g[���=�V�X�_c���qTO@Jm�Ĉ�[���j��c\�Ѹ�J]$�ޞ�%dQ�]��JOT�T��Wrq+�v�^�+�-�+��vpN�OE�U�5y;\
�vt�R0l���Y� �=�廞N���U�@�-��
��X(�c��@�/dE &�D=�0�;�pmb��8'��XZ�^N�1C�`]Y��>i�f0��Ey���^�/l�N`�B�3(��)W*����``i��s =�§I7��;��n� W2���Ρ���gd�f��D?X�b��q��FZ:\@����e��7����� ��f�����P3�,�����|S��&����C����ЯYu��|����ov����ʢ%_,0v�d�����z�H	�*�ZyE��X]uV;Y��3h�y�+�����=�w}
6gZ+� 1˿�N=pI�Z��f�)���'_Q[��g�k��Wי�Wi�1`d9ZIw{�������$0Ԁ86@ecQ��>7�k]h���lqo�o�}����	G=.i;�i�.�yNP��G�ո�ڰ!�mA_ęo�P�~0��T�;��N�j �� T�h��b{����������+���`-
�`Kt�J@� ,��iT���C�A�ҷ��X�N;���)B�!���B2��X �e|�X������X�#���9h���U����1�Ĵ�L�%Pt��@.�ޮ���_+�T�*�9`�}���%B��I\#M �4[�+pVU�D��_'(�[H����>�i�=l���M2�p�I/���*�[HI�J���Cg�gc[`��#jH�j�*��$x�E������2�n�"Um�B��z����&�AU��6Pm�1�{��#�L�l/�F'ߐv=�p�X������<��y��=�y���j��I�2�g��;�jp��*K��W�.zC:;�9��L$?O��]�g>���6$���~wݪÀlR
�ZL��8YȘDY�ߛ�/Lύ656�S~,Q�W��,���
�����Ӈ�n [hf�����Dލ�Lky�O!*�X��a�N�`kbι�^�g~�F�C��Z0R?��F�7z��N��o͓i�����'~�4R�W=�G�*��g�h>V. ��?�A��Nw�o�����j�l/�	c�i��C�&�H��%/ eӕ6}m�ٖ��E%�eC��n��O33b��Ql�k��%���T �`��V�3+e*Vd�t�g�Ok�8��@`�����UѠBWs*�Z�s�����} IqFz� ���^�`��q��~�#�nyT5�&�N<�����C*�;n��c���~��+��)?��EFiW��yp�]
l���>�������{��z��|zy�d<k��ߣ'}�\��8]�;#׭�����>;&�ׯN�a��xc�={�ua*�������k�������K�A�Ӭ��Ӷ�C+t9���κ5�P���50������Ũ���ϖ��r��]�)���\����(��?(��K�x��o���Uf��;O߄�{��%�n�%Y�Y'Z��\��@E��"JK©��ϝk����_�2�1�rW��0ΑIp�Q^����5�-2�ᒃ����}T4����1���Q*��}{�w�x�=�c�b@@{��-�cZ�ֱ}�T@�n�:ކ!f<�"����Ç�1%��U��g�*�][��3��+��%��>�����@��Xc���_���6�k9@�Z��.��6�j9��ЍD��@��������QkcFރ�X۽����
ծ;�����v���.O�
s�Rs*A���`��K���H��L���rm\ ���X̪8�2�uu;t����r�/Qe;�*�,pl�n]L�
y�������4��&�� ��9�93B���!6��{�H��Z���{���/�?L�}�c��`�^��uc*>�#�=� ��\�z�E��b;��҉a�͠�\�� ��[7&����\��_~������?z��
]hZԋ5�H����(/�0�Dg�)�u3�ƍ>݁�9/0�vH�jb��;�����OX=�Mim�n{zW��5 ��^�}���������'՛r,�~m?��u.1��n�m�A^�k�2��36�`��`���_�g�)�$3Nl���v�X�'�~v��b.�k#��4@]͎�V|s����/�c	n��A�|�z�f�kʄK�g������"�
 	ۉ+7EG�ќ;�U��'�Lo�W�
7�|��鑵/�z:}�c�i5KaU�e�o@}���;�]��M�r4�o�7�j�N^5�
���X����#�3��H]��L��E�ձn���v3��Q3y��]N���4}̟`��4�ZXL�f�K�ݙ���"S�������{������U, -T�+.	T������cF��ߺ*���w���H�Z�K+
�mT���|.\50�������E���{"��M�r�����t=7��p��[60mgp� D�jz�na�����.����Ed�;���V0����]�%�M�g�F;v��dy���C�!���� n��y���flth�\.��/1�:��q��u�=�n���~�E�Z�T�^�h���4��]�vTs��g��w��E�gX���o�.��-��9�뿘����ݥ��p7V���x�y�t�}[X: .s� �*���o�q�������[V����J��_�M?"���SwJ�h��9�72�=tuj����s�F����	�����}�:�V9�}�����%��;�7i���_��ڇ�,��b�&�3�S�����>� U���z#6`� ��"��uoŎ,�D�na�b�-��s�:���D{�58`�3���d[D`X��e/
���;3Ĺ�w��F�J�c1b-��ь�k\˰ž˂�z��P�,�������l]y�}!����c��c�2�xN�2�nGV_w��T�Z#�٤��"aծC;��#(��F�o������̨��X\����+�<m��̷w�o�c����B��w����J����Iv�l�>������������ϑ�[f=�|�}N�.��������8-Ĉ��vR�σ��EI�{��=ABp]��u��!-J���zp�S�W���[ r_�|�ۭ��w��r�d����ڮ���Я.�W������x��2pu�
�6��51�b��y���-��(��!i[V+�M�����9/P�s�R)��'����)���O��F``�R��1[��<�;�˗A���@ԯ�����j��ˁ���ȣm�*L@ʝ��W��*��r�fEBT���e1��C]տ]u�bbw�����Xc���a��0|�wi�P��]�Z����³�(,��������c����q�ms����}Gە�[�u���v�૟��897C�A	¹Ɯ���[d8��ȧ.?�`}�Zc`��O�E`��yS{9a�U�e+z�U�\LY��`��W��75o$ �j�t+[����͗Q~5�j��|�Pz0-t"��F�j�'�12��8��
&�N���Kl�LX���ٌw����c!�.l�BL*��J���V�=���:�*����-cv��29x�ccB/  �����B��Բ:Әg�9^�_-a+)�헒kunj�NJ����������s*�YP���		�\���>S�F]ME��qU9UJ��P.}nk��Ab������m$�����<zN�2��ل+�ހ������v5 H�(�����< Nb������ kc�E>.����>�t����o������3��\�8�wv�����^e��Tb7IN��i ���?dZܣ$����؄��RQ��ٙ��fw#vl9����zp+���UCM�q�� 6�(4
3��G⪪á����	xE;���3V�u�.v���-��k�ݕP�(��e�8.]��Eˋ�g��`�D�G��2-�]Q�Em�W�|7u��g��A<����2>��Ѥ$5q���p���ʁZ� �sTuq���rU���^9���2�X,j�<cx��d�σM��zCJ�2���+�޵����p�Z�t����j:��-��}&��>�����n*���~c*��$�p\�]K �R�'D���aR�5����v�͊�v}jc��d�1�N�WpTp�XH��m�� �*��[�MQ8�2�J�6_�Rwѡ��7��;{�}3��#�6Ϥ �;`�h��Z�K:GW�v�O��x��{�R��h[����{a��}3T�G�6�PS�1����8~����gU��ms�XR�.���G�i�H��/�dgt�������g�/j������#�\�W���:�&��Ogۆ�U/�΀��&�K��lj��E��\��>��.<?|$���1X\`ɭ���`v|Yڶ���쭉�/o�u�h�S${>%�������������wkq&�c��.^&4o����p�����"������Ex������/H�8�'�eҤ�20�]^���̠��h��ʄpu���q���]�Z`ld��ܶ��a���{%Gr#Kԁ 3�!�V�l������Ϊ��+3� .�q��,M�ĒmH�YI�8܏�U8@ ,@w��}¦5�S��;$��h�<��񝱞M@�rz< �=�E��� 0=�f�v��W����S�\ƶ򐌠���������I�xr�T��"���k�����D�q�}�Մ8
�5I�{c����N�I�����w�P������#f���%�*�zѹ�wʏ-��T�<ָD� ⻲����Y�N��_Re�Xp��"5�<�̭���i��Q��x�Q/�ԅɳi��hA�
}DV`a��߽O�Zr��>�����L���D�X����0h�v�zT��&�s�{���w��`��wǺN�-�s��ui�|jFB�db��"����O�g���i�վ�	X��YkϢ:x��d^j�{J��1�Jjf�e���X��qZ��j�LL����b��9�Za|[����w���ݫ��ze�H��� u�4�m0��/Lc�9���G�j�Э5��q��)Cb��\����V��f��r=�Ȑ�V�g&~6� ̧�c;�ۑ�����p�V"�k�~�}G���5+Zk��p,�u~1�1�Z��*r�G ����|(#�a[�ږ�Oڊq"[	�������-��>wJ��� �L�ZI:/a�Y���W���f��X�|#i)�}�����?��4�]0�>@�BZC�����$C����BM��^�SU7����=��������j�@�-�giS/�9�Q�㎭��Z{1���A��q�{��_%���G����t*��GeK�Ico��h?@j�B�1~>���΄��$����q�����H�`{��2:ZG9�ɲ׊i�v�j�M�Kp�dܹ6N��l"�ÿ�N���չ�U�%��;L�V����b?l?��d����y����#�X
� 6K��j*���K3i9�((<ͨ��)���W*;jl�K���I��nG�m�@B*�I�I�EN��E�o秣�Q.�3UC�vR���l)U������`,͸`��1��{��Hd�M�f\B��A�aQ���Rsq�	�~�0P��G�<H(�TK��wa�u��7�u�U��"�8��N�����=�E�{�/�AL~��v�,�(h�{��,��J/�3%W���@�r��'�s

�U�j�N���Z�%Q��iR�^���G}�lB�r�Ip;��>���6�7���Bm��d���i����h��T��~o��$2��@��g�^s��8��D�LkX
߃Z��jؘ�r�'�?�6�����Vb4\Y�Sj��[��e�X]}��jKH�ԇՈad�I��S�z��x��&�!<����5��N�U�@(��\����/��<��Q\�.*$���6do}	y�㬦j��1�B���$��"L�V�{1)܏c��N�*23�r��,����7�L��(M�iu>.6�Exa|3�]&���`s�"���G���Xk��и��e��{+
��za�����a��gp��3���K���m]��B��~����P<9�k����  ��cE��"�'�k�Q9����O���(�:�Q,ˤ�0U����M^��sR���/fm|���U�����H؀�$�~�h�*T��".i��&#�͛LkF8
�b���b"��L���Q>�V��.����mc��`bC�(�Z_�܌�IM߷����y�$��;�����\��I-/���Jz���w Sf�1�J׸�1a	n��������۵��#��.��{�E��L�A�ެ2W�QI�l` �U�����X�v�u��v��(2��}��6�e������bNɷ"��W�'��7n^����}<ǆ���&������Յ�S͑ʨ�
�ZI�-*Qi[(ۄs�q{�Rx���70�t���yTG�3���^�+)��y|��I*"�9��V4�����Y�� �A��JUs�O	-������l�B�5V6o��`�]�����LİZY��C�"7Z��B��^���C�����z�(+�\�JK58$�4G��F=Gjh��r���k��f�^�_sONQSԻ�J�vL�'l�,��o:3��i��G��en�$��$��Ϊ��A�e6%ڵkCL�k�سW��a�4�﯅�Fd0sRԂ%V:��v�%l>��[>�(�xBՑxg0Z��m:��=���%��v�3�}�ĩ���KcLw�ڍ��Z�O �	_r�n�$��l���~|��[l(�u�V&��j��)�s�U6(ԃt"�BUb�S�bNP�lP�Z��F+�����f���H� ��Yc��,-�ZoG��J<T�����wҵD�B�P�l.�h8�ÀyB���e��_����&��63�df{k52�9[OmhQ��h�}{~ƈ�]��
$ߐ�y�qS��T鞽�z��/��X�����������=k���Gҩ]�	�E4��ۛ�i�t���o{���Ŋ��X����{��_/5&'��f�d�����7����SK�Z�>��L�Y�K�-�t|����9�^^_�ӧOr�g�U���&|��;��:��M^^NV�ں"�3�'KZ9����k��;0��m|��07����T��!�r
�wmG�N��A�A$�!7\���6�T��uz5B���_��w��VE��D���߫��,4	zG7�f�m�y�MR,��/���`c��,4�"��4!ݍw�c'���^�ظ��^��8O@P��ٵw����*��
��4i8�<yoɮ�Ld�-y�zQ4H�#��
6����ؔD�\m}��3F1+� ��l�p�}�yie�H�bƯ%!����U�g�;A�0F�r��[T�z��K_�@!`��G�S��=����ˊ�� ��C�}�4�)Qyͅ�Ҭ>����_`���oz��ps(:���3yAͦ�8�<��ps�_�^ߡ��/��4���/���t��/Z�D�����ϛϹ2Y��oo�o~����}̴�� ��}���<��_�H�<�!0���������&��$���I�f�������_3��6�mC�Y��m�Mb����i�D�3�M��FToe�l��E���I����s#�Y9�P7��{��D�(vGi�ȉ��*�����JG뺵�0v�V�0��v��C�p�s���Z79D��(z����z��gĚ(��z���1�N -�W�O�s$R<:#2 ��������م�^EC`v`�X������y�<i�I2�i�饞��n�l�1����1�i^����,뿝]00�%R�l]�U�F� �m��I����l�0:�{�i�؜���u�UD5=;�b���2��.�f{E�k;}�kdE�����"[pX�I��LM+�y�@Ż�Eȃ&�O�C���0�@%	)��*{��ρN�^�I��4������\�3�7��g�̐��HCM{M�\���*�;3}��Պv[�]�#��[xK���dT��e�M���UyV��	���WL�f4��V*��Ԗ9�kê
�g�����F�����	�G�O"�d����팢�V,�Rm@03�_�"�e����
���^��'4d��58u�U[�4�Q�����ov>��(i�ʊ�C#镡Dy�3��6!�-D�n��|;/l�aO԰ ���{u��B��5���iϢ(ۃ�ִL�����r���CF���ߣH2��ެ��_TX�X�aBL�/vړ����o��L��q��,uq����)xΩ��cOa�4���8��煢�V�Τ�#����U���k��4�'G��d3#S�)�Đ����,��3�j�ى�������!3;���]M��s�n�b#�.s�E2ӈZ	/
H_w�w��	���N�
�҈�<���߃�ڒ�^�K��U�-�p��q��3Ckn�G�C��v5�T��)
V�!��X&lԉ�i�l�I�3�[��R����0A�}��3�3Z��Cڳ���C@}��M�1�Se�jDQ��0b�p�>v�7�-���T	�"W
r-!���4��O�� 
�(E�<,�p`���Nr���������L��a��ٜf�7�c������TU/�^h)��|;λ�x��6ҭ��?#��_Ɲ��-B�L}�V��j�
ڍXA��g�>쬎>x�oK�KCH�B8T;=�����n���hvE����q��JHƊPS5��~�	x���A��tH�i�\S�8�ܼ��嚵M�I2H�I�a�X ���@�(y�{7�W*�),�Sf�ؔHw����r;�0�)^�����,s5g2���c>ug�[T0J�4��q������F�^G���5o;�'�K]���3,s eH΋,�y<Ӝs4��������6[�N���OO���4����y@��P^!Tx䏵9��[�C�N��=�Ǿ��>8sU`�-�n���r��-z���l��|[0�:/��r�V��3�'��#�� o]L�3��T� �&h'R�Z��$Z�(�M�����J6�w*l}z�߫%��Ή��w���[=ې_I�P	�a�+㶷6��YP��LZА�{8=2A!��c��9+KL����͝R9�z��<��;��<�%�L�b_��Gٯ�(�[7�{$�M�060쩯���A��W�LFg���:�2vzn&?թ�#T�O�gl�&�s�D�(,,��ζ>�7���v��2���2��)�W5ѢP>��)�	���1���r|�JAN+��z��_Lêh�`���mP8�F�`�ҋ0�'�{�����w+��&85��5m��i�!��j�|?���+���	��֒���#���X�Y���5��8���=�k�iA��m���5j�YǓj�X�ǿ)�$�k��q��1g����(���m���j�ͷKm��/��Mj� .�P���R���q�(eu�Ӓ�ȀL���Cj�`�p1����]��TX�,�:S�$S���c�j�C�w�+�r�%oB�2�tQ+љ09y��G�B�5��B��5#��%\�~ؼ�L*?>���@�����
��j�F��=l|V.��g������M0ӭ��Sv�d���5�k[6�N�����i��B�%�����mM��Gj@r��{�e��c3��x�xo8S`�GѲ��S�	�\����X��O����,�=��z�מ��	) ���ڈO�]������"Q_v&](B�����2��o��VP�S��x�DT�o��>C�����o�gx��4㪳2�vc������	7Uo��e���P��0�8�M��	Ǟm5Vw���`5X�iZ�B��P��Q�U�pT�獵��1�w	�z�����=���'����i��I���(��߹Q4���7[x񝙽$1��f7A8BOD-R��u�xO�cF�u��$t�
�C
/��U���ڜ5��zcHoo��[��ǯ�����c7���P��6<�/%�5�R�&�L�ړ`,�<�Y7�j	��hc�0D}�}b���/�ݷ�#���QZ���D��L5��a����K�/6��6G��{}���;&�R���輡�Mi�RƐz��m[/�ւ>��i�8\�ſ�x������[�-%�H؍�{a�<gþS2EB7�M�~�r[�ͥ�� l���4Tx*�C�|dTGa7�T[�&��N��mj:���3V�6�{��&Ҝk{�@ja�(��߭��0Uf�D��C�1Kk06{��3e[6�M��iv"��S��EL�2�mX�:��i<��'���*�S�O���m[�P�0���L�Ż�l��Ce�۸h���9g����X;�;1�B��d�����:'Za*v�`'mY];��r�P�T�����5Uu�WiQ_L��i(6�Z��53�Ն<BS��0ܾ}K���+Ғ>�_t쟔aFFR�L �����k�rU ��g��~|.G2b0���p��SM���W��=�T3��p.�~�1Oz��,�.�t
�-�)�sꂖ����F��gI˰i�<�`n�p��za��s��(A�W�Af6Tk�tđ�$�bW�j���ͷ_������G��6�ʗ��"�(R���g0�r.������I�y����_H5v'�(�Z7Fe��D���X�$�#̇�=g���M�<���k��D�;���?"LƑ(TK=`��8��g�W�з�9w�����o[y�q�o=�J��7�jo���FǋJ�g$�󫲠�b#���h.d���&�gf��S�`��hP��%Z�Jt�t\<|��9����N�1g[ B�G�F��e���P\i��rU3T�s�&�;��˟�l�X���]�5����C.>F7AM�Ȩ3t��j�1�������I�銨ܟ�Q���؎f!��6W`�����A�v�i��F��Y��v�K��f��2I���#��RR+#�8�풽�/N�����o��/����o��j�H���C]�0��Sf��1����V��)<�(e�N��{�5�s�%_Z�gƆ�{��m��87ŞiXD,�M�y������k SS��Tbi�a��f���L�
s��}u[��	L5��BBQ�h�l��L9F�3��Q&�Gr�]	�3=lz�6#�_r�Z�?i9;L4@s&@"�l�HM�a��Ĕ�K5�6����尛 �s���eV���f�H�L]	%�����,�Xl�b�;-%�
�$�����n�C�"~���tfꜼ��/7���?�I�����_n?�T�I�e4���4	f���7	�|��zW�iZ�6���{�sjz���S?�4�Vm�5� k`���i6��H�L�,�DbQb��������*2�DnA4Z�K���T��M^N��Vr��ڢ�H/g7���ę�:���
�� @E���9
�����2�Tһ�>�IY���E��|m�y�*N6ôU.�L��Jl�@��?���ȕPR2Iu Fv��ӏ5 �� ��'a�kɀu��H�S���6�=*s��]#eѢm�2�C��� jz�����y�w:%��
[s��qW����ζ5���fF�*�{�)�d^��p��<�J̯3�f ��S7(l	� �[9�n�r���E�ts*9"D|���12�`�k�">t���ט0�=5KS�����p����s@�� 0�}c�z|܄ɷ)�h�|c�_���A�wۗ�M4��sP$PMr�駛'e�[����n?���>��`��s
|�� UU�Y�?�P/�a�t�&�%�^CUDq�l��z������E��?o4�'fD[�Z8�F���|�0@�VL��Qh�����|��k.�)BJ���x`c�6)��Cc�om�`0ր�6pGf�VjV�Q��:l�S��цei�T��oB/bB�NhL�����;)�PKXpV֦%} �����u?�����F	=v�&��b��W)~�S�������m|Pm��2ȼ!�ZJa趒Z��t����R��p>LIn�F�݈����Yk�Ջߩ��j]@�z@ڂ�B��S8i����<"V�Q�٫�j�.�h�fe�+LM9}����f�WE���eH��އ'�d��tA��Dߛ�|�rB#ە�jv�2y���wg�a����E��gON=��(�X�������h_�����y����'���~.��`{�)0�36��2cp�HZS �^֙�~�cR4����禮�}-�����_1�U���1�?.6'���B�p
mɨq_f�u���-Y� �B���3;����,�:ԥF�J"΢} �x�1�J�s����s�
��/�?�g���o+���Q9�p����8Y�����-�3{uKsBn=l�`�ծ�����H�(���c���̠ab᳾[e*��@�Y\C��d���wW����bw�X�*��ZD�����֓�~�kG�F	����k0�1:E�~I���y��::�XQg��ժyЀԇ����a�p��^��~~���l��R~b�tC����
d�f�-��.��u�I]P�0�d�M���
�iբC���5�U���.�����s9�����*�RҌ��YW`Ǆ�Y-�0�8�u�0��w�
��S����9�3�D��;���  ��IDATr��l3�@m��'��N�q��57<�5ig�+���;�DX$KCz�B��x��F�|�?�|G����s{���TO�P
�{0��80.����B�f�M2/y���]9��"h:kg-!n2�`�-R�cwh!�.u퐺Z������z�o��җ�����Z�۞7��A.�ORV}3,�3�k� R�}�_s2U`<��.s���5й�$3%��`w�3U	���w�!�����ΰr���#-�S=<�΃#��1����=�_��6.a�)R6�Pw�;��0�CG�@���5�VB�l�D'Q66��
�$��9��$Ђc�9���b�F~��F�lyF��1�\��2�����%4>�_���`a!�6p1R>*ԩM�I���t�}��A�	< )�:1�ޛ_9�$Q>։��:;��3�i5�LY<zx�������a���2�-jJ`�N/^e��zx_��r���D)xA䌎ÊI�)��%����KE���ό%��P���Z�z����5��������ҙ���s�8��T�ڭ �8��b�j�9��sǑa��r���� B6D9N�3�U/G��vg"���"Ҳ���vH!H�3'#ז���#$!���-��f��������&:"�ڜ̐,�!B��>��{X�2�;{�9-�!�:��f��;4H�� [��M��B�[��q��}��u}R�|�@h��;,L�A��[��Ѻ,�Y�3`��"�;����ٛaH3M0hr��yFM��@�x�?�h��<��zO/t4�]MOm�њ�*���Z��6�J�	���	�:cN��%����~���;V+�@y]�&��b��c�P�O5��P!�8��c��d@�2�K���;<Ȩp���.�p�B*�}\����]R���I�ʄ���6n���b�8�g�[n�����,L�̔e���T��8��`�/[,f�]}D��YG�߁�b�
�T�i�]{h�PY���U�f����r�Cd$Sda�G��&6����.�67�XW����'8�I �%��l���M^`�c�`��e:�)��I��{Tݵe};�-��L�h�`>p�P��6�oJvG�v�"���) �f�:�b��:�lC�2�@'�C�|�!d?���lA����["0έF����j����\9)[W�B�ИDE�=T'sqĢ��8j)7�<��	�$�;򖺮����g��	g��9	fӋ��a'>��[�{��~D#w��6C��-T��qSZh��K��ؘ>7�m��Y��#�����X%�1��(4�3&�<ۣ�HYf+l�Y�aᕠ%����մ���	�Ff��;3�w�hf�Nkez*!̕�<g~H��T����^md!�|7e|ӝ�Kdh|wF
Ĺثc�\�����s8�f+.�.p��wYZJ��򈐰k�%fX�J�:��6҄p򠅃��_�H5�$��U3V��R��
y*R�Ҥ��_vGlK�"])��]	aGp�1gyfc��ha�a!�;`�=3�8�o!�djQQ������)%R謌�������`��^�BM�l0�`�>w�3���m������5v������d�/3�c��FMv��L�u��Y	!�-��e�T����X�v��ח5������Mp!A6���lŗݚS���~E�~����c��s�k�0�=e�Ul
�=��}��b5.4�c'(���F%��^M�V�3n���#[P�m�ݘ*��Q��2ir�����y��y@M�*�"f^F�22,��-��Õ�6��]26QB�>�g읅�T�j��Hp�#���
�f��vP�dl��gs�`si�:̎<%��� �H�.��� �&f�U��xOܢ�Ƹ��� 칹	c ��ܕ��	��cA�0��%�Kk���oe��jn����� K����L4�����@}������J�W�t'�7Ӄn"��J�wD�s�?���
�+9�:�nDӘ��+�"H(J�E�%P̹��@�jK�1���C�v.���.�`ȡ������[q7W+�"��j����1B]�B��ݰc4á����4�m��D������=xh�,��#K��8���od?����������ן�r#3B^�
LT��y�wN)�F�QS`��)U�w�\�G� �s��N:�����e[��Cu;-*+C���sr�]SeQ��5�e����gG-���O��l�1� bZ|o���0	a�^�z/d#���Z>�u�#{,��3����ujRskH��Sؕ@b(r�1�����.=��Gh8�L$i�j��-�V�3ή���f��%�F+��%v�
�Qr�p���@��(�}m7��B��o�U���y^���U��sHK�eBK_N��t	E�0^�·Q���jˁ���\6)�w���ply���]�y�//�m�(�6g�2!�y�yZ`v/�#�������N)���71����̭(��B"[ե��lf�\גQI�Ǿ1����/d���U5m�����cʕ�qsN�:r4b�ք��afվ}��[`3!�YL��]���Ȓ܀��	�?L������&r����;�p(�9� ��Sr�X��=�K����ƒ�GV������Z{��h�cxф{��ZOt���d�]�Qe���,p��ʠ.�)����G4����P4� �� �Ϙ%`���h���ט�>�>��t�
�ޡ�`��)�F�\�I��d:+��E��(��y( /M(TR�qd�r�	��2� �i%s%SQM(��ExX�/���	fR�f�Z���Һ�Jƃ���}�nP���`����=&cQ�$72#-�w�)���Pl�"c��������B+�H�J[he�(�9	��%�}�a�k�<�UVgJX3���zh�����ѽI]w:�90TC�}�Z�����j��َ4�NSn#�*fG�����R[�~Z&I��@{ �f�M�L)I�Vrg \hQ�i$����Ʊt�X�?�a�zT���ɀ-쨺o5K�i������ŵ2h��������g/���$O9<2<?aG�`�x�rg{��3��;K��(�W�$QL�@�m�h�����Ьj�T!�(��jʜF7h��Qu�}��7;�I�*5�(��m��ܛ�sCyB�T�!���c��Ĉ�Pk�&T(����"�(;�2rrf��q�U�9��6���%[*r�{X�K@�k�̠�d�LkW�����[K"� �C;n�/�է�CȎH=�I�K����허��`�L�18^YP[t��=�[��#p���1��
[���mbX�H  @����H��~�o9#a����jo��~��k%>���[�g�����T�:�%|+BH{��ԺS�Hަ��(��g; �G�
��c<0������t�Uk5�*��	����V��8����`�R��̈́qe'Ȭҙ�&���+�M�&�Dj�@UsD���v�=e���5*/%g�-T9p���Y��D�dڐD�3|�QMH�ՃF����m���Dq����pAN$�4�<����F�D�I_#��bg�v��^׊��QH������1�H�����^�l�B��w�����`�B����D��-�0�(��b�H���-ь�k1���,L��Q��T�hu~EU�����b,2+17YE��h�.SJ'�Ҡ5�-��G�xj����r�O���Xb�ff��*d���YդLɃgI�#r��9�V��
�ԯ?'��.�'쯤jQ�cUw*X:i�X���s��м�'ߣIV��?W
�����!Z�J���)�_�g� 3d^#u���%S���408����95KN81�d�ް�{����0^3� �l���;�NŃ<L�1i�ֻ5_ p\;�^������&����4��j,<4��Gj���T�֑ tc��^����X���i�:�-����kV��,�K��6��1���G�(�j�#t���`o�3u��s�L*G� P�f��'�R����d�~ �D� )]��	�R�u��ѧ'G�DA��<����I4P��݈�����X�Љ�bZ}��IK@Ay@#0�=��N�&� &
�DFt��A�K�ʕ�1�et,G)D8��erՂ�#���ω���PQ�6����q�)�7�ݮ�ӊJ����s"��9�-��cF�xv�?R����6䶎%=�1��z�'�P�;q��FEķNz;��sGy�SÊ�W!'e�'�8l��52���lR�zE�e��������J�č�l�N�ړ�����ik]��L��}��B�*��
�W�2 ��S�'ơ΢9����L��;#�E��f2ҖP���LF�y�|�z|��4RR���m�?ҖiDH� U���\��ѱ�eF�JZ.�8�2��瓘i��9�lF�z���qx]�)�(�Z��!	'X2B��]3}lx_��e���@��3^��a�d	�,ox��L��:	%��q�֭߅T�i �f���B�`�+ݝ�G�9l|ي��1�It���b�Z�T"���g�{sr�5�A*aв����F�}+��u����O�s� ��=��(^�xо�0u[z�(��J	]L�ǜ{��k2U"���İ)Y�����o�*��v�=?�j$���8x#OY!�5�*�ã�O�a]0���q����Y�l0�h�z\�¨�:��c����G}1TV�	蕀.��Uy̎YS#���8�̀�)�F���5��)4��Ǽ��9~%�(gD�ȠeǺrP=r�=����L1��sedh��Lԙ��a�<g�Q�z-;
����'B�`�s�\n"�l�4s2�N[֖]�]�^�-�<��+Ѝ��v�&��e�ˬ$i)�Q!��0�E���@�n�W/Z}�Qb�6h�ދ��5;j84mZ��em�3v�ș~����(�A��� *eV�I�O1z�{s77�{��G�bc�P���s$�1I�A����bV����ۦ�;Ɍ���,79�1��s%pOT��S�ww�66h(��Os��|~?�X����-ո-��hMJ��^gć����;�o�^�XR���r�Ek?-�� -6�;>��`F*"�Z���Xx2����&�+&a@>�}T]۵�sI4Θ_U Y���|������+ex�߃h��zB�j�T�eV�Bd��0�)�ܕ4���z�1�!�>���Ԟ@�����������zV�I��!�1���2	���1�ѵ���@����}���L����nӖ�J�o�
��br6�IU�/��F�����Xh@gL��C_����D�(��K&$�>l*l�L����T�gc�H��5-o�*?�Ę-�[J�+�B�gm��awAJ+��J
�Z7�8#,���n�I�*�Ph�}�#*�0G��N�'�h"�r��O-�z�#�;�T�4#�Zi!M��Fg���=� �U�� �ۼ��=�z��8���r���XLQ��u�|ִ�UCʽ���SS�'�+�`K�i��R
O����;V��.eG���0U��,@d�1�c��`koO��H��
"ܼ�s�'v=-Dz�\�l���:��W()��zŋ�ֆ|[H�G���PjyKZ{<i�r�hG�{���t$�� ج����K���.�"m�_� �Ň<K�e8�O�<Nz�[�{	�n əaD�4�e�{j� {�=$�_��� ҄� I�q�9���"��������iQ�'!f:�a�����-��(,Q�L,xQ�:��I�Ë\t�3C������F
ft�B�);3�`x�M��@bf��F��p<�"����aګ�z��\��6Μ���_��]�
S'�o�iZ�r�.�[��<�	�ט?󙠋%�7�뢮2O��fWJ~G}B= ����AՂ�����M����a�aN�oKą��e)u�o�����;ў������V?j�{m�]r������3�t�I�T9��������UU��Ȁ��6V�(�%QCi`a[ۑ%�Hx]��嬜ڔ�f0����a����c�ґ�YB8,6�D��d��H�ſ������˘�2�Vy���9����*AEɎy.f'-��-��`ʸӬx�Ș�,�B�bF��Ϙ���f�^�"�T�x�V)��*���Z�%��*y"���F
�L��䈙�Hb���C� �2Ė\�&�=��aK�佣���?���'B-����x�`I�=�ϑͤ��;�l���G����w=��������L��3k|�TU����y�|���5{
^�vM(�+2M����f�M���@&��-���;bky=F�%ڕVhЇ^齹~�Cg�`K�X)D�B�CHI�V�6-���Kdui��&Q�#���q��f���Ɨ㨮�l�ߗ�+zX
�@(S���,��ֲ�ƒ:S�t�l�A�;Xh5���C���C���W��ڍ6��Ҩ$du����[ݙ�f�B	+h�l�`�#�V�E�		��PB����-�7��l�iHJg@����~��UFbV��7�Q�I(߱p
q�ݴ�f�
5ģ�~�M�N@?���e-}��E^_�2�{����-x�N��2gb�=��B�zeb�~��G�#� U�ɲ�ߩ^<������Vu+�{�T!D	��?l��Vɽ8�����F��0�5��}��e�~�6��a`�y���[z�3w�*xN͢
�1a׍2�H?F�S3�w׬jU�1?���R�]�} ��1�����h�]��F��L`!��+j'�LHܜ57$��}g�0ټRZ���u/H"6g#й���������%�,kج`;���QK'=�A/Z�ǽ��R���F�%��c�6���H�m��. ��qڪ���Յ%�zΖ�{C��-ҼkO$o�9nYt�E��e��N�s᳧����#s����f��ǜ�Z��"�6y�j�-coh�Ã�g;٢M�J��(��rc��������O�׿����"�������&�����R��lW�x�$Ę�64�Z�Pa��PeK*��2\��ϑS�ꦤ�b�`�U7����P�0c��a�c�|b�e?���g2�Iւ �왁u�I*����~��':�33@��q�v�wF�u�γƼ�l�F�T������V�������t�X&��:���s���{�T�h��ɰ��ryex�&�g�ڄy��f#��B�7��Q�&����˩���V9״��p���CC�8YB��n���ݛ��5՚�����1>��r@{�`��jS�~� we�z��i��D���b�/o麻���A]�^Ob��^QŮ�2�`�I�j��g|��}+� �|���?F�QI= �>+ݹ��J-2��T-�3~h\��ss��!�s�s������ÊR[�Sx�o����j��`O��v_�뇿��I���/�r�����������l_sR}I���%�Dɵ��~�xμ�%1�a[T���q�-tH�:��og�WG�R-�bBV��+?�X��ɾI��:;>Α�_]mw&P���)�z7��|�����xF8�H5#,6������6�Ѭ}��|=o�Q��lE���\��.��C�$���̃#���G;
���wG��M@�w�.�q�����`/#���A�2�E�Y�L�eӄ@���6z���wS��{+L�8ɟ���L��Ͼ:B�� "3�?ф��ތ1�J�kv�S�s��7k	�����0L^�A��9킩���3t���|t��+Ԣ��ti���#0F��׾��%J%ު����ߺ�/�iW�>Qj��}�\�&����{����kŭKz���Ǔ2�fN�]s�ؘ @��yф�Ƶ���P��n�d���g����b�6���R��2�.����y�T)Wv�
MB��2�z���=Yb�j�,��;Q�X��� {�_Y'6�ΝW�r�(��̮�P�%:Uޮ��QVlct$��	��CVk�*�f[U��xC�����PO~�}������^�={�o�a�s�mm[y�˦�m�m��Q�OY����`ӂ���d!��Bbm=� ч$Cu��b��|����Mϻ\^�ǳp�jr:8���6Yvjj\�Ր���XO_�-i� �
�t�i�V$�ҜeV�15�;S����Aޣ*��$�{�Jl�; ��;ã`�Ɍ�F{I�l�: G�<��p(� ��cߏ��oN��%���j�9C�z�gOrJôA�u˙���dSS0�/�5R�t�t�������S�D!�����XN����\$ ��\╊Q��RH�F�eʪBP���q�*H�}].��Ԑu���eQ����b��!Uc����k��jHZ�:{�?�n5���_�8��K}C�q��ض�*�]J��ʣ�i�8�4�d�������Po�Cf��q�����\s�o���x_bf��JsY+�q&Qg2#�Z�r�ԧ��Z�hqp#�C�Ȕ��蘰f6ψ��%(��@躮�XKx�\VdG���Xr *M�>�Ⱦbe%��A��o�ccG-#p����u�����&�1�~��}-�ǳ���rEHc����J�x�S�6� <ae�#�@�k�i��D��:	/���,�+��hq��:�<����}���S��)X��F���aCɬjA\�GDh�7C�^��1���-|,��P���	�f�͋�|���!x��VO�y)BUY�~������%Լ/�µ�=�2�;`~ "��mANa��0����3Ҹ�('5tb��y�)��������x�9x��oĳ�Y�U
�s|o��l���A�`�(�c4����)�w�5���G_6�j�Rh�Ҡ�%i�
Ҙ@�X\ˉ�<����A��N$bWǎ��p~�		NW彃9��Xl33X�D�s��n� 8�Tg���=�5��<gYh�_��S ��x^`?-`��ZdBx��>�Sr���fz^]%���Ү�^��� ψ�Azά�BN�B���
���wW�Y�۽�5�E��.��������\��qԧ�p��|:%�(jP�@U3�v��M����[t/��$���mp�z�lF.suK��H:�	qL��
��C�#��#m��&��s��P#C��87VHQ��+TdV��.�v���s��;�v��r�Z�9�t����v
��W�68Ɩ�"��!H��0�T�����Z�SM˜�ӧ�3�շW8��е�̏���TO�����iN�V���;���$�]�xdC	��)�XȚPo�t�I����[h�lr������~]�=@V5�H@�:W��s �B�r�$���&���m�����ǹ*ĭy������7ԧ�)�D��I��v��0b���~c ר֎���B��1�^j��W��v�3Tr?�3�sy�>��9�(J�A��g��l�zkU�(C�"QWR2�-�o��f����������l��Q�_�}�<j��U�@�L��Jǐ�҈y� ���/���U.t*ر㎦�����sn粙 V�גr�FvWk��aP��h�(wH5mx=KNц�B$��vur��S�+����dT���R��� 
t�uRL!��^����_?]Q+���k�ֻ���`�ޡ�B����w3�x͌%	 �T��G�`��S��Eӌ�5��(�d1㛵G���m\Ɯ[�������4a�'O-0=���'���STw[�=�+�"�T�{/�_o���&ѿ�.����:�eš����6x>���vZjeذ���03=��9�B~Z�4��*9�1P������J1cQ��V'�������j7�b�a�s���1���Dt���	@�ʄ�P9�a�iK�Su5�4��W7E8�TO�X�����_=�Ω;a�1�f���{�Tb"�0���ֽ˥.λg�8��,�U{cd���g�| �2�&؍Q�Log�h���a.lNj��Pe�_.�S �TW�v�N����X 4 �OO������/�g!���f�)訜����.�}����C����<4�L���g m=� j��>��-�p9�<�Ϫn��i���ۃ	�g-�NM��rc�/b�H�}�ta���V��aX��vc*���M��T���oa����MU�c��V��Ve�[�Cf���y,޴X5�1��m|@|K7�h5&UvZ���{�����c�����n���r��.��4Y��u���r��-��bv��s?�=�;�\C��%�Ԃ2;���M�}1eؖ�Y�c�pG��Y�X�[�c�����b{_6p;�mh7H)�zFE].3AiKP�m.Ȅ���-��Bbp��E�3��Ȱ��k�Ac^>�<,nӆ�7���d�S�y�߄�u��	�ZڍC��F�8�<�KSg3����YVRUв@9j�:hra%S� S�T���z{�n``�*��&� ����4�Z�MI���!�!T�@�>�ΰs��RÀ>L*{<�nD���b�jۘBL�K��"9[�Kr5��+\���s��g���`;��3�S��p�Սi�W9�_ѦH�B-�����6v�^��d
���G{ثA<p`c-�b�x�&d�z2FU$��2=ӄ��(q�M�t3�.fȎ$}���vm�3)u�v�Kh��q]�t~��I�'�F�@�_��Qf��vИ���e?g��I�#��!�̴r�C�Bp��Q{?�!��$*�{F��{`s�d�+��l*)���ZF�	����A�1���)�о�+7�TaJ��Y~�:�:�Q�*0pV_�{��3�'V�����i���E7m��������[��rMd���H���'��Ӧ��=C����Lc��PU��О=ԯ�����U��1��tAe�YTD(�@jc�{(C���	���db{H^SK�>��/�򓈲E�X�һ^#��4ML]!D<�U�!L�*�%p�mے���6�&3B ����f�YMf�á�͕e���>�bzڱݡV��fatD�P��Ib���t�j�c�!Ԯ��l��=b��KA&�@���;�[��%
չ3 	!7��x��U@�_�NQ�m�+:C��	�˞_2��o1�1������_����{&���J
d<3u�>0�9ɐ����sHa;��<�fC5��#ưU��ܔ�U�FS�ͻ�)n ^uF�=�~�*�>}�K�xX$��
U���3��m����*�5-s�>"�deo��Y�۵j۴X?犀n�yli�
ݳp��^�%;m��c0�1C��x��$@��B�'��Y��SѮ;�Z�%�<c+�%�-N$�.xw�8�KĂ�)9|��k��0f�zrRH�%zw��Q�^sh4` +K����oI��/��f"Z2�M5bl�s/����� �P,$����B�~a�D=���D�P���npzҹ���s0]~P��瞪�)��έ%#��)�*�av����=��]��s�4m�*�� -�6����xK�m��(8�fh(0���A��Y��R�����rc?�[�������_b�ZnvS]�J��9��������zH�(E_#Ii[6,lb���Ü֓*z���%��|�9z/E|�p�z5;���jɣ�86.��*���qd�
�odS	u��3�\��6�(�G֔\�|��m96����3<Ƀ���<���f�A7V��4�L>9����ʩ�	Ɔ����'�@�1�
(uA��I/3�Ia�hPt}��fS�( �5��B�M�"�|u�9���0-��s�b#�`��y�����8���萴&C}��u�v6˼C@h��v1T~c��P�R2����<�l���.ծ pV�W���ݬP�6+�X�l���ﭴ
�α�{&{.�}^��۸^N�:x'h]hm7���~�I�O�d�#�z�}w2i��v������ʧM��^q�|FR��c�����Z�X}� �c�����n�Z �wc�w�7�����B8x�,[�U�>RE[�4>����Qm��K�*�Ɉ�e�פPQ���8]>���Z�L(1J�s	��\��u����;4�6TMd�*ԩ�.�j��lf,r��}�y����^��m��3(�t��6�A�����Q�s�@Fv�1�y8R]>����T�1��'3_ܔ>X0�
7kɉ��ywεU5��&�m�!"&�dsgYq1ޗh7a�1�J���ʞ8���Vf%�&��������~�.�o�{\(yش��e��l�HPX�#�S�h۵Ǒ!l"%�8d�Y��
L�$��1R���>�^�x�|���b��[������������m�E6F�0/����V�u����YE�B�붴����<;��-j�*r�}�p�����ZK4e���n�7��d�L)��.���+U
��*ӹɸ��Vrs�9��{�H2��cǋ u2d��,���k�� �IA�E��TZ�#f�d97�={
�0Ex�����͛,�f�>���p��b���z9�Vz�脣P��(��Xh�v�x\:����?mT�c~Q�ϲ��p�kZD����4kiZ�@����-�ԏ�V5`�����gOsJ�;(O��/�?�6�{fI9W	��]���v*���]oj�6����8�bd&�6-�����������rcb�ʋ�\j�i�I�$�Enq��^�C��0��	{1����M��*�~�.�?��@����D�@l�D����֝䎂Q*�8����������Ϊ��H1�Sڔ���#�s4V�wBsp0�q�	J�akY�ž􋬵먧�L��#�զ�uj���[
�$��/HJ��⾡C5��ݎ�#�� ��BoD� �Ղä`�����#9��Vx.L+��y����W�jfBH�Qг%M���kz[��q��K
��e��&�px��"1�O8���}�wA��-����!)���)M��q�\Z�s���TsuVM��d��&��9�*ZJ����� ��q�[~�z��TץA�7�۹ǉ�ܤo؄�l:y�:g��Xm���3��W�r����k����rC"g|���ɶ���M,5�d'��,ccܹ�I�J���"��?��ΟP�X-vM\�ʄ0�A�pTqv�W����L�oOr(�#�7��y<�.�.��0	!�%��{E�`�DUaUC�n��l�s�T���iqb�
ķu���+.[�ŗF��D�'Z���w٣��T��i��$��w��3*`BЎ��t��\/-�MЉx��nnib �O�x>��װ+c�����ѣI��K����E�(��:��6d�]ӣJNz�jxM���Ԟ�Z1�
\�V�d �/%���>�V1���E�c{�Q�#��0w�/��LO��q
o>�X8�]"����a�8���%J%�՚��Uz�ƥ���<������R�@93�����TBZ(Ũ`�T{ْ�.�07/ �b�L�`�PF(��&M����L8�I*o=�փ�z_�v���sO��>�A��e��A�=6S�ˮB5�|r�d�V�!4!��4�*����%�o��ڒ|Y�Ghf(����f��6�n��I��6ԝ���0�}�q��r���$�����¦��2�����Eo��	�p��HA�/����g�},-�ix�3i�0�\�g���b��b3�:��%K,$�mj]�V��L�,�s��=z�g��D�t�y���>%b�E�!@̄r�l��s�<|���gڔ��C(�\w�ѯ_�S�s�!*K�>0��{�ƅV�fWьq'Cd���njo�)Nzfن��8�ZT8M�J0v��0��=��N�b���ky"�P����ƶڻ��,�Z\+S�7�:%�K�q�f0��7팡��h�6��q[{h�'Z�x�&~�w���{���L���D{@��� <q����ٍ�?ec���@CGԴ=�m8*jC��c|w���ǿ�P�������O!-�:��o�*$3t���&y��o�������D� �{nv S��l�'T��k��|/L�B��7s�z,E=Z�	�;G�Α�	
4wKI;��##Z<�4[�$f��|�����ג��a��)�P�ܭ=ƞaF����9��zCh�`�(�2@/��C�{���c���T�Z��#j4�J�p�M.�~~@ �f��L�:zF[fq��!F���D�n���z�*`�traЭ2ّ~1c��n[��Ϥ/жx,�%����D�V�U�r}�kj��UX�W�M���.mt�}]�L� ������GtW�ydf泏'"�N%g('S�o��&c,W��[�XS'͑Wf������ݠ�	�"T��*?��Tl��\�ʉ��e i��ˊ:=�ef�2+	�BJ�M�4"�g�0&SCR�)�i�Be�w!'�M��D�T#�'�lR�ہ�Vj_�hI����c��.����o_Ƒ�/­�;��!�9�`�q2�3���v�v<W����x[[穑1�0߁@�ڄ۽����ƚk�K� �Ƒ��8����ct�b:���6���&�Y����#XMP���C�MM-h��ϣ���`v�[7�w8%�@��}��5��Q��2��r#���eQ��&�����|&��Z��S�ߠ�svޜwk5b}��$�J�^�Iy��k�>��eor�+�L�SÉ�� �a�sV�@���]^O/7��dt:mKк�$���A�>�ڧ��Dᑮ�o�R{��B%{�����裸�`51�
�^0�6�Z�x�BB,�Pm���ϰ�'�3	�>����^�2'�v]<��h@��0A��.�0�S<��N�J�-!�2c�є����S�C�M�����%���n~N��vJ:ט<#�Ӻ-��*j��.L�~W,k,����\I)Nw�44�ƃ��F�ן��N6�|B�n�
 ,�R������l!R`����r�)-Ju����_I{�um�R�4��Uh�5��Wc�:X��?ds�7Oc�`��w{�/_>�_��Wc��?���}����3�ώ(���dFe�V6U�K ���zDB$���MՏlh�۟&��5���S9v��>���=�3l"H"d�I�b��&I�Mb+ƚG[~�y��ACh�1y���T��V-旑�5����9$/<�=$�ޙ����G��1�a�Y�|��ފ��m�٫�?�4�v<IA�-|�����o�.Lǁ�ؘ���5��6�����eO�|2i�Yo�1՞��N�h�j/�����P�4���l�,݉�*�]3��5W�!ñ5�`^�fE��1"��h�?LZj����`��MH�����9����.�U�	��N�ׯ_������o��K��M��g�x�~S��E�l�筧֙�
&�8�fÆ�{�f%��V���b#	*-A����*<C��=�&���d�$}����s&p@��k��t�FJ�*RڗZԎ�J BVw�s���A�(�����/rp��zK��f|`F̘E����.zd���mf�`��n;���}��]�T�X�,� ���f����dt��xl��]6�N�R�,��g�6�pr���-��K��0���W�2T��SU���S[4�0�{��o��;��Z�
a�qn����YǷ	����*�=�<�qKhH(`�sG��e��,3Vi%-du�׎�?�xC526�(;�Oʟ�|���bR��uJn����^���j�6ۓ�=��ç�9YϤ�ʯNU/�a]�����y�0�^:�Q��$DJR9��\L�ɞD��vs-��v�S �\D��6q2�Y��;jq{�ޭr�s�Sի���c�!�I՝噕 X��3����A"�pږ�R!m	�
�Ea��4Q��_���Nh����A�X����`\�(�c�V!`�{x���������6�hO!�A�`Vq������xA�~~+FL�0��N�̈b;����$�-��5�^N�6W����e���c<��� =j�A���n��jw�#��K�-���=�[C+rMo�g8�,��Ѕ� P���'���C:z�񴮧3�K}s��P�/J#��t��t6O��ɻ9K^n3u���.��ʷ�{�+a��~��ח �Ѫ��(c�t�,H��c3�����6"!��H4�y�^�����*ŘPJ�blD�gb*X^;g�G,6�*�=y+�?݆��Y4�qڌ�D�Y�(�0#Pm&2�#���
��*����'Q�1���A��;�H��/�/֑ޅ�v]�tDɊH�b'�MA�z���a���9�IC��k��s�?͢9��R �
�$W�ې�(&^ڂ�nhk!hB��
 ���ɵ1�� z��LD�W��g8t=j�`��y��4q��(^y�s�i�*�n�y�t��j@�]k��}��=G�`���_��̄���_���X��y*b���̟����E�Ү�����[����P6M7��Xp��o7)�.V$EQ��6��/��;i��3
�4R��I��q�)"e82I�j������n�mA��F�ql�"TI�b_�����Bh����N���FfDa�ޣ�����E(�?C�)
�p�G�;QV�����=2rz�:S�*��m��Lʖ,���^��HF��ϲ���Ÿ�wH����X�9*�!�@o����I��J�-8j�#�@	�*�m�ns0��	�z]�iT�5�,��B�84.V�"<��Τ#���q�PG̱;�|"N�f�\k4�έ4�V�Q�(�,y�-�'�
��)v�E�%2jiD!�	a�ӱj����w/�t;O��_@�W����Oϫ�/���Ž�ׇ�@��v�W�h�*S�p�C�*In���_n��f��ʤ�y��m�n��8�nz`�5 WS;!�ň}`��y�n@��w�A.����a�nj"P+���s`d��-�����`#���	1,���l�T�?�/� ��w@�@�@b��ñ���lF�t�̾R����G�"��*�͌�_0 � �����t��;#�]��������@�{��V�]��*��F�y�"?��V�M�^�W���,aO��N��:�FGW�_�����2������Lj{~%�˙n����#yMԹ�EO�p��u�ۼD�X�uBG4G���6����8TV/����ۛw�Ժ�C껕�R8ne������]=9N�ʤ��P�n*B�`���'����q1#���;0�#3�q�aD�t�;^'���?�����ױ�@�"�os=nA}��~�N�Az�N9������k���
�����t��`?���i��}�d���]V��u�}�]���9�������oɬ��Y��yB,,~�j9�ܑ|�`Ӷ�Hj7�����Q��0W�92��P�=P&�}�uX�ބP�xw��o��!��0%�uJڱƂ�l�}��������f~�]B�}<-��%���B>� �U�iqZc��k�b�I��Y�ۏ3�k��K5�Í�&����/�F��ɔ�߸���M�ο�X$�x�ܰ��f2]�i�`��E�����9���Cf�Ϧ��G0J0�R�ټ!˳�lm@��y���屧�u�-,��4�L�ĄV�YϲwcL�8c�����%[�0����V�
�g8�u�ю��Hr�:���0:�4O�}=¼����lˍ��<+��>��x�E����>4��̬h��֞�-�G��p��S�-+���E����:���*��{�C�o�P?�B�ۍ,C����s�ַ(ͦ�e�t������c��B(�p���B�CHU�� @?˵"�p����x����=�S�%�z$���#���Ah�8� ���#�q�~to�g��.��+d3�]�s(1]'Q��z0+`)~�m��uS�����@�yA4��3��VF�
��0�r�Y��N���!i��d+�?�׼�%��!��)�T	�l�3=�����F��"P,8��?'�0�����:��7>�[�3�<�x��/E��R��-�b��]틭Z����u��q����ƪ�.V;U�E%���2Ģ��A��G(�Pdkɴ�x����#X�1ڊ��w��[؈`�����d
Ta�3#�[4+�(6�:�՞��]�s*�9�����	1�dic��r�C�6�-��$���9����#��K�k	xyL�����ga�a&$�4�D�j��4�g��V�9^ZEs葎�N5_K0SC�X;r�,:hXc�1���v���[�{��[��������xC�#	`Qbb�`�~�gu�-Q����fZ�V7$�����&#�ǂ��J�f���m�E};2;����������ʊ`q<�C�Z��Xyc��~�~�� �Ŗj�l��CF�LzA����]�W�f��bF����o����6x:��Ӌ�8�:3r^�a���y>2�ܼ�1��Q������q'ظ�̱$ Z������Av����B�$�=��Q!��L�"J�%�R��`�M����Wj7P�)Lo�9�s����D\U�+�F��߁fb6����A�5m���l��<�x*C�NJ���e�/��� �k��Ѱ��i@\Y����OH_�m���u@�G�d��2�g�6g���5!�)t_�{a��s�Җ�k�PwvC;�$[�G�{'���ɇ��JU������ILuf|��G�:����(��\����Ym�Z�����7�k�wPM9yd���lS�P�%߇�F���G��Q<�1���q��F���L!\�Y��_�(���[;�kFM�m�����%jO�j��rOt����_Y�W)��*IχM�Z������2T��A�T��E���Ơ�+fT��أ[��sTOW��P�:���o���B�#�=��Oz��<&�H4�����|�7^	~a�"9j��[�^�A����1���� �C"S�;Uf(�`	�pf��;�I��8w����=0] �����\�=%�4ց���Z{�~5+�]2hdL�U��<"y����9���w�1'�Ě/����x3���y�Ƙ�бO0g�EtNIg�q|�yW�z��c���ؾ�|�.-�f�L0q�b�8�
��b�#��;�(O>��Pk���@������'���f1��o��N?�ꔵ���x����xQ-�G�/D,t͑�.���kB�|O|wDw��4�2�.������T����31;9O0/"k&����`��Ӏ��9�J�x�3zVn���e�?��nd#���ֽ��4�Ŧ,�'��GJ�ǌ)�n�q��]�l�
Si^��53��>�%5�4#D3B�߲		��XX
�{Y���7�<I�345�._���u�;��FH9R��� ú6I�5:�{����`�ǵ|��\�J�tL���P�a!W��m����o'}R[�����Q�rC��k�^�����礣���k�X���7y�l�����c�G?z.�X>������Y��8	h�����9D�����z	S*;�z���c>�V?B-��������N���ȸ)�bT����G��Fs��̿�<'&�4�qެ�'�$h!�=jǲ��($�����%	AS���4�Qs8�֘7�Bљ\�(p�댽�eS��xwjQ���0����֏;{7�0��8G쥺�7A�MIC�����*�ќ�i�����ʈ���tЙTy\�O�9u�2c���;��ʱ��������ϙw��(����|:����!ʯÁ}��}�L�Xr��C��db6Iح��w�ϱ�\�>`��꽔sCH�3������>
�0��xE���.s��4+c��Z7�"��D�b`>_U�"��nxF}��FrO?����j2T��,�+��tODo�]aYYR
�F�t� �*g6�9؎�bb˂3�̰��Q�,"�Vh�Sc��X1o� YA��& `���3��W��h}���0�SSO�Ӗ��/�G��f�����*�\Ė����^�O����M���낼}��Ջ��.ݔ�K����[b�H�-��{iQh%7\��&][�Ϳ0���)f�`1!��0�'�H]%�g�ji����GS 490�c���I�[=�-��r��c,���_r1i�y1+qU�P�+z>3����fF�?֙�ޡ-���"���dz:
�@jo�sTV���*-�V�y�O�}���١յ�nk�6���G����Tf��&��ZJa�e!��a�$���Z��=�?E�	=.QuL�=�$ kݲgq��GfT8�Z`�|)j�/_�9ޒ�iD=��~
�TA?�n��x<�����jQ�L��^#�z�w��0u�2^��h{�{<��-l�����p>�5%?��%��F� ����=���Ẽb�D�w2:����q���m Hvp�րg���b��K:��d��� ɽ����Nt
4F�Ȃ%.��B�|��7͛�/�����Ѽ�G�q���x/��#E�L[���ڦ�Xe`*�����B�
�3�D������&�2$�-h���<��a�e��l$��0�i���
�У�iP�֭:V&������O��/�y�1�v<7l*(>5��i �ZF�<[�~6��p[�H{ǰ�FS�?�,�ڠ�	F��p�ad�j�MUs�Ck�w��J�X�
�����9�D��	�S���#��jc��a�V�!����0f~7�L�{p��3M���}��y�L���gX�����h���q`v�j�z��5ң��(���(�OR3{�d��8l="���	ƼtCC��Q�}xI/6u�s�c=��,Hԗ�4��tL=�Ǚ�a����^�����쨪�&��,�[T�������i�H���㩙R��؋L�6��PE�Q�rS�O7��!"��7���L+�XRE�h@�#����z�TE� 3e��bb�!&�,BY�]�e�B��w��o��L���V����R� ��XO�'fu����'�ȉm�@N���� �Z�q��|������\3��4�l�MB�nn��A~w�e#��L-^}�!28�~\��>!Gs.y\�v��I	�`<TM�����@�G�奔��I/��V�j���G��;���s0�J��e�!����u�`boHn�C���E�%�Zo����W����Y5�(ş´�Ê��K����X����lD�r��\�Y����61�:�PI����^��؟}��YH82N#�;0��j!3�f�l�19@f9M����p����&@(1��Ʋv<�sTap�[��;b|Y߀���P��9�4���Q���x_�25��=�o
�����q}�������ݽ��KMW|N��MUo�g!�يwm�[���؟�8�kZ��2������ {n�边1�S�Fq8fM��
 ǒ����3� �n*��z6ț׬�d�N����ސ�ke��z��6m�;�t@$�p�c��v�V�B��S�;�&�/��̔�U&�7W�������S��m\����� �9sSa�e��,�'TH̛�W#���L�Z~����լhGC�q@���=鞌RM]G��i�87��fj��<�u�E�ѻ�3H`�z�7Ơ���&�4��IQ<��Ԣ�9�]���9���֨����=��3Tܛ��.к,5�O���V� ��a���S;�L�	|&R���7̗~��|�*d)	MV"C�n�E����7m�$ǱAUs�Ȭ�s�WfegDvV�����/-�[]��nJ��x�#M=�,�.��0wӋ�� ��'Q9���z�/��~��1+���X��wl�f$�ʥo�>�	��d���2�EY����4����ֻ����-��"��_3�>J���Q.���$�����|�o]�2�E����Fj?��.�Σͅd��m��U���T�zO��K�%#(d��7T}�V�)3E4������E9�^X1P� ��lYϕ�s
Skn�����Z�
2�iv} �4�L�ԗw���_�f��O>����r2p9 >�A�^;)|Q�{<~-s�{'�q����i�@K�S�1����I�Z�gq׎���}G�L��[k5��Z���@` �qm[�13Cߍ 2�2�r �aiפ~�!)!����[������(��7�4��|��E3��c}����:>�
�Yq2���̀v����5������AN�;��'9	Y��������DJ�#4�P;���&��^��FP�1�V�F��Ms�V)�u��6����A��瞌Ż�]!�~O�w�@����F�$�ĪKJ�r[џ�~o|}x������j��\�:Q�l�=��Ou*�ڟ�wtD�dҺ������PG2X��0�0��
I�f2 �@m-լ��4h�����ێ5 $�*���Oq�Nm�1��Ll�'s9K�$T-��n;�lx�	�uxO��H�_(g�vi�s� � �V�V����0f�A���W�+ege��g<��N"6k[K�8kw�{�%�^�%��C��&��ڔ��	I[~�4)[�?�����2н|2���o5.!R��ֱ�c�_��n�����`q嗽�MQ�}�K?0c���%������� ����^WG=?=�����'�N��*ǵO�(�� L�Z��R:�����300h�#�,B���@E����}.��{�8f�u��7�֖�Ƴ�E �=\fފ�6��O��SF@̘�R���}��ڌq7a��'�[��uQ
h�S����oj��9��6�8���/X#�M���іvD4E���ܟ��"9��[lm��"B-��`��%�g��퉊�R۞�Q�\��=�)��RwUP_��ǧm�9F�G���c�Ɔ�QG���d���L~�֮.�����N�,'�n�DW5���0ѡ�)�V �{�;lS֬ G���<��]�dCN����VF8��-�֨�YN���0)Q�	h����vt�]K�]N�=#�˛�-�)0��)�W�� GL��w����D�ԶV�D�v[�e���L2�h���u`E��t��4�Q�^i����$�k����!-�K�3�'���߷��$	َ����n-��P��E6�O��<�L�8��Pp����#��n��5��J�� `��>�V9r�Z�h"6Նw�l�O�`:�k�����PUt��ņ�w����E���g�x����P��\7�e3��y�@m��| "�(�7��:؟&�
�h;��Ŧ~B�u�cnqO �1��`o<��](����6�m��C�o�ɪX�f�C�w4����KO�.̡γ�K���hp�����d� +|����SK��RP&�`��)O2�3�{J�]f��*�ʐd�C�@���"��`C��;���[��o�\+71�Y�s�)�k;z���V��~f��W��Ɲ`l� Þ�4jX
������PEr�O����\V���r�ɻ2�����EtA�F�;X�wX?�r�<���FZz����ouݲ���;J�
�1��ۍ��T�H���[��w��F`Nt�EQ��"���2�<)�����>.�a[��5בZٻ|l�bʭֺ��z1���XƠ77R#�x�*p�]0���
�xDֹrhj=8�b��O�3P�-�(!W�E�x�6�?�X����@��H�V�,`20���r��=Y����H �3���g�[��*�G����{I�)&C$��E�^K+
`�L{���Jd0�T�h�\p�c %�� ��oQ8��z&��!�~ޥA�7�ҭ��e����!O�����7���x1�*;� G�
���E����٦ܤ3�
 U��T&H8������Z��~��b�PL�/��ɦ��Ŧb ��YC�w�[�D����`��C& �%���C$�V�7<�XFp���-rN� �ȸUf*��{:�����-�^`ΰv��hL*�i�rU6�9�y����O��V޴e�`�,�ˁ�F��������q�նX��ʄ��>)<n�2���(B�q�@�%�h�� �>O� >����̲=�����&�)�&�v�C���*�p��u��K�� }��)�h�z�u��KZS�-A2�}+vkq���F�`yx�])��GyE�\�u歲Y�$����9��8^�W�y�H�ǫm�䶔������WTe=���F��t<؇ھ�7A���"��Q돓 B��N�z���ec�,�7�>J��ĳ�|&�D��4؍�n:���<��qO���Tl���w�b5> n��e�pzrh�i���2�m�u�p�o�0��G��"�P��4��=��QέWZ�������[b&Bmπ% �g�<=�zP�|�M*���M�1��0���ց���S�vMfo����KC�5�[��� �}Ꞃ��]0h��m~~d7+�k'��7Y?�d�Q�N�wf[�  ����RkU�5ν��0�:���Z����(�u�;������'��p�X���t�98��3�4�^/��d'd���p~/�/'��?)�ټ�^�%s�u쉠�/5wh�-Ι��;��	+���F	 N������ ��]��{�I+�3�ۿ���:�&��c�Zi�㘵��hp�����\3,��Z��I�Mv�\�	�$�}:Y�|����aWKٓ�M�-ӳ�v�]b@eG�1��\]���.��y|�DDƘ�g����+�N05<����;|�b�Gl�����f4'2�Xt��C]7����9��M��鎌P�*�?;�����ZI��X�M~���%�M;4.��,�o��ᬕAe���}fQ�Ҧ ��� 8�A�
���;��D3��9]��`����&v97�4����2�ao��$�yӷ��Y-MH|�A�e��^D��"��H�¬9AjL���v:��ky�e%��(�Hƴ�Uu��lyUz{N��n��SΊm��̴3[�db��������tM��z����W�~1mYb��d�ɀ�rPnx����g+����i�*qF��?��������]�z����.͇�w�ٲ��L�-�S��2T` Xِ3�w����e�;L"��� V� -;��)D��E���BG2�d�����&v����)4�X���v�9F�K��1��4��2[X������P:������w�3�΂٨��Z�N�" �EAL��2)B��	���8a`Q��ދ5��S���\UE��`���U�6~r�{j���k�*7`���`ڻ���US�кD���Cū�.����Yx����.`'���w����P�VT�DZ��q��p����_0 b�<�u�؊�1��f�]V�A�Rm}-�x1�͉0�$�/��WK���z2���t��ܒ��g0����m����k� P�g��/�a@��l��
z^g?h�����j�1��*A�v��0�򚼾M�����#�!�(� #�a��%���*7����>]"'�IfS�.��1�Ysf���T�q�w})�s*Ѩ�M�"R���'�30���',𴰠��l�+@��?혌��v(��p7/������] �k��FoM�Y�>t��G��ܯmk2LҌ|����>t�$v[BR���:�=eֱ����Ɉ�o�3�w�l��v. ��b��q�M;��6T�4��;���� F�u���lW�I	�`M���^{	 �׎�O3'(m�����"�i�KXY��d���	Р��]N1�}޷4*��Mr��U�3����CF�����Y�	cN\�/�o�jQ�Q)��<c�Jj�ű8o0���'�=?������?1!��<}�%�N�u���m�����y����_�������7;��; Nq��`� �b�.�|C �j��!e&O�X$3-h���>Y�ȇ[K�53�;v���& K������f���ğ&t�l�V��=� ��X���D]�=��\����B��}���QC��2b2��X	�rZ���O`�:�(p����.�⩏����\�Ʒ�bL9X-���.r̊tʭ��O�!8����h�1� ���fb��M.�3�%��ju���O�q�f�.[.$l�.9{�{ #G��÷E���O{�����r����Z��1���ƌ٦ZQal1�flF�@j$��!���`����X\i�ü���ϗ��@�@m�Yv7�갆�轶�]Kϭ���Q�l0��j���J�I�����*��i� [A�9��^�2��2K�@�&�F]|Y)�&e�g��zD���O�9Uq��{1_3=W\)�1Pb�k�۳BΊ���3�����u��I��#�qY3(�ƨ1�ST��q��K���[(�d���UuC�r^��Qɢ��!x���e�O[xq��c ���ɻ�@��oU��j�w�������o�1��^�������@i-3&Z|�zTCJ��r��E;��H`٠�z�C]���l��9U���2�uǢd�O`�� t��x�	kzN8k�s���S��3r���i���z$c�2k�j�~%nEBqg�^~<��6��S�9�Q�6�"��޵���#㉹�0�� )�� cjGza���K��dF)�T�'L����xّ��s�=<�E���wV�-���YX�yi�ڲ��Nr7�-Zz�w2yz�@Yd,[� \�
��4d�B�������>_���
�����2�=�8�����p3����z�O7@�W �FPƪf�L������̥�H%g�`�� ��S��Ҽf���gґ�������d~.bb��`�cl TKge�2�i ��b�CdV��ic~6�J<#��
���0p#s[��?�\�a�H�/����X��%�����t��������Ƌ�և�¨��-�4�)�AZu_���@��J����ב�B0�(k	���h����t��6)��Kfl��Q6}��mTm�"�j��	��=���K��6�/����CC(�P��Q�gf����l�K���u':4Gd�ǀǡ�+{t���2�{���H���i�Rl�­��,��Ԏ��ކ$��O�z����/gv��P�^-���� �Nޑ�&�C˚��Q�x�� OA������--vG�z$��M9m+�������e[A��|�`ZM����M��^r��!�i�a���ؠ��p�Ȗ�^"W�wZ��ϲ���Q��]�=��bnۼ������u��^�J�(q�#�4��-��?ͺ��.`3_*a3�܅`m�T�B����[i,�c�fL8�k��s8ɸ�RtS=�9�64��۾l���a�Pͽ�W�rn<��]`t阱�h(h���_��_��zr?��k�?|�`����%߹�V��vmHc���̰��˝� 4�����g��L�B�>b?e7�,o@1;d�����`�о����?")�iO�������Y�3gw-tu��s����`��k����v����X��9�0b�k�&��waHZ�xͼ>cw+�z�
����R����Q߻��d[:��׼�A����Gkol�zry0Y���Q�BvF$4����ۈ��'e��0��k���k����=¯��6f8Y�ʤʌޯk�5��k�K�j��"ë]�+� <���Ɗ�=�xX�>�A��<�RG.�y@64	���}�{�0_�R�#ˍ`^�"W�O���9�ڗ]??�^~���|����|��1� �M}����~;�%�h���'�Vp1�D�4O���~'�?}�O7�_����Z�8��u���.����A�蕱�M�D3�ׄ�ff���lG������4uA�-ٔ�Z$Wix�5�c���)�Q�
oa���������a�)�@lqu	`�M���6<8��t����6��WD��з�m)�s��7���C���I�U(�'�m���������r��038�Y%F�z�r�F!OVOu�ȞTj��=1F�#/��	
	�m�Bж���K��J�\v�+Rl���Y����`�8^JD����3u�[n�V���
�{��r����Z��70�駟�_�/���Nf�;m�'	D 3Y����W+��S���u��Q�><��T�4���곏��fd��߈=f��B����qy�LL s�̀b�Ȯd�rL@���#������ut�Y��'��0L�'�������F�=�N�i+6���6�`��]�	�[��#32��H�����C��6�
�TQ�TD�k�L>OE��:R����^"��t��^m�u���!����2m�A�bJυi�	KL�Z�5��I�G��>����~�muln9j�JLeėh>�X���� ʓ�D|�@��M
e	��$��$c�zd�!V���dۏ��E�)�y���H+��r�en1yc���K�D��Տ?�(?������SǑZ:ۍ]�5c�0�A?L��{�,��uLɉ��~������Z_~���z��%�U�f�_<��эYKm8ͫ
�a�3o%�Sd�cM��7i�~���`��ɿ����X�T}����R�L�&k�$pp;�v��J�� ���u�9[�|�	ܟ �_�TRIրxКq%�Ef	��W)?�}�"���[3�]��\�YY�D􀸩8�/g�"�۷wA#����y����&�M�����E��y���00ԉ��t1D9�H� �zk��;����l�9h8@�Y �2�y�)�^��%���{�7�C�D�0������8o����T(6.Z���� (�u�-,����U)�*�� ���}��'>�x,CM�)s1�{7m��/y\z�j��?Z��(7`��9(O�p��ˋ�[�s16����X�#)�w�Tb�;�5�94�A[��4 5P$fQ�>U(��L���lD���{�k��
[!���ڰW��Lu�v�(s�A�%�޻|����=�MLJ[�O�D��Fɜ���Sk �������~)6������K�,g����ǹ�.�����L�l=��}`ma��ǧʻ�Գ�Ve*B�Ko5Q���R��vL@\*��.-X�Y<� <��u<�ˇ�:��}}Ѽ����H���s�{����_�"���nf��L�y����=��*���2�͟�U�L=xR�Çg��
�zaR
�NU��ٝ�,  俑�؉�=�� >�W��{|#ޕ3��~�΂Tۙv>�Qp��bFu�k]~�����Ͽ�kL8���8E�h�_C���f �R�a~�1��G]20��� �Fu=b�'�ۼJ�M@�&����I�`�2·z՜�G�0Σ}� ���o�ư�
�G*eg��&td�9B1`��5�!E2]K����G����
P��[�m'ś�d��-�7��!�}FiuW�߶��|@y#c�o�rM_#�M
32���ǋ'��v�P�j����s�b"��@=�-#���-�c���&�p^��[D��j�mQ�n${�	�n�o����?�Q���?��~�Ӎ��NfHf�͞�wy��.>T�$��6�D"�1���/	P#g�L�F��&�	��r�F��&��_���iY�(@dF�kƅ���[�yY1�d��0��	-���3�T��׿&y��G�m�#�p��[��=?�W�;����(W��Җ�,��1`�x�"}}Hл���V�+(1;�c����D�	��C3�Orc.�mL;.�k���>���K*ƙ� 4�e����͔��Tq_(�c��n������	�IBӊaAi�d+&�%,��}��po �n��D�����r��[={ж��`�0劾G�VZ�Yv��R�k����n7�e�"��ҥ�y��
�7V �
�����At�,��2����(}�+���x�Z�!�[鉝l㻣��nbW�5���L=�=N�����>%���,��s��fb�dZ��[�#���!��u�U��-}��Y.7!�=r��{��x���ۋ�X��0H�|��/dM��~:hC������0	1���9?�>^��ۜ4ʦ��P����.�$.���*��)���-���'V��?����>b��7���Bv�:	��A��> �q�~Ы:M�x���4cj�}�iԘH9b$�1��IW��t�^#d~��;�c��OX��{�T��8U8��l&7z~�2�@ 8U#X���[�3�"�%���� ��X0ѭ���}���-A���E)�:�ź����PaΤ9�NZ�D�M"��VB�{7Vb��n�x龥���1�þ�
ѩ	�|�	x��*���x۠�R�u&�gQ�ıZ&�Nˎ ^��;|GLU4��_b�g�%Z������_)��4� 0�@���R9Z@���Mq���ͱ�~O��No��� �T�aJ���p��l:��v%�]@�@EÃw'HB
��|�%���7��bl$�Lvo�����8 ��-��}ߣX��}�2��"��{�w�P����SNX~7�X?~���P�b�[�"MĘ���lQ�R���z��~z�~�}qM�0��^�V�ɂ���l5�<��s�#8~�SAh���X[�ϛ�d�*��t�������3�5�&"%���>`���M�� ��1��i�h��/������m!A��b�\ N��Ñb[0��N��l�J�[,�Y>���g�WZ�ä0�rv�����l6���`�L�r92�6A�C��V *�䃵ޞpH<����td#�9�_0zS\:)�O)���E�j�a �� F7')W;BݐTje'l�x�s�|)�P��dF_6�J&������i��\*�3X�a��)�������)�j��2�g[��-a�� -��o��W�Ev~V�bm�Cc����ꁥ2qw�ڿ>�]"�@�Ј�7�l���wa��&�������?=C}�H�%)" �'{
��l2�� z��塝\��%X�M�f�+�:�߉���u �Bbi������,��h˲�>r��ol9	#1���`گ1S�W&��,��ɟ�gmU�S�OF�0��E�{�G)3�i�����
nֵh+X��Oqk�5l_�L�rZ�@��/�J��R�p�J(�A���	��$�i�Ba6Y�A���3��L(^f5�:Vd�Ǭ@'��N�V�ma�(������� ��	�KȒ��_srJ�2�s�ٔy)�`���,��)Y=&�J�L�#�D�weވ����GY&��~Y�-rY`��0z�oO���G���<m3�ȝ�+����gy_t<P��߭W��Z4n�T8��S�2�hWQfLw?)h��=X0X$/��!��8γ���N>"W�������6�b��~T�7��H���l>T�~C�����o�Q�#�F+0�@�6��Jw-^Mv�A�z,��-�9`>{�k����P�b��bx�Э4�9h4@�XR���&�L&��ď\��Q��^�����q�5�T��>$4G=W�jZ��Ǝ�XI�ڴ �-�ϖ^ޔ�-�?��z��R�}>"w�.��e��T����֯�ڏ#5���9WI��Ji�rD�%�O-���3-?iL.AywX�=Z����j>��{Y#V�"i�+I��.�'��[�	� g-B��#՚&@�g� �=��/ C���vb��V�'�L#�>�2�`_Ua�m��o��l?n[��?������C�$�:�#�]�,E�i�&
�A�S�m���V0�\���8�>b�U^>J���� �ۓ%H22k�`6D�ꮥ��m $7$�˛AD҄�?vd��<� ��K�_u��
 O�3"���&�D��=����.�dܣ����X�>࿌o�߷dN
����m��h���X)
 m�=��1mh��Z�xt�G����-��8�����<��Y������ ��P�'5��}s��=�e�vT��Řn�;��C_�j��vuM���L���\��e�q�K$p�c�����rR�'���x�݀�2Q���򹹠�l�p�x�̱y�||��?J0ܩKZ\C��5SO��´��ڬi�W
kÄR�&|�L�2+�U əq�>L�"|y\��K���XP�n�Pf�__�z�[���~�Y]����?��#�����CM?+c�ml)mF����%���5�]�Of,�0�e�$׼{-�abD<]��wmg��4_F[^��x�0T����0�NN�%�O2N2������Ϥ#M߯�uŀ� �n�k�L�M�lP��b\lUˣ���YT롷?�,��o��[��n�:!��_>锸<}|����g{�^>^rr������[���K
��
��J4_��$!��S��aB���qX��{�xk�  ��6�, ���C.s%˷=�MԵ\�x$y2���� P}��?�:��������,�z@�i����OI�5����r�3���7�)��Pp�qWҬq�u�qhUfU�~���r�3De�b�.�Cs��LQӹ7f}���7�Kۻ2���P��Dx\*G�A�N�6�3���e��2*	x��d�,K;�p8;�tg䤤�O�(Hs0�b�c�l�ltd[�qD���"���duO99��_��l7�K(�`���]��BH�&��CN��q�p�7�y� ����e�w��C���b�C*��C��,�~Ǆ�*U�6�g�q0i�Д6��[���[����1F� ӿp� /c���O6�(*���N�Q�MD�%���v���P[�F�gs�0	h��1�>؜�h�Q��M�M��F����E�p)	ځ.p��i�����x�
�u�eD�0`LW*���ā��Z"v�8�ov��j0�+�)���ƭ��9�2f�	wd��W�����'�cw��xҎ��C��M����el^���P�seߊd
��Ou��%�(�swv�d"��}����e̴E��q����$*zN���
��^�7�W���L�)���� �J���
���	��I��MMFJ���x*=>[�g�;�)b\�pg��r���X���cxR����iqǠQB$�qj�1r��czy\�}��o4��.4m��O�4W���Z8�A�4�4�,1�l"�{�HYA,������N�����$����$5�DVҧd��^�	�fϋ�W)�)��Z�}�l���@ 0���}�
4{���>����F@���/��n��SB;>�ܐ��%��!`�(Y�ٲN�v�N�35�yS�u(]�U��z�/ٴ�~[��j	��
i��U�31z�4֖�i�\9�e�ZZ�T�@��)Ֆc������\�%#sw�N߅%�vAR��G�6Ř�?�
S�P�V�T���(4�)q�歲]z�Y��fo�f	|��ӊ�w���˖gK���h�uR ���U�=�������w���"`c�?�ی,:�5�&ǐ�fb��a�}����s�-1N���f�����H�{Td��(�+52��z�$�$ܬ�Kю���i놶x|��K����ƌ�v�K$}���`���_�`s��U�_4]���~�T��@�ա�2lj�i�`��P �rN>�6;��M�V���GI�O���VXkyO�O)v*�9'M����a>T>��K�T8��g�a�όr�.�Y_���q~T�$i�x�̿�,�O0���c�T���Yٷ�~O��>��� %X�H��	0�w{H��Ђu�b��I��w�!��V��ZxT[`��1n�&׾Is{��ϩL��&n2	ڒ�e�\��7ڣ���heV4
�sJF��{��SA��2�~��޳��we���KvI���V�~dK���LGd��c�2ލ�7
�"�&�j���RC��"c��� �(?L�ON&���MKd���~��n���[���B��:0f�G�f�X`o�Ȭ3�ԁУ�G+�ͯ�$���3P��Hv`�|����16�	,�.�HZ�Ͷ�r1KY�-n@��-At���6�g��!�y �s�l{��ʑ�U��\Yy	��ٶ�Й�-:Q>y�dbuh;����I��
�i?	ψ�(��j�d��PC�݈��n��� ��lB�@^�y0�g��?a��r�o���˃H�)�8q���'�h�<�
 ���ol���d��&��9,&���=e1����\�w5ի��w����^����XFL}4+��8�q�Ԥ[B������j�B��Z�����k��$�	� D^ő-s��<NsN�AY������׳9��I�� D�U�Q1�l�js\�=����]�ek`�������˂u�>Мa��bk��z{n�,0h"���V�%�[X�=�[d g#ʭnfm�i��|X�٭�ks��+/%5���w�J�r�
�΋U&7J%_�s�����s]=�6�@?��y�%�˒�MQ��j�{ �iS}�%����kӸԝl��1��1���lp¥J�D���f�{j�xn�V.�b��zy����K<i�l�XfI��Q�d�U?9�G4*��Yj���윯!fg�nQz�~4�#�@$H�|��M4�S0��v��=Ǒ^�r������P�2cP��͗lJ�ٌE�(`�iy� ��\���Y�$�# �����beQ ꁄݡ�l���zS�k�i��ڗ�f���T�%%Z���,e��P��ᰬ��4����Y��~��a��K�h+� #÷^^�n�s�ܙ���9���!3B��|r�[�yj��^	��8񁞱>6�n.G�+��${��&p�f��ɩ[�C���/6�B}(��<���-r �Z�Dg^��b�s}���]����c��������lU���<O�\�%�W��'{5bIqH�.lGq{�܏I��̧�jj%�C`F�#�����x�s;�P�ρH���y����&��~'3��e��IF�HfK��]X��|�k�:�@��F�����>��T�X�i�j���/o�^�4��O-Y("!��_(��(T�*���nB�UJ� �IRIf5c�A�%KjOj
iS��{�b4)���a��NʀL�*�:N~7�Z�:�t$'@�f���X�7K�[�S����_��W<���}����nu�keл7q���y��ny!c)g��2�A\g�J&3tO2��!@�^��N�<�>���
ж�o:�[
W7��S�CU�� ̪�G��E�\��O-�'�z�(}v��|BaP9+/��;�Q�;���rԝ��c��lS�Ӷ։XrF�<�Wq��i��RK?_9��A`�UL��gZ�%��֦��)	�aTCr�����_�MG��#by"�w��B��P���Թ�,�͘�^��x@msC�A�	_0��3�7~<f�W���HK0��ݲ�<���2�s6����e�Dy�e����E��eF|Z	`�)�v�6���qJ	����|��ܥ���ȺCY���䚯�nI<�2;��	���i۔`:��ɥy��ew�D�s�cpc���n	x�h�q4f�3A�V�� ����#��CHqp_CK��%�KB��,�Q�N��I� [�GMe۰b�l�M/�n�]4ź���+�aX)�R���( ��b�����8�+�D$`� Q�\�������?#��D�@[����ʻ�)l�P���J���vq�i�B7*L��d����R�F���`�&�G��.�?@��"3���G��|C���f������lY�MJ��?�W������hP�%�؄���]�E�QҲ�1�m�X�^��e=
���v�����U�`�'�t���{�<b��p��}��P>���Y � ,������.,~r��` ��m�/��d�p�S�pgF�1j}~k�3���XU�ٟ �H ��/�T�������+g��ե}!I�A�8ʗۨ�����{����`{������G������t�п���	D������[�וS���V��MjAI��+��HhK�����r[ka�gT��2@=}��a�>��Ta�ǱL>>�x(C2&A����U��<M00��ޜ���x4����:����k���C&I6��9�ybߝ�Bt��&pY}�S���-�f�/��:����ac��U�!�]k -r@n��:D$3#A��Ռ0��Xjys���|�w��ff"��I���@J��} �y�L��ni���|�;c)�B��̽��	-��w׼�$&� ?�H�� ��Q=�k����m�ݏi��K�A��4g�&Q�����M��6����~�а��[�ٵ�l�ܠ�q*vT��	�(&���<d7,z�>Ѧ;��-�=b�͓��r�k9����ö@9��VOJΌ~�9�t�񉤟	��I�{m���z`����P��Lxlu�A�Ln5APsO����� '�(� lY��O|�u�:��Hz�IMh �k �MƄd��Y4`m�fɑ�@�|$�负ԆN�S�T���cv���i	+^E�4�����;��1�	Pl� �u+���"_ \��3ʣ��ϱ�9 �mNf1h��^�nAn����摫ہ��z}=,K�ʲ���r���dr�[�h��g5�2W�0)
?q���Ѕ��)\,3H6�Gs�ۡL�(����2�X�
������b֣ѿU�w����>ԅ�np�7c�Ok=�A��k=�v,�LT%Vs��6гG��~��!�5���#�)��ւI�?y�o5�l�*$���
���#c2H�j���`T	s�X,����I��wm��gΦ��������"Q�ͩ�s�c�`�8G�B�e[b���H�Y��X#��?c��f
����ONn�. 	����L,��*#���c0�#w�d��}�X�&��A�-)~�M��bsIn��05�e�ޱM�J�{������LҒ��<����G�T��{�t�b������Qm({�n�r�y�Ǌ�_�9��@n��i0Pkئ_�����dV� *�?&>{m�0_}4X���1{G���۟��Z�~����J�T�gGX�:-��<��ÿ:l"�cKs�aH!�g
�}��k�jŉQp6��:�.&��h$$[݄�s�/��i�I�"�bR� �^;��]�OZ�	�Q������PX��6�H�av���d
��_2X� ����+���[f��b�N���M�[�4�#_8���ٕ�Q߻�,*eQ��j	%?W���UMS����=��P	��wvn�Hb���N�k�����Li	���\~����'��Ɔ`�N�k`�`^nά@���3���*;������pO�%���m`lr՝0M'֩e�4�Gf�J��9��3��C$ �fj���
�z�}��7�`���<��P8�'���9�*SQ5+Dn}�>T+�.l�x
��]���Nƻm��7�F�@E�p�	�K�1�)�~��������{�7O�|5���cm)2g��OO�kw�בE�|��b]��=�.�P,��7��*&� ���n�J�婯eq+c�?C�ۋ	 b��c}��ܯ��y��y��dIR��I���@����d���Ԃ�5�`d�V��b��k�V��E�z�e��ּ]�x<���=����J���3-�����P6=g�����=+��41)7�17}[��C�JM�
��$��R�:
��"c_*��1�y=~'V;m�H}���L��٪PyEJ��U�K={O���a�;%�n��'9�~ �m�~�.$��J�~�|�7P�P~����2�k�
~���n�!1������Ϙe�Y�����Z� ��{�E��`\�7�/c��5�25�;͇
3�˹�+�3�fq��}�%�����I�D*"sg��3ۓ�Aφk�10�}���<��C!@ Y^��Q����M o�'�.>@���Lt�O.�!J�@;�
YN�# �1�H���^�حu���v�k=��M���n�rpу,#\N�t	93Wj[�W萵��b�b��ݗ�ɤOD09�|檼ը%6�ji�O�=����u�dɗx�M\Ҹ�����P�E4���8���Q�@<y7�/�&�OX,�w@��O�zg�S��2�A�A�``��H��¦�����11S��4'��i��X�[�\öԩ��ͥGG;\noU�
0�`�}���#��{�0t/��g��P*n���F ᭘(�!4�=���b	k�k�dzU���a�L�� O뛊bnD$����rX �=�#M�YL�bgcG�Z-�n�`���`����2��_�& o);�h�q�E �{�HN&=�_t�������_���C�˿�k,E}2k��ɨ5|�.�Cf~Ac��NA��6��p��/ ��X4�����aHL��V$�W0Ƨ ��K���U�E�σ�*چ����5��:ޘ�ҿ\��4��	�+�����>-7�A	�f��2��l����V[���I�a;��D����S�kr?]\�	*��Q)S�#�m��P_lL���t�T�RR� �M�L�%3������g@�r��4ݖ�ʾQ X��2��#�v��y=f��>�&.k! G�tD�ղ�Ȅ׋��z�L�_v�����b�c8�{@E鮟������7y��9��&�W(7�' J{���~G���#�=4�2���[������/�;
�N�Q���J��̬��OY�$7��j˘3��0贳}�`I����f��A,����KY(���t M���R,8�*.��u ȅ��/�N�({��jG��m��Ѹ�}x2S�Cb��C.�oc��Mr?%����#�dkB�eKc=�+L�9� i�JDHȣo'm5��o-c��g�
��+�J��M�8O�a.��?l��<���/��W���:�e�����<�P��lsȱ���Z) �e�C��ld����T1+F��z����ϟl7T0�U���|����1���"�1+�)țm!'�?,R�Ɣi�?HB�%E�ဵ�~h���Ϝ�٪��+��O�P��H�в�x�8e
v������c�������M�hb�-����7�x�
ժI���NT�*-��p_ni�T3�����
��s�Ǒ���Iۛ�|�~�}E\7��\��.��w @B�_�ը�����h�d�+r�h����y��߂jmd�� �ag@�G�����ׂI#����o7��P=|�{�l���==���o�ٷ0Yd��^�����ADRf��	m�;3F�Lyt�n��3�(ܐ�=|�:Q��s�*dy �V�8��M�I�-w��� ��n��k)G�����B
>Lwƈ�15�6�x/4�����c$� +���	p+X�T�%c��Tq|�Џ��a�<������G~���ڒ��M5��8�:�����ˣU��x��R���HM��Z��2���GE���cR%��mO� e��*��d6w�W+3v[7��@(�;�m��\���rGo��>{�j�l	�h��<�����[�6��w�K�ơ��X����r���]r�'��R'�3��>��GM$����Ķbc)� 1�<	f�z��b]V�dZ��Q~�����z��26Н�t�^���0ہ�c�v�5eq�u ɉ��a�(w,��*Y�6|���B/tO�n�L��� D�gV�w8�&�������K@GL������p.��ʞJ:!��a�X��#��
��*�ɏ��rla=����D�?+{����M�oh�H��	H1P,w�2ӟW�;]sX��5تO\R�9��|z�0P����������Bb�����O��T5]��0�J�vݓ��"��;���E��nޮ��5Շ�9:/�{Ӷl��p��9e�"KF�����GBO����;LC�ij�?<ˇ�oe|�Y{=.����G(�-�ـW|�����Y�4	)����G]/����ֆK�X��QO�+	e�ˍ����wD"쑦P��w���7Vz1e����A~����í�?o�l�0�E������F�6f����5��?i�F�\�+������ ��f\�')�"U�e����'��uI�"�͔��T<����/=%����'�O���m��葆�XҀ� ��@����1`6�@��l+w��m�z&��X�A�b	|:F�D��V�)Z�׮�$7�V���6����~���>9�{��5�c$�k[CVx�nf�-&Rz�%��n��Fɉ��<�s�������R�I@��*��l���[.X���8M�FX�D�n��KK?n�-h��7�1*d����I�,z"����ω��|��Ű���t vA�����,1g��/���V�9�t<~Qύ^�|9��..�<?��O�!�r2G~�P4���D���˵�O۳|`߹�X�o�}٩��z؆�����_1f�I��WS}���֢m��_]߻�ڦw���/�A�p���,���#/k-�v���g�G��bp{Y���'�tR<ify+���16���k�tJ1�f�H�<��b���}���HN��E�c�D��ܒh�jg�$����4�]�Ok�����V�]m���P{�S8l�h�� ��MCy�@��=�Uw���c�g%5R��n��K��ܽd�1��m9!ŘC�y���LSge`�r�b�)��,���)_���B�`����^#K�g�G�?�	��&�<��m8�����;�S=6ſ�b�1|����o�0z
+�0絭h>_�}�fT=Ty�Oa�?c|T��u��)=7"tg�����j�G 8|x��'}n��3g��̃��t#ԍ���L��
Y��Fyx%(=���g��<	��.���n�5C�Y���j�I�����7u-��^(���H��~m����>.99v��@��p��b���40�Azn!M� ���ߟEˁ�N����;{O��k���������R����Y*?��ٳ��b�ϟ�bG�38j31�e\.�&�su�������>���-/*��|�x����=�D���<�Q�� pАok��a�}'l�������5�.V�VPi�]��&1��	�
6=�Ć�f-���?pIR�L�vA�L�=��+�>�9���w���X	��7q++�LP���#�^�zA�L�ⱥ� IY����1"ݑA��PQ^��Ї�P����&�5'dz����8̌�%`����L�X��~��$���w�d+]�| �����dT�ǹ,m9h�K�3g�㎥<+��s��f��a�,P��ɽ���8`������L�
d䝎w�Sj�Ռ��A$�`��Ⱦ�nbTY5��_�Y���jm:�ae!:��I���(�_�ݘ��V�����`�V&^�������q��X3e��o��lJ�l�[m!�ף���>�\���
���r��M%&��'��X������3�[�:�������ἢ�Hz��T�`�yyy����n����W�\��{��
sb��|���l�P�-��a�Ԕ���"͠�k�5v������?�����/�������l�Ĥ���Q��%K4π�m�@����W�_�Ch�SP��k�6��)�v�x����qo�>�x?j6j�Bq�7X�{�S8�5�� ����4��^��c�P�mw�|�,�� -�{��FK<�B�hi�xh�2 �X����C�Y���#6���k�)���x���/��5j�Yg�:|rN�\�4%���V"J��>�g��z�i�=�`C�&��^{���F\�� h��:y���w�!��;)p�O����	�H5;hs�*(zT����R���5%��.���e��ʺ��<E��ʢ_����������������������h�!^&�*�H���Eo�&�� �WJ霅��u@��H�J	�-�>��<�u<8l�?�m�	X2vf�a˝p*(��t�V�������o�MCɢ��ϴ��g"4P�ӬOHkE�<���ұ�a1�J
-�b����`�H2�s�\��%�J6�J1��V�����b��ƌ�8�=�&7�#���NN���o>Ɂ/�(r�Gн4��G�}�ԺXl#dn ��}ϹB��,z((V�([��ٛ�B��W}|�a�!\�r�� �ǃ^�Ƚ���n��al�������	���͟���KL�����|�&s%�a7җw97�HL�nYP�=�n�s���@���0-ө���i��\
n
?�<b�<h�O�����X�(�Jf�u�rxW� �S��{*u#-=�H��A�C/���ƊP�����>$L���*�X_5�3�naJl��� �t���q� ��H���i@ ��S������[�F�Y����	3��%��=��+������1�F�����Y�d�
����ev��?�g���"
�Br�*����>kl�Zv�E
��Gism)��>���N|��[-j�TW<>#2���|TA�|� �>����(�ۗ�<�xj!jI �� av�kH�
���"�d�b���J����C�}�9\�/D���E&;�L�2a$#nss+÷zΰ���U�,w��Z��Z)Å$�N���U4
J��K\sPK06Q�n�yOuʲ�!�x��Y}#P傶�|�ɉ2�;��o�g�S_���,XB�jqt`]$T�̻H�����XL��,�,�?��N�z�����E��{��au�]�=T?�\��f���/�?�᏶��y���
7r"�?�ʚjh�N�F���Պ\&�ڊ�sb�LØ�WLP��͖�[��b�se�������)a��`�Tg��A����r���"��:�]g������L���Y�����g�ڋ�����e&;5H�x���P��ˠx��#Y��?�����&�c�7��9��ho�C�2�평�N�jԏS9�v�����y�P��Z*���Vc�b�(a�9K���"$
�t$s-�:��Em���XQ�G�i�-�ǝ[��;�a���#.sB%b�i�i=�&@3�Ҝ�e�~Uf���Gc���J=�j��,���_X�Lu:���ҷ��
��ɀ
��~��H�U��*�Y%�����G�4)�Ȅ�����"a��O �i�e����;?1����.�u@�k��ו�рX�#���+Y��h�j-�(��������Q �/�9ُ0l�V�������B��e�ڹI�mMD���Zk��Vb�NC(�F�Ő)a��5Lv]�#S�Q��v���Vr_���������K[�g�2��ҷ��[]|Ǆ!^z\_��%S��G����E���EM���6�+ە�N�0)N/v�'�1Iu<�2��W�E��)�X����f�>=d���~�� �2�����Y�������fj�ځD�KF��H���.q���H�nL
*����Z���K��N����Fو)���60^�3�/0����{������"j[H�&
��:t�β�Xĵ{^S�F�����ܛ��9���z묿�U`��A`ŋ���^I&@׌K�x��p�� ��	M�c��	���JX-<£)�P�(�)��>%�UL?��{s��J:����'J�@?/�U;����a�Bs�2��f��:��^��+�E��T5��ӧO2�7��7t�j��p�ڟ�\`��h�א-~��u|��������RI�O5�Lw�ٛ��-���EV�w�
���=��Kǻ0Tf�8�����l�4�a��gڞ~�$����Y
����';;�0m��g'���*�kW�q�O��KT��Ύ���T���PsSB6���_��Cks��~SS��}A�%�p!�ـ�������Y���G��c�䯗��#.�\ѻYP�v� E�BPY<��7����+a_�Z�������� r�C�Q/��TTƜ��n�Wg�B�&�`s��P�W�J��<_����zTf���6P���vj]�Ӓl���J?�~���|��,&�4(_T��ȱ�(����L�O'��*ok_��K����-��*�i̇0�����>����m };E�?rR웯�������$�4��t7�"�����Cү��$8/fAw&��*��g�==��a\�����qH)|<,�4�&�%5r+Qwp�,�5�Vtbm�I������,�\I��Ԣ �$�n0�e@+͚����.߇z��0Ϭ����ϻa��u��F#H%ްs����w�F�߭T~����B�X^amK�i�@60q�nZ���2�9�- �m��Nm��*���	�ԊѾ��o�����}�HW�l��'���f�`�ʻw��M�0�y2 ɍ6ިYa�H`�{�	�9ج�����;5��濥.%M�¹��M��I�[
*̟�6����M��=�����o�%Y��K����}_��y�,�|�Ym� ��1(�L�'�nsX �	,1�\�"�u�q�O&�{��e.S�K_�V�[�?�w�rr5�c���Ԙ��~˷�E��R��5>�x8�z��r�g=c��3��|�c�drHK����z/L��2�q�rG4O��pG�Iz�m��W��٘63N��N����ⴉ�� �������� �Nڋ�&�{|�,�Dݿ�:����YiDn#
�b>T]Ǐ-_�����-}�>�X�7ط(�ob�wJ����e�\S��(S�i㲒�)�"o�9N��ǻ��F]��h�F��/R�� &���䠬V�L���3���~�3����ڣ�vg�zS�F�d�,y�=�	����b�t�#�����_����L���$���V�PJY�(08�X�_\
D,��:��ϺI�����?#dL`�I�U����������X� yv^f�������l�U���R��x�?)�Ɂ�d&��ZN�4�;��9�i���vD�g��M҅�f�J8�޴���yO�7ah��{,�j|�!�u����kQ1��1����d��mS��j�a!�3��Te�����s�%Q� �f�L2V���L1��s_9��S��xC�S�|���c�����]L~;H�Wy͠�C��|0K\g%gߩ$��$��}�� 	�˯��mN�,��)��r�"�#*��΅0��o�&��GlY����M��w�d�׎oQ���]�o{�L��kW�X$�w��O�n��E�ۈ5-B@\o ���.?gvg`z�P���^W�^E��$� �	D���tz|Q����C��1J�%�{��)��5ƈ��a��	h��nsX�T������zNB�T���tA� ��������[�7��̉����g���`�}/ ��ߛ�#��s��"�l�.��	hM`�� �_��A�,v�E+���PK��% ����.�&Y��N��|6+�/�1��òM�/3(b��8cP�	���}d��P�9p�G�����e~��-�n��",�A��۰���A9%aX�ܘ�� �~'Zv����<��=�K'Zkg��=P����)��215�`��x�j9��n��>?[T�� H
,=�m�.]X��.�[�6�epBV& ms��_]o��6���;(
2�J�:�)�Y|�n��wZά4'��3uޘ��e�{w�`Zg���\�%}_���<�N�|YJK����<zF� 4r��3��ݝ����A]�=ǺG�W��������w��廉'o0@����'Gyz�,S��'��F(X2D�ݶ�C]�-��)[߼�O����� ���O�=�x�-P�}���� �](3MS��Iӷ�$�fj�+���ٖ�-Lt�.��TW���Tm`�< (�7��%m�aY*�(��M��v��٨f�Ζ©�|Q�_�dtP��-�U{�N;o"S�&R,`HP ��ūz��P���b�(9�d/���k��14o*��Y�K��1R���5=�D%'M�49�'Ӊ��rjKN��$R�7�h� 1��t~ �V�Н�Zm8ϰO��c&(�N��o�)�`�gj/�?kz�|'���؂>TG��c�B̎T4�?�R*q��v�>��P�n�Q�=��Q�&�Z>��4�D��i`���r�R�^h�t4�2�,���d��/�D�]��%����o�S�ޏ�����S� ���������ݳJYr�[2��]��1֔�hǻ8胈$�=��L�@���鍲K���Z.�k�|���ȷ�@Ւ0E�{�,䙖l����k� ;�2w}E��-^?����)
0���WK4�5|��,m�r{�9f�2<m�냶��Wxz�4���U��daV���I���s�[������y� ��v�
���C~��g���_n�_3s��njh�[jG�,�J+9&�E;��0m$��]��d�&y�j2�R;��!g0,6m������.�ůͽ�z)@�wh����m���Z;5<�x�6�-��k�����v���d�N�������~�w�m�^���)��,{�1{a���-H
Z6��պ|L�B���>Y�J�0�g�bܽ]���A��9�"9���L-�~/�lsV��N"C���xBj��#<gT���"~bɀ�
�9�U�8��?P�d(6�!�2 ��su+?����o	l�M*3���m��
\�\ƒ��^�.n�	mf_g%BbdR�(�x2�����e��Q+��ӯ��*��~>�|����]߯ϵD�1a$)��;
��e�H^����R��s
��-:�e��Fd"��I~�Z�ҏ�^�z����x�O�~!A?��5�f��|;�0�����i���ѥ6ak� "L����A���M ��&S60������ngL"XH]�-A:['�J�4�E�ҷ��2����z"3-����-G�o�nN�?bc�މ���6dR���9���ۜ�n7�X�r52�m;hݤ�����2����i�r�9{?�(��$�Q_o�P�en"�<i_��,d����A��K��})�-`_�c<&�?��O�lþ��I.�ob��u������9���6������ �i�Q�����T��)�Οl1�$vg�ήS��l{��x����@уX�	���2�{��э�J.;��n�i]�:3�kU�מ�$�	?T�@��!��{�UE#���B��7j0���:�~==�ܦS3�(<�� =��o�GQ	���i�6�Q�Oi���|G٩Y+�>IMOU(=��w7$in�Ʀ���5�&��yޞ"#=v�[�:Aig��e�-�v�G~�0c�����-��=�_��OrV\<u��8��k \/���3�������Tn�]�۞�X�rV�q��͖��5 �T"�+,�K��k4.'�-����@�o��el=�����WVɆ-���ҒӼ�b�ǆM�1�n����ۜ�x�q ��mo���&�[l0�l�-�W��Ү���Á��v�߃��:E���б얉X���ڴ�r���ۄ:�C�V�Zl	r�,�P����P�q:N��O�jq���dy��y"��`.2K# �9�xH_��E�!�G��:o�{"%[2��LK#�rumn�MJ̶��^t�V%����R]<�C}�d�KO��p!��#�b�u$c�F��ʟ-X�����]>	�}�-@�.R�M_#��
�K���)�v���P�)��K�R
 ��ԨM�i'���Y��k����Ï?�>0f6���N'�eN�V��^��ַ�>7��Lz�lR����b��l/�r3q�
�tp�391�P�X���_�7]�Cgj�!<��6�;\����6o�6���)і	��H���wAMfv=r��xiZl���Ep��a��-m��8�y�ة�Mm��]�ιJl2��`A���sX/���l�u��P��I��")3�#��&}���F��c>?��C�"�p�e��Ω+�� }�}����m|��֜��1b��]c�����t�������Lh&yI�/E�촱���$�2�d��jO�1*ы4�%#�c솀�G�����q�x���
|<.ub#7^cߐs3^�}�"��r  ��mވ�����L�덥�fd�?��lG�`8Oi����C�|@���[�g��1N�����"KP����#ho#�Kg�{C�U�wO�6|�zs�V�P>ͬk��". a�{�����}���q�,^c�U'����(��ۺO����b�W��V�F��@�>h���K0qc/��Զw������hZ�I˗�%+ꦼ"��,Y�T]��Ii��z�O�_��0�5�H��H�/=�7�kYO ڶѿ�W*�:�"�>a֧"⢂�r�� �
Y�����yA�v����ˬ_�ge�C����q����W��߾v`��)v�	���3��>�`�n�������Ϋ����g
�Y�b4�p҉�����e������!����=���k2��~o�&:]�hhO΢u��{21����Z��AZ�P��'3�} 7�����ox'��Z���_���ɖ�5׉�ushm�훼��r�2���ɮ������ ���O[S�r�N������HR���s��۶ |8b�����!0d�����=��r��6B�ox*���BP��3���-���$Euqߜ�H&Y�ET|�S_/?�.�sn�����=?��E�h��]����\�R�ۅIR�:��,$�p�ڲ:=�/�_r���t~���Br֨g7�ⅽ�r��Z���2)4g���1�{�K��ߐ[�60T��܈����M�v��S0��?�AxfWcZ���`�f3�b�]ˣ�tD�5�<��V��%ƚ~2�b�I4���Ckx0��&�v��D{i[�!+�^�v��5�
P� ��걟-�qa5D���5�����P�#�LUɘ_(�ُ�c$�t�b�&��6��,&��R�x�{��J~�|PJpo|����ܶ����q���9<&$\Z�6�+���������W���#�]"�6��2LOv$�?}������=&&��gR �vODHM?��7*�%.�g3�u��3�}��!w��=�/1C���F~m���EJD\$�4�w�Y�;A&㙕�3��������`�W2cq�$ޣ6�O �k�xO�"�xR	�o�h�э<8-����̔�hSh���.zJpԨ������zZ�6�}��V³<a�k<,��]� n�}��de����� %�	>�� �+�	]�W��[]�L{�$+�.;,�+kD�f���5TNj���w��o�`P�E��[�8z~~��u2�Q�c u��(�N����!��¨���Ev��0�K9�}�P�j�`�M��R�~�Q y���L���5����_��gf{��|��n�z��q������RJG$�T�W��@���~?������pU����tL]u�	-��Dyz��{��\-�,_�|P�+	$�1�UϜ�[�_��/qyA;9xG�V���4���W;&q ;l�16=o����4��b��Zb�'Fm+�����e�~�v���s�_�j)8���S&{֍M��j~f)Lf�UXIާ�,ZȻ.�e��Ɵbyj�v�Յ!���<���n���Y~���w*��X��|�z0��Ӊ�\s����?ޮ?|@��(z?�'���|G����'�Zjݯ�E��GF;p�j�x�va��k���et���A��p�q����}���f텕O�{�[^vg@�%�Ĺ�������~�*�>~4�v�^�}N`/^X������pSD�>��|f�?�S����	��{�����M�cf�!3/�/7`�l�g?ŒDw��i�8�n�����r~���ϯQ�٥37]����X.9+�j(/���*ps����A�5"�r��Ty�$)���m���)��Y!(6΍��e��ݴ�k2�d��#�>:�P��=F,Z�k3ޗ�FFz|�U���Y��AZŰԫyX
��ZP���~�����Ab�)���w�����7GY����su0������	���o�e:����ӧF�,�# ��dn�|}}- ���MaX��f�0����"$�.eM����"(K���Lz���N���V�+����q���>�"D.av�8��a����f���O�b�33oS�[�x>M��r�����(�_Uu�2۠%wX�H0��xy9ne�怷�_d��\ ������1�j%�w����v�E-W�7o����ٶ4�>���.;�~P��������/�����)���7 K(]$I)e9����l�����J�$��b��)�4f�W�e�[(���/n���Ė-�^`��ճ�[~uW8i���@]_VY�v<P������M�iyhC��Y˦)�j�
�'ty]%�)�a�Aq�����\kv� >���=Y+]H���zl0G�R�6q��*c0G�>/�gω�.3�'H���|?XZ��! ���䰜4ۍL�kG�X
-�7����?�=���+���f���؞I1<�!�	�Hs�w�-�ݞ=��H�($��*�,�ʘ�͎r�[c &��{\�\�	%lq'@�G�'��M� X�R�빏?� �˟����[����2��V<_���i �d�d�Pg0m�l��O��3���e��߷�*9� .��n���ܑ �D�E!e���p�xĽܟ��^oZ"t<4۔�6sxG�MF|=l�@�?��Ҡ��'�����QW[������A�N0,���Y��ߡd����a�ϙZ� �-�}�?�|Ѕ��E��9�U`�.�|�V7թ]#��|�b����L~��G`�kL���.(�(f2�

'� ӋL��L-d��%}�sj�su���{� ['���ʜ�]@�cf��-�|: ���7M�	�fj��:/�A���b2�wm\��m��Y���]�}��2|����\���"0?��,��.j�z�{���N������^�q��Ly�왏����u`��o���ӧO��.������ARP_˨�o}�g���R���>�x�]OG	����;ף��]$��q��k��P�;ԇ�/����!��L��Mɡ8��N���!R&�?�|�2���ό������ߙ��F렀�"�ھ�K�Oa����zY�A)oY.�Қ�kk�Nq�`I&�?��r��՟ح��O�)�<|��j>+�&���,���U��%&&����%u]��[ ]$J�m5dcXa��o����"�@M�D���@*'V.M
aBJ�<Uw��H�!F�\�x�+E]0��C �͑�.r���<� 0^�j)�2���+�>�eda
t���잫��R���Q6m�	P[�T���Rx]�a���nz�Z��� ���zcC�&@=�n/��8�l�e����(@U����>|�魁���?f�bU�ޓ��&b���O�ی1oS�����.-�����	�b�D[�:m
��m��M��7�`O�.mK�<�J�a �����`'�F�>�=�����d��5�"\
}
�>�&�~ʃދ	DǣRu$�4�/��5?��G(����6MX�m�v4[4�Ҭ+��:.2L�=b�`e���Ƣ.����pLn�WP$����m|�؂��������������B��ax�3E��)W��,�,:�x�L��
���_��oa��\�; �іקk�M ,�����_q<v��/�r����
e�G����i2_����`>�£��㊀_͡X��ͽ�N]>�we�4
��h��ta�e��i8��C���	�X@>���	�m$@^CȲ���� �W������ �F2�Ƭ�f��l3C��l�Y�/�E�B̞��q$�Pn��z��i�N3�)Gcfj� �k�=+��~����ܽg��F�-\� 9A��׻���x���zoڵ-+It��p��Ar<���h8$4:�>��e~.s��yPY`�����d�������(돺��ct����n���q�_]��Lm�SZ](�W$�#�K�L���޷=�O>�CZ<�7�|����#�D7Z^�,�3�B�W �����`�� ��gÌ�kh�m	���q<]�)a����X�F>���p8��o0�m� �1���X�y���G٬<���&�0ܚh��$��������H+fg 1Y�p�Q�=�����l����ͪVpm����	���sr�D���DT a� ������
Pm �XЙ���x�{��@�ʰHC7x�ͩ��-��<���y�vJ����x�s�ٍ?r_���<N�]��-�G�Wtc�l#�,W��q�{
��{,/61��m�A�D���/�� id�ϛ����jVi�N��> �@t�oҔg�����8)��(���1�+���zg�
5MÁ@�I�77$������~��ɌR8`��0I��S�͘`��N�b\���&���kw���$םf�D1�7��3ʜۤT ��PQ�8��N0�e��`W!�/ �*�%5�9�c�bRc���֮V`3�4����-`�G���Q�%3-V�稳�үݒ5�~���ɋ�Z�����p0ө�T��%���!p�a��@���9iÕHK_�k7��X;�槊�H-�槚���o�/�`����X��M����J�6��  �E�-l�
�
Ⱥ�H|R��9�-u�����l����ø��P��k7;�K�o�O�f�$ui[|�~"ڎ��h�vH�ҀQI�nqI��k˜	_	Q�c��$�@�'�aă�K<�1W[Pj�*\mT����"l��ȝ�Ӝ�3����6ǚ<�[{G�k4[�*(��B�7�C��4��"q��%��0� k>�<��h��q=�?����c�at��f�N�IeQ(��Ĳu�'V��-�1�=׍�{T,��_�(B·'+��SU��sAp{X�]fC ��J��`���8n$��a �k�����Rv5�6�C���A����>g0�5���;a�07F�$V�Z}ײ�:��CuT
��T�_Ir���9Q�,g���&�$�c]I=XO5� ���J��O�CŢw�O��OU�zA��,����9�m�gg��.��ґ7�K�|��'qƿɞ�[�.�����t��@O���Zw��o1��,�a_j�2_qs����L� $aj���{r����0���.m��x�k�z)�q\�4 Xy���n�:D���Е���;��Wu1��
z2uR
F�qǳ��#��"��]��c����� �F�I)xF�֜�KiPYg]��/XI:�I`@]2g� ��Z���ޖ����+��z��zLm�o��5qP��+�滑=C^[!!���`骔�w���PXH����:V��;��qV ՟d��X��늡��J �_�"��+�f�8AA�f`�j�%�Wv��d$�Rl�B�v�٣Ǣ��;��"?�@WZ������*�@Kh���������S��y;�.���&����0%*��:��>�~�)�zѵ� �z?�'���z�؃����)�IZV�C��i��ֹ��<G�C�⤌���7>?٠�8zQ�i����)�k�xt�A�Y?�ǌ��?V��"�/zs�������T7MH�ϴ>PӼPE'�@��9Wp�<�b�C��理�y�<��$��}��5�$�ZǓ�P��Hҡ�+*�NV�g=1�DEˮ��)���a�ѩܻ�j6w�FC�ʍ�H�=�����Ħ��i���Y��I�4}���C�G�дv_KX��t���M�H�\)�	؉�)�#ё�,����zI�Y�V阘�F��EC׆тfb�(X�l��/sc��zCaz]֣�>�`t�H/g9W�;!:�%�Z5�Y��X������ꂲ�`i2��_�R<24fU$zoV��p8Ж�����'���֭o6�\�+MT� w����8��ã���XEu�F�E��R;ߠC�w��3Q *P�t�u>�e�x�s11T;0�[�Թ�㑠~X�Ծi:�C�v�=���O9).L�3��������A�K��]�o���&��>&P #����>�t���ضu)+Q/S���1��Q�Xr+�]�2�j̍��Z�b�?n^z�"��h��D���-D���3%R�aqw��FH�]� U>���z���0�K�)�	H�>�?�{�.8?9#���=�����R��5[څ���$�6�܋��!�y��o���!x�j��9��|H�-�,RB��v~d��~�[X�#136w"p|J(�ٸ@$PK
��~c�E�Z�M���x>�2�~>ᚥ��5㋶�E������u��rDK#� �mǙA����X��=��u-^a��bQ����VNa(�/Ʃ���"�݌S-� �b��L�?5'�>�uuC����/����%�lt��9;���?�z�d�	U0=X�+&Ʃ�����?��d���]�] I���/�k�3a�fK��l!!:�;�i�?�ĸ{�>��Bd֏"�/���u�J0Sb����"=Ug�
��z �Js5R�YUOj�9ct*Bvc
����Ƴ�i�۵{�х4@���Pq��h������ZҬ`E����W��U.y+�U�1� &�?�Iن�Ap6V�5Gvv|G$��X�h���U#ł�#�$K(�����U(N<����Y�Y�:����A�$�SjQ`���qo��0b�*�Mޯ�Әd��D��R�O{�?r<����O��}�C�R�	�� `W��u!���s{�w�����ҹ>�D�33��h�f�jb��=��'�+�C�s���%���	b	?"��c�ú}N)��"�E^���G�ᶂ�ԓ���IQ @�� �_D}�n���y�J+��d'{¢��k���hѕ��{��b\٘�d 
k?Q0�<�zPΞ������d�Z��%g0��@�i�Du�B���e�%"V�p`�=����6R1nR6�$&��B~���iu8�����N�cC��s��h��9M��g��{�ܦ�����H���4�£?���}�� �I�x��Q�� ����'%5ା��	�hq��be�����"�~���X���Y֍J�b����rm+��EL�P����Ը��C1)a��Ϻ�'R5A! �&/XI���EX���E�p#2�X`,Ib\bɞ�luOe-����i!:��t�K>#B�s�Ƈ�˳%�R])��b��k����0¯�Ũ��+��p���T��4����U��{�����u1����w���W�䱾���V�SW-�����y!K+�����g�	"0��L��'>�C� �T�@�%�{2	�5��1/�r�Dp��K���� �t�>���h��!\����ښJ=�>B�J&� �U=�de�Ln������,�NZ��%6WA}\s��	��C��U�R�7i�����i����ˇ�Ws)h�^�|��秤�}��s*�fV@���ռfp�����B$q�~2�1gρi>7��i����`�>�	��f/� !�5���d��i�+j��x�BlK,!���~�Im��ζf.�|o�
;"��_%-7}�8;��U.L!([ �T'�����&�����8dMW�b�U����8�R���<mp	h�Y�����!��,i��v����kx9�$��OnM��1(>2�{�����J�u��2��S��p���9WE�:�`��|<c~m�Ε�L�=���uS{��[�����W��睼��yG��΀���������'�F��N�4�eLpוs�§���v����䀊��u]Q����C�u:��.�X��,.>�H�K�Ɏ���k�|d�}�.�(���xY'��?s��s/X���=�&n=vF�Yl���`���!~?w\����@/��F6(0�������%bi�8��}�����p�EgK_`d��w6M�����T6���Ikn�G�')����ף�n	�����i;��&�zr����F���U�-p�S��'��� K�GY�Q�R�^�8y>�^}?w�@\>���� A��o��@�<�����Tj@��ɮ��ȯ~_��1�S�<+��KF�0̈�`���
���ݡ�������i��=.V��#�Ùa�uTCĊ�e`l�Y�X��a��9�Ԧ�2�˓�A5OȒ��	�-_3��n�؊��^QT9��z!e��Y_�[�X%�=bsЗ�(\�F�P�����_^g	�}x>��Xm�]��@)�=I4��y�5�Z ���:��f�j�hh�{g ʕ<��Ͽa	�����-���P�S�2t҅~:sLu����÷�&o|�m�ŹV���6��j*]�B�>c1@��v#��%��!�̇A��~��$��q�P�g�Z�I/7�$�oov.���g�Y�Wi�|������n�W+Q��#L�`���"4Ry�D}�#%��=��t�x�>��2Eǆ*
DBP�8����6r�,QE��g93�&kvĞ}��:�,�����QA�ޑ͘�Ԛ���B��ԧi/H��S�i���ς�mXH�c�/E!)�!���b�:�����B�Z����i)�4я�6�DL��i�\)uJ������
T�{� � ���2I#�XM�����x��� �Uu�2&�aT�5��Nl�4`eQ�'�*�N����"���NI ���ꬉ��ᥞ���ک!~���-gT��
�KY��. �ޑ��G�9~P��p�j&.���k�S@(9䷴ W�����
B�'9F����d����J�*��?l �`��'9��x�͐�,���V�����u}��[��!5߭䈾g�x��g�+6���)�ˆ�)�G�{X�EG��k@��O�j8�>[��z��n�E2em[�<0耑�'�څ��X�'�������4e;�	��XtJ�v���}S���u\W�'�V&b�:��L�=[�,)� �gq��/KU����H�%� ��>�%���B��+e�������tk��}����|D�A߆8s~S�2�;@(+�]�/J���DQW5wm��rw'w5M�[��:�=���U���
�hub|�%X(��`���X���8\X�v��R�t��Z%��N�g-�3��i�A�}?A�<�$�Q �)9"ɧn���h�h�^�0ɸ�F��ū�$��g ���7OO|bٙ���D���Lі�B�Z�ɛ���,��W���ՊřGٔg��R�$n9E��#�.(��˺I,��yn
�z�m�g(eN�k�4|~�c��gu�2�&�;�[�oXP9�R,�}� nB$��Y�oO�Uҕ�Euf�W�nJ��üYte���B�M�:oO�A6'�K��k��=0$<�<�*�0�ƛ������J
�-�9�����ՐB��A
�I��)l��.DPlH5��\��6D;<�R�v�?t����5�<��h���.
�|���������Ȕ?}@��XCh��E2iO
�9SO>�t��8��6E�̡&����Z�]c�9�T��0 8��Q�Ĵ$�9Y��7��vf 
 y>DdG�t�#��3��"kӲ�?��0���R,֤x�k �7��0���3۬�P��h��JHzQV�I ��p�g�2S���1�O�i5�OI-��Pd�j#���.�T;e�RW�x�lM1���:s�bB��6�xjY��sd�b}Lih��� 
�hPa5�b���-u��:	 j m��?'�&���	�pԬ��y��rT�|D�="�)���Xڠq���8��kU��~�������]���\*����N�\╕��$�
�C��c]c�E�j�w��3�߶ ��關u�Ǧ��.����b�d����m��`C���|��Z!I6�/��ވ�lՄ�`T�V�d�*�����O��2��&�4apq�����{h���H�W(>1nS� _Y��	�?H?�\�V��܄������Ϥ����X���tgo[d�y	h�S@��nc���9��R��n˕,SXuP��Ml�'O��3�O����,�V�E+ �x��^�xIϞ=�g�'1��n�}�Jz鰹��:ҧ:Ч��{6�6!�X6������:��s&�zUu.������Z��p��ݤZ0���.�sD
#�7�/媞��eT^�=�3�����ҝ������ș٩����'��}�;݊��p���kB!3�-H�*f�\x��E���H�b�Zwj�{XY֣�t�iQ#uZ�.H5@3\�lx��d���g�{�_���a���b���(0'j��M�����-^[�'���AI-��j�(�j�H���bN�q8�%kް1OLY��bg�ϑ�i����"%�9\DR��p��"'�P�7@�|Vm����W��A)I���V�|������*60U5����W��j0�2y�d���u��2VشJ���cŃ����/#��6���nQ͢�@��\ֺ����C]c|�MŲ�|$�,V6 (�}8�'�8b�)�2�{d_�:��܄8y+q̓�~�@�u��q�<iv�L:�y]�C��.}TLWfI!����=�ٳ!��%[{�ۖ�7�� �.l���E���A�G�&`����.p��Dy,L�#���k�׻�N�j�n�4ۅ��\��Xf�mtk�z��d�>���5�t��B�6�m�%]vK:I��#_O1'�b���
Qܲ<��\�0���B݂��dL����V����I�;���߃�))��1��G2.�^�&�й�p^
�&���
��n�Y�R���]�!�M���_c����5�'֡��"KSY\E;ec���]ۆ��-��F%�XT�ŇE7�J��'� z���3�L�Ѓ����4I�pd0]��ho����%[�$	��3�EȮ��#�M�"c�3S��$c(�i;6{��,�����`Z�I�.=���نl�L�g�*
����TUY�����$R����K���TQ��LQ�"�&n�ʘ9��h���������<�)��������Tf��C<���G��DY�#m���@��\�ҭ�qZ�U���F1�E{Lݬ֨��2�M�<�:k����� �w��3��$�fn�]]�b��V�p�<5Xm�l�5�'�6�	Q�0��:@aP�OYLlb��
ȁ�&@��BXJ��:�2���w
���K}õ�O"������~��=��R׸O�](����V�Qt�ƨ����=`	�N�p1O>���l5� �˝[��I}����	���d�H���`0F}t7:��댈ն�9k2u����j�����4u0��Q��G��ȯ@�F28ro���ˬ�*������]HL,ʓ͢n5�PҚ]�p2�1� ���Y��@3�J� ���#:P�	��/{ɻ���Ztp&$G\;�\T��j���s��,��f�5���/�����
��4)|Mx������O�C5�oB�b��wZ��_&׀��[&[-�ң��X�^� &����,���$b���zFta���u ��Pu@�=e�����|�xAo��:?f0��3t�E�����K�:g���Xl� ��YDg����)L���^�Hs��-�ˌa.:�H��z8��Vl20��j�j�,�qvp%?ޔb�j5�sϭL�Gu�i���6[$S>J)���KaH�}~uT0bf~�����bLB͔tq�� )��6S�z9��(�U�n��ʂF()�@r��ڮ���З $n	�)�vA�����l?2k���;�:��liʳY�����A�綳�c�TH|��1CTv�J��HHt��	E��>�>��ɻ��gN�,�rˎ��(և����iG�2����y���Dq��ҧ���b��?2��\Z�\�OU��:�R�i��j�n�Ӽ�L&�ju3����X��$u�>�`e��!���[S��;6,�c�B�:N���nS-0�t�L��3� ��d�~ϋ�5K\B%0zP�نd�# @�I��E�9S�4곗-�ʙ\�4�Ҩ��Q�( ���`)����A�
���,Ku�&r.��Ȃ��  �vS�X�|����z�5�=��A�E����:��\΋�_#�]໗�@֝����)n��%j�;�(�X�|��`�sM:�kq�'s��p��ź�e�eFԷ�j�1oTg�O���V5�>���	!TT
�2�'C/��˻֥�~|z�0??��1��5��A�������Jiz���[� ��wZ�n��1Ƃ6��"�Z�u<nnvt�ۺ���y{�}��="O��������J��h&$����h�ju"W��J�0����ʶ�OK�16D,��#�R�c[zh�L;ϕ-ϕ���@�����!�+�/���O6*�N�Dh0a��c�Xך)F@@�$c����R���'�rMXUmЛz�" �\��<� �m�b�4	`���{;�j�}��͟g����+D���_����E�������a���AL�E��z�ֺT~v��5Z2�T�#ܹ!;.`N#��L���|��k�|��a�ј�sc傭�P����:3���� R<�,�,��uH���Z9�a� u��Z��o�F^3q4���GE�I@��>����H�E�&D%!�td|¹���3-#b����c����7 <��p`oD����Xd����g����>Gˀ��I>��K����nS^���!?c�;�ͬ嶇hu�̶ �_�������7�y~OϞ?���s��̆:�73�G�Ry�Q�C~����	����v!�7�zӕ��a�Sr��`
��5�'w���P<�-
.���}�-��M�	S���% `K%����Ui�&���@�LU���`�5�{5��~�^�C�P`d�"}��	�Q��F/�=\����,��X-�US������Q�;䡸����e��.��`l~����V{�bඁ�FS�F5�)�7�7��u�R$ON������\��Hn�Ɵ.�;��I���؞�*͋��u��U@�{��Y��r��PE�g@��O�?��g�R7+IrT#,�����[�[��E� ��:���N�*�`�q<~�`��?�E�/���2�p��Ct�Yep"����PY&���k�X�g��@Tc�����3a��ذ�o���4~��0Z]l��_�t�� ͪ�h�$��Y���dB�KX�����	�ʋ�q�OϓE���Y0]o��snl'�_v���;")��d*��o���+:�!ΛP���U���mߨ^ja��������	]�����~Ɂ}5Yݰ+l���~�B/���u�a��J��~p�KL�0�@���� �X�ӹ��@����`�E�65���IJjj_m4�]�ޛi+��ס�`����nׇTy�H��Tc��˳r�_fG<n�'��ғә6A�i2^���s{�G�@�)�������?�����_�Ub9<��x���^g�	�3�G��Z��y���;�9�0��2�oL���t�s`몏�Z�qp�ٹ��7����ryy�	F�Y*D`��W��nF�y�M$�jނ�lu����k0��9\{L�?{F?<!N�3H� ��(2�YD�	�oŀbu+:V��y��D��7����y��F~�G54��'� �7�n.�d�e�g�YU��c��471t��u��`qxw������}�糓���2ag^�6�2��\���f{�Ev2]�9���~�z�)��[��
3ݙsx���Le�Gug�m�wwN
��Vwi#3c�:?�n"��9K<No߾�òq������b-��ۚ�¯�ڝ����7:���f�-� TW��|�׉lVI�~���J���S��0\���8�F)�\�)3����t��gB����rQR�T���?M�E�d����9d\�A���͎��z�90B !�=y�e1�u_7l����
�b{NR�; �@MQP(���N�Ɩ��7�5W���S,|R�� �E���ea2���je ��$��f4$cj,�N�ɢ�\�nv<�XT��{r{�V˞�!`J<)��C��yب�"����~E���&h���Ƭ� B-e� {�ۘW�����W@�W���'�M!:��;��[ `ll��!5���ʖE�17W%�Q�K?I�R��L� ��Qu��@vA\���~?�}Om��醙$y1��� ��N��	Rq�u�eǣ��S�-e]1�;ټV"`�)�r8*L@]�b�<����\��w�x@�<t�6@�pg��h�cs�6��<tQ@�|�߆J�]C��''�SL$��j��9��u���a�X%�̓18�2�ԇO�#^���y�}4��Uˬ$�(
�Ӭ��ܕ���ީ�<��4���ivI�q���,/4u�Zؕ��V~w;_�Q�
�,�o��a�wd�64DH�D�\�Z9��r��ˢ����]��2��6\W��g.���Dt��[%��I��m�♹�������.�D�M]�dc���i`
b�7eK7�D=T��
�Z�V��f�D ��g�J~���Ƭ	���"�*g��np�|8�k�K����e�dâJ��v���1��Qڏԁ��A�nry������zX��F+ٸ��l@&���m�d�E�l�Yja��Jgq��h8�d	괱���?�x*|�(p�G��FbRc�$�-��G���Y)���uS�n�w@9�2�o���+�����+gX��wLt$cJ>����.��6�{a`�vL]rDVw�8#��0�2�e@BVl11�r�R,�h�E�N�˅^T'�2D�"_�T�W�SQ�U��E51{4
����Z_�f���c�X.Ѯm��{�χX<e���� ��9/;�֘���.l�ls.������A(�򨮏���iލ�*�Wѹ�.�5O�VUtc"��0�am�u|nӘP�nr��^LJv<�K/�6jȔkU2�{U�ٌ!�,�F��QZ���T}�ǧ�u������K�٠24R&U����'䀥HR3��7�ڝ߰gJvm;�zA.V�gO��M�~Կpv)�8Ku��X�9�GϏ"6ts���J-L�"qG,P��]��t����78��b�E��l㉊�\fTuv�w����&$�@(^M��ٜؗ\y�n��q��z��?�T��g�"���j�gb7�ɼ��	�bfU4ۖ�O����!n�n���V�c� ��!/�"�
IgfH;I�dpٰBs��ތUBs|8X�z-����)*u�O�~0jw�*����4��3�2���tR�A��ƨ1�Q7�$�;�aсۤŬ[�RY0҆��}͈gƺK����x����،|����i̔uF9��,<C~�
Nlc�/H��r	;z<��vJ1	;~��ǿ���ْ-�9sR��g�|��+P�r�� ���z�4ՠL���4^[�SUْ����h&����aʟ��`Y�
��kYj:=I-�v0,1 YD��8;;���N�=�2��֨�:U��k	�2��9J)%��y� �gS�9�!����g_Y�gHL��&-���}YM�@��R23���}Q������[�y�<��-�:�c�{�>�ޚ=s����[s�Ƴ��?�ט!#�U�^����m��s ��k�@^�����N6r1����v�Ͷ�Ͷ�cSiU#�	�'�z��2:`��6�h�|���x��N�\��2�|���1�A��D���۝֡�92aQ�����lq��Lo�����¦�%\��!i��m����6��#M\gUX�p)��f5}\�|Ý<�Ϳ�M���x���%���sS���ԧ(��P&��Ȳ�$v5�P�@���9�7���-�qf�k�kULܰT'FL�q�hE$z����-	ΤI�(�Y�;�F��s�nsD7�"��A(mRkd��Ki��
������sHR���IJ��c&B���3������k�5l���@�i�R=D�������� EВ������E~a���
�r@��t����4�؜D�f�����؍���/�&.Tᇉ� T��?Q�,vu�C���Z,|�~�i�������hѩ��л�_u�����P���~�4�6Mgø�ȼ�������!%���|!����sb��|T��f*� 0�^|^����9�!��<ϰZ��!�b�_{$�Λ�˹��*�҈jl��=ȮCXs��e�`�)@}ނ��'t�,06������W�M���
���5g)�S��9+r��Ćŀ�<j��yI'�ҩ��cǓ�Ps��)c���?P������ �+�� QˎPgF�6N��N3C�������3m���Ѽz�#�B�n_J�yә5S>�<k�.)�+� s��V=��������� ��߮)�����"��f�$�|��Z:�����u���������6�ʁ;��I0�M�� ]�	�`�>�x1��(E��~������\�*�����LyH`+��f�}�7خ"����ə6�38"N>��������|��Pnonh�F���O�4>6:����5��i
w.��Q#��=O�qS<�ϛ�*�c`��{:��OV�����QYUCA̬�/f�m��odk�B�G1�I����8�v��|�$��L��V%�j������]8�.����hWl�!������G&��˺�����M������dD>L<rV#�W:��I���X���-V$��Q R-C��\/�T�W�4*�����BEgl��C��Ǯ�∇��:Z�Q'��^מ4,�6��̮'�rS������S�=Þ_Jd�"��+,�^�]L��c��vwt��^\�$\��z-Th�܂�{����.]4_w���~����O�qf1|M|pb�,���}�sַ����5�t��mr$�zv����F��
��ki��v�p��M�yއ�9�`��6��dP�����\�����J eG��i7�=DLdg����r;2dv��?���/D����{z��wz��A �'���UdɟS;Ң]���z-��;  ��IDAT�1�7��]m��(R���&���b��c��G�(���7�h�1�`A���͚?� B�U���tr�@H	��,������h�&�P���F8d57 u|�X�/� }��:Q�w
�Яථ���h5�b��)f�P��=��C�s������Y�*j6��k-�ؔN�O���wǍ'f�({�X{0od,��ou�>�]:0�p�� ?�Hד�p�-�.���a�t'�F���9��	,�l���A�H������L<�3��g��U� �^�37[|6	
��� �駟�?��?������_�)��>~�h�4��Q3Hi{�=e0��ή
Y��`���71+�d���.��NV��jl�ŏ?��ϥ���eC`�q��t>0�r"��>Їe�������A��� �
�	�i>����I����ؼ!o�n�!�*�D�i��`#�KKjܣ$Ll6yc�Pa�Y��0,�3U�}Y:�R-Tzj�eo	�����9���=����1��6�2�nen�"��W��K~/��D'N�	�����pU��h�����5��e��cQ��OL��DS��@G$��&�"�]�O�6���4:�QߓD!��ᢨ1qy��*܈�'���4���	���r��mޥX�)'�`@���/�3YM�Yj܃�Ag��9~CL�c+�� ]�׻��Ɯ]���D}P֥�X�g�������������^-m�_�6뻎ǘIv������	�������[a��Z��A]�}	0@߷x|S���M.m>z!���$Pͬ-��Pb H�L�z�{_[�')iy�iS��5��73�>(��e.�a�
xgF�.t��6|$R���l��^���	J�z��ӧW�I:�X�Q��N�X��ײ�>C)�)\�������(��S��U=M{P��<c3������`a�Y�L[���nS�;��͖���lmA�ގR��BYG���KZ$v�LR�'2#�8Ri֔u�[7�wv�0�����naq�jR���0�h���'�T�8�>&�`4Q��_C����|��o�/_���Dw���/�+��?�.�=v��m��ۅ}�c�-tr=ٝdq����w�R��oۅ�oTE�1���˛��7$a	}a$YF�%�gt����A	wr��9
��,�d	��SھR^-�l��d�}��}��%G�*�������;�÷l�_4fN%�1m���u���cp����Ա]G�6���p�#d��5h J\�kIa�H�y�?�ГW�p��:pˢ��,���A�S��ά��A��x|p�{�o�A:����8���4�?�M��F�h%�|��qX�I�3�p>lB]�BJk櫉�����|�.>��G�â�ra��bAG��6Y�s�I�S�I��J%�KG_��� @��F��ǵ���j�~��.�����/��?ӋW?J���ہ7��L��Us���lWm9��ݝ��N�����X���;�>-������CwC!D3N�eL=�-lr��"��1zB`1� �y�CB#�=:��U����w��T����Y��a�Ho�ͦNQ7��l�9��%=$��^��'��+��H�Z��/������_H�-`U�v�^��GJĴ�$"N���ħ��q5�v3��3��?x���!��V}Sf 2��	�=�N�(�s���^���x��2玲��_�d��U�u�{X7i�1f+(� �F܁̐�L����$�^W�)v�a0��n����⪢��H�]l$�ߣ���yk��8����n���{�*T5�f�1(-�a� ��/�����B?��[�L�n�:Q5����ו}T$��S�
��xX�^/����$�������Ŋ��5�#�D�2 �R'���9,m`0)S+ئ��h�2��c<�����"J5�>�6w���Hq��e�}X�����$��P��%���-.g�qq��_�du��_8�/�S%B5<`�2@�e���ܯտ�-j2$PO�:�o�#y�}�>�u5��E�&�ȏ&�آ����,��߬O�w>�j�]��>���=��Àŷ\�l�3�ήY�L�E�׆T��B֣&�7֘
:�f��I>�����t�q,��9�ߜ���˗�Ï?.L�N��n_�ϖ����w��n��#MM��2��\����NRrb��FY;�����),"g�o�`L�:[o\e�4���K��;6��hd7�d���}�	0,��{�w1��>�R���F���)����ԉ��L)�o��b�>~�����g�M ��B_�{��x��Rr����X��`�6VE�{�ۈ	Bq��!���;֍~���/ΤS5Tq�����w�1��ݓl��[����s3V��G�wVE��ӱ����^�u)Ooױ�c�1�� ꋗ?��W��3�?c��Ç��?�Z���;z��ɏ�O)�Y�z+������]*� ��x)̃= �%�f�w���|E)�"ꤍ~�)R�q{��ޒX��-%�	FUa�U{�0��X1"���h#uB+�W�5��6��^���[���'��q���F����ơS.��oi��5>5��9p�6'�=,��,Wҡ�b�(�)0/����t1����_����ckf���B!���ߺ/�Dm��I4�z��D���(L�8�j��Y�*���M��x����0� ��s����,�����P9���� I=�.��ͻ�"��{�û���ﴵ�/�����;1lqC�v���N������~j5~��^X�$"�^��Qny^��ifwS���'������e_$YK�"4�������~����'��r�}aHhu1h�Ƴ,�kC�M��u	k|=>����ȂT�~�Bš�6gr���N��ϟ�
�v�y�;+��VwT��E�j��hUh\�}��9E>�UJ;��� Z7o���LꮔG�h��K���uO%DɬwS����L�\uo�C'9��A�����{:uH��n32&UW9*��z���ؕ�`�>.�ݛ���۷�G�Y�v�;�������lt��`�U �K%R��i�&��0�ْ`��T+����>����Hr���.i�,�D��|Ĺg˹�%�K^q}6X��7�c���:e�
 i*z?�4��Ȝ7\�����IH/�3���b�8�1=��zb��pi��#���|�5���U"3�6�pD��B]��="�X��+�3�P��[��̊���s�P���.���3!&Q���Qk��θ���$
�a��2��J�G{�;���."I�:y z��i5�V�����ҁ�����fgڿ�ce�XYDg4��,�?,�9�b�A���}����k�Hu�qN�
�m�X���p���֮���Ǐz��g ��)�M��/���3�>G���?ο���/��~x�R�wʃ��.u���?Ї�=6�! e7��?Ej��C#�X�q��kw&
�$�tYl�p]�y���H�(�*Dm���|�:Y��6s��%%�g�ZTq=o�-]:��ʙ��@4O�z2\Y[��m8���c�1R K������)�P�_���1�(>�v-%2�h]�^罨�~�(� }���U�it؁^��Z���UN�]�����%��V �YT�X{", z����퍈�B��TR]��e9�[�=�U�5�J����U-��/��Y�|rӺR�;U�y`�1|�W?��~z���a��g�-�[z��+��_�B?/?\�Hr���Qˑ�;ֿ��Oɚ��eX�׫�(�'��zQ���nN(�p`]�K����A���t?R��6���/�	G���Sǚ��~���U����=��&�u�L��u�v;߅�0����U���I��/��`�N/���h��{t���n�������E|�&�ƹ�y��{��7�����
�ƺ�Xh�s/�E�_����O�M�z��=m9Z��ZB7��\���!�e�A�Esf�H�'��G�2ڵ�)��<T���@��\���u�|�:㴀�Ze�O6�I������N��@���y��ai���.u��r(��i7Z�!��g�-����7td_W��m�����u7s@�������&� �rõ��b�A/���!�a]��T���g���=3��Lh�	�4��q�Zv��}%9��0�v�R��Z��'��7��jx@�6�H]��F��1�kӛO"�P��o�H�:��u�ܧ:霸?4�ʈz�`�M�s�l|8ung��8��4ي����Eey��F�⯃U�F#��HW���j9eu�귱�[*�h#i����3?�S��u�D�QU��}GI$n��Uo*�_vYj��Y�iv��JF�=w��٘�(�L*��o/'^a���.�xU�����إ����
��`50{m��z%l�:U6)�N��j�D>�*6�`��T�[��Zt�@�o	��L�y�g�/iiڛ���Ԕ/>L�_Ʒ�a�i e	PͲp7���%n��Sc����<�q]@-&�z�� �o�
��+t�-1�W��@����@��XX̲$z�-�R�I�3�l��<!�I=)��m4�X�K.�����%�)f��%���ɶ����lm�Z����ŪX�}��!>�rC31/�]�� �g/ ��*Vt����V]��E���`_v�Z�^���}���C
;QhRI��4!K_�zo�������o^����&�/��-�����}����ꕰQ6��'��U�^���,��%�����$�AZ�=��!�K��ʄ@�c����e���ӉQ78��y���#"����A�w��g8g,�|ӹ��h]3#s��a�7�kWT��#��0��yH��IZf^�6��n4�Q��ҵ���dH�5�%K�T+-�PgMO'�+�qJʻ�T�mqT����1%+�b4��|��.�-aխ�m�$��?���o�cf�_~�E�0�����3���K=d�Jyd�w1�a�N���]9Xa���o	�.�n����g�x��J�m.9��\T�)	.�p<����^k�����"�Y������������ͭ�g�A�̏�h	T&�aK��K�,i��/�$�"r=��%�+�yJ$���2���!����1w��ԡ��^���S��8a���I�M��X�%�紞t���
p�Sm�+ �n���OQC�13s�������|V�f�'\�>-?�0�i�k~������O?���L'�dP�2s;j�T1@�������M�,��0sk�a:�����~_�ux����$ᓤy4y�;�D�ɢn`�_�Z\I�9����̐���׀R0��l��f�a�h�݆u�U�`��%����͎�E�X�+����N����<�N����n���"�k�o
�l�������K�������"��⸿���/��˦�x�Qc{x
��4ӽT@�͌�%�*�p��ټ��	\�YB��϶l����A*kACN����
lkv�c�LMf�g.��>z�ӥ�V�R=��ڤ1j�1�g�ʹ�{�R_�����uy�N�?� Y�G���_�C�:̯�e��'n#؝[�������
�k����ʜ����Ή6�m}\������H$Bf��Y��r'GՑ�c�xf�9K;�/׭|�#�!�[�^t��Ã��3����v��;w�ADg��E�?d�� Ơ>�Z���4��ncm�R*�f�|F*���	�g�LH�\a��W��N�$�f�E�,�|�*����|��#? ���@����~�о�����3�m�;�&����h���A����l����5s�	���^,��$3K_�����X��ŋ�!�a�G����� ���k��/�htZ =*���d����x%{3nV}�{(�rf����,�'�����Pf��}M���z��G���Z�G�D��Z�7Y�[;�S��݁?-���� ���Tr������ >g_��uܓ��U+O.W3��6�c�5FJH�p֮[�;D��?\�PK��N�U���a߀�Bq� |i҃b�{��ݹ��W0�>��R��u��[t��G�~�eb�Qc��	�g�"O���OT]"��u������(�L��לQ���<O�1����F3Rx���	�E�.�l��p61���l��,Ϊ���Htas��յgn��y[0���~|�ra�7bH�<�&*`q�Bl�)+~Z�]9�M�����x4-`��r,?�K;-����a����A,9�y= T$+��^6�ya�}BI���s�����d�X�ᨎ���EQֻI�թk��Ŝ�E����R��:�������r�J/*�	�,nw����uM$��s$#��b��{��(#���әK��O��~�̕>�W���t���*ْ?��1a�4�qC�}~�Bexb��9Wԡ�Owܙ�<�X�EK�^Q�"��(6W���Hì��󶋲RK��'
J�^7�ךg8��kdng B�9>�����T��EX����%��+}`�[�$;�W�ɺ٪.��C�F�A7@���Tːp;�Z��������0�0����D)�(��R��2l!{;�Ja�8�s}����̢�Yg����E��\r7��X�$B��a�Kx\��8��r?��A�'�>M����{��n ������Tn�\a{v�ɒA����H)8����q�.z{+Ǽ
���J�sF�D|ͱ�ޟ�]���c�3������=q�����2���Ó��q�j|<��4DTm��qmͩl�vY�ۦ[0/pI?g���j�?����P���ލ̊�`�`q5�N�ͭ���C�P����Z���t�I�?OC���g{c�0���w�_���۷�����>g�bc��t�d�5y����S��{jv�W�u���7���\��o��￳�� ��L��4j�>�;�/���4'K�̌Y�Q�$�nj�3�dvX�{��ӼF.e���a��y�d�=a�v/��(�f�r��]��1�:�N��_��� 5�'�4W��T�r�6}F��(����`�U��yR=���${�l�C72�O�??����.��e�'�
�-��M5��(k�K��U[���ナ�K���Tn��1ES�9wf��r�ׯ_�o�={���$`���+r��{	�/�6)��M���N�����?K�(����L߾}Co߼�2)�3J=�(�nn&"[�@3��T)�E���Y�1z���m��=W�[�^Kd ��@s�=t���Hɧ�X�}�`sQƖ3u����Uu��й]b���n ;{�r�+����W�~uP�S Uu�%��I��'˖��?}�׀��س�n�%r���%y10k<�iY�d�-щ���r�[�͵����{��[�p����3��I-��*c>���|�������X����c�z��-������/��ka˓뢊e/i�J���o.Ë߾yK���?���N2N��?W�����`�ZQ�e`��S��bs�u9�)����wz��K9_\θ��l�|9��:�[�>�b�$ђ�(`�[xC�T#�jUDo$�JuF�8��k���G��p�S��L����F)q�1Cc6Ja^�iJ1���\#=����Çq�z�����^���r��j)��!EOs���g�q�����K���h3Y�Љ�_f�r�P;BG��)�2�
S�O��;>E�2��5Q�9�8���_n�s���3sb��W|)�k��b�}�å��`]��IJ4QI��L�p�����޾}G�?��$��,�`�����x��Փ1V�C��ϹPQ����������"���0�����=�%�t�����GN�'b��������n�Z[��϶�h[*�5�2�@�sO+}b�0�f+9PA�~�z?�:�rξ�N�`��<hU+�Y-��2y��O��IU���XDV.Q90�먏Ɯ=F�&��w��Կg�����|{�ABa�#:���B����O֡Q�����B�M��������sV�i 3���a���\i%JX����g����Pa�қE�eQ�l:c���Yٷ��@��,�KUؙ <��G�����TU7#Ts}/Xi�zl��x�)��$L��y�LA�c�=�75�����m�ע�e�0ڽC�hφ*n����񱱠Tv7���X��oLdb|�R<bh[>�]��>a�$�I����l�ɇlBEY��)
�����/�Qr��,f�3ʦ��JV�6~�o碠�Yl��RhC�����QNfN߄�Q曟s��>Ѿr�w1AO����O]Ӟ���t�&�k9��ܥ��
���8�/���-i���k0���j�rf
�vR�7iȺ��=ji�ٮ��T�c6�믿��k6gIz��6��ɽ� ��4x���쁪`40�I����-l�/�?����K�Ø���~��>�ua�N�,��j�%_�#���7��]���h�Qo�YQ>�f��}N����2T��k)+�^X�d�@�Ռ�Q��j1B��L\�,�ڴ	�%&�����Uy�j��~�L�":�In�6-�cH)ARV�lPxY, ��s���Fj@�w��f'��򳡳�w��wd)���}�����L�ͩ:�|��x��O�2��d��ku�_�=�_I?�b�:�SP����s���>���P�x�Jl����q�Ȑ�&�9Z�Hܧ��0A�hm�M��)Q-��.V����ۖ�.5:����q���'Θ%���Z4�h>�
�R�u�G'q�7�ԃ���8�:��S.o"%��/r��^Q�����hY��۱�b��i.�acU�,W|����]� k��ހ#���0vnR����b�o�H�ctPu�V��6�K��'<2N�I��4g`�~�zq�]���9#�qH$@횈�{;ʥ���gx���]f�eP��u�r��N9́8|�1�Z+�~������zȴY ��j��&sC���32H%}.Gѐ�w;S�ӽ\�`~���=�u���Qf�a �f�������f�����FJ�����A�\~�H4ł&&���8��fY�A��E��I�|����8_��]�
�^PH3���ndH�Dv�&Uu�j`����7+V����_�=�V��+~���\�["�����#��:O�U-�q5A��u�llj�pi�r����z�ێ�R�v�pr+P��Ƥ�a�t���8��� ���>��h��x�l�*�{�|��u�Ϯg��.�P?u�n1:r`���ȹ���D��o���;���
@��#?"_��8�]�ɝ�'�	��C��AFM`\��� �=�wM����
*���O��f\3��,�}4�1����r��H/��7��x�#n�'�(�Ժ�y�PK�(`��A]�` c�Ȁ5Ih�$?��@�N������obo1F�?���r�j���[���-V�Hf�"Sw+Y�Vtn˯��|�&��fŒ2p����\�e#�}LC�ס���Q =��� 2�VuG�{ݯ	���/��,*�{Pݱ��u�d�4�v�@�����}��ga��-�`���Q�ZA8m*ד���P����;ϰ���x2���ԯKyt���LCN��3��+�3�c��� qy&��
c��KX�ԅ�9�c1V�(�^���t��#�]4E?�Ə�f��_eD,i\9�٠_;J6�f@��i�)oV�ْ�0��uH�
�J>��w_MSW}u�lX w�g�SRNS�V�
T��a��`ѕ|��V7�Y2��e���Z\����G73�f�O���	�gҙR�T:ݔ,ξ�{.�ۃ�yJ<�5%J^2��̱�#���.�#�fdӭ�i����O?����<�-��=0��)���5���wǺT�5��_�����lLZ���L2�yR����4��󎧏�wq��S�IT�@�IYR��9�2�_`�1���c�P�.J �N�v�Gݤ{�v@'�N��^?��=#����ǺV�e'�ɬi3����1=��Є�8��c@|%�
�W
�qi���ZMdA���`�q� ���&�*����X����Ⲇ��ߩ��=��DYч02��F�l��2�-Z��P��H�y7�Y��� �32�g��bQ��u�7�к��>zUU��ꀍ}��S� � �9����W�/��H�GRBہ,*�J�E�9kRdۘ�*���.�<��~c�Y�\��x_�|A�����^RQ�i%�<o!g�O�K	�����G����>1*��}��(k]r���>ڹnkGM.9�Y���6>��&"��T���uTRjg�S�;�������>>�k�T{�_���P!@�(��.��	����T1qb ��H�`��`�&]�<����}�>U�?�7���~LBWg�G����h4���~f��U�w�R�s�GQ��~����,P:�6c�_A�\���>G{z�'%7�eB���r�J:���7RD�U��VM'��
���u@��u��N�d�P��3�U�~v�7��J�/��l���3f��Iz�㉜]^��N�?�29
�?��ӟ�f�3�����=��SW��b"��}�I�ɔ,Z�~r��	s�u��`Qg���5�uDu��#��K�ʧ��KٖK
��q��,5�zc�1V�bg��@i��1rhC��	E�YcsDJ:QUxi&&V���䉶E��ZqcS�a�~�MR�'a逃�"�:���q��{H�7��؞�@U����P'��M#"���)Ƴ��@�C4�Y�]�$�?��ru�[M=�H�in�}������[�di|�j�⨂������y�߯�Ǐ��PO^؟��_u�X��=X�EsN�����"N�V�����Qt1.̏��f=���G�ߧ<��2/�Y�It���>1d�	9ky~�P�"`(���rR��st=��� ���	�ì�>��iP%Wqh&��9�e��1���� ��@��W�
Ʒ�����"�A���V+��J���0ZIy#K}B�|���jE֫�U`�`��r͂�����Ү��()�@\��6m���Z�+�]����ck������b����.N�Ǉ�o�/l�WO��������εU��=9�|�~�ޕD�p#á�5)��gK� Y���6�e���Ա�H�<���}��>�S=��jē�9���J������:�&���ۄN��a
�����Uݨ��Z�?|�����J��p��F�9nY�� *3�唽��-B����������b�c܂E����Zϻ�`�FF+���|r��ì����c�4?�,8aw5*oJ6�Deqa�mf!)�{2}���l0fjnT����O\��A)޿�:��CM@
p���y*��MJ}P\nW3%�g�������(�P`u�D'�W\��틸���>D��}q���fBz��,��U4�����L&��Wύ-=�bd\4�ڨ�z���ٓ��)��鬟�l;�5��fFn�C%�dȚ�}h��Ǵ����^�Y%J��ל�폢ED�G�ݭp_���ђΐ�+!���e����v�����*k� �kx�H	�5�v&�Ƙ�����7�fٖ߳I��c�Y��-Ue���"ϭE}yt�%i�"�+ï/b�_A�x�8���~��.�Pb�W����(�n��t}��>u��K��|�B�c}����x�/�����k�|wV@�o.�Y�	p��Յ,�B�2���,�0�M�ϲ����A��w��ʠpX��^͢�*ڧ�;��!�T�E���'���Kx��Ef�&nw�( Gv��d~��(��+v�}*[����b�J�=)�P�5��iL����������)�@Zn}`���^d~����Y��D��v���j
�t�S�<�^,?�3�����p5CʛO �݁���P�4D&=���5g��3��}��ƀ`���w���/��ң�vح�-$� ՏQ���~�*�av$1]�Zq ��E t�ł��r������m#Gͭ���,T�OV��b`Y,� �Z`j���~���;�p�I7�'zţ��2k�U ���-�D��-���I�zo�*�I�>�ǫ�כ|㾼�������:ՓOqL~x%�c��U���c
��_�Ṯ��'p8n�A�>��r��%�}��M%�;aϫ��{a��7f��r�e��j�z�p�n�e ]�G�t[O|Ĥt!D`�x����hCAu:�;�`���5���L)g��E�ʐPC��7*��^/c��5@��9E^u^��SO
��0��ȹ~��V��&>f
p͇I�=�Y3E15��A* �½�Ĺ]X�����ˋLu�?x��V�w�`�G�戅^qARg�5pe���Nic�)�ЌY|
�Ւ�=��z�|�a�@�Il-ᓯ�USӃ^��>�*u���@z��������*�"����~x��;��s�aB~�~��PĞ�ͦ�zT묊��NM ) ̟U�%`5nXkZ��b1.�Y ��tw��'� 	�:�r4 v�YB�57���-RI�6������h��[�� ��O�r���N�� �`��R�����>O@����s�bUC�%�u���3 ���D���#��x��?R�@YM�yN%�*���<I�׻w��Cl��Gv�-0�=�[Hx#��~��4��������J`�'$ ���u�o����!Ɇ��?��a�<���|?���eӗ�N��~��s��X���?n���}�0��߫��I�Y�a�
�!X��ܱ_�������	o"JO�@]�LV�Bd� �q��u�7YL��P�ذ��?�����|�H�Y9GE�":b�^nû�k�D~A�c�tw}���=��*L��K��u�T��栏sX'���\�K<,�Cƨ@j�C��Kw-'��u��ߎY�&+���v^���񍒣�G��񱮇?�/۾�X��L0q��MpzI_�F������ǧ�� �:�c,��,4c��1*��g�]f�7<�X��Lf�𧫓e���ȯ�DZ㪻�
��,2�����ߟA�"ƭEyLm1�3#t�t���%g�'b�;T�4;QS���U����m9���bO*1M�|�}ڪ���_�|z��+��G��yXj���*�-'�L)MXa��Fɓ� ���eSDj�;"�-�����]�D��f���-��2��2���ܩґ�蒬�h�.}�X�1��;~ן�>��P׺'w��NnL	��z��ĳ>B�+[�VF�փU95������������ɏw����%2���㰹�;�?,�$(��%�>��zS�(��"��ja�E�+�v4�����P�6+�B͢�����bg�h7c��;d���c�
:�4�<ߦ�9�YP��3�Vu%��9�S��&�ɲX�վ��α%C����#AT�=k���۲��NR��X��,�ME��nj�R�h/ύ��60��/b���Ħ�����̲�H�,�l��n�~;rV�㞞��ԅ�a��.XE��J	�)���@�}x�3�����y���SqY�]��I��: �q�ń�[s�o�q�z�@����m}<�� �ݖ0�N=|3��Rz/]<�$Q�fYTY�k�%2�%���_����wfӗ ��t����C�U<�=��t�A��ňK���#�.@����PEN)���A���2����	�݀(w��=* ���0�y�h�R��Y�T�:U�)�S�V;���Р9ϯ�G4�1�i���|R�����o7-��T�!�����qb�c�����
_H�C~U��x83MBd79�����2��v�5e��)���_��K�)��)��.ǧ?2I�G�p2%q�0�Q�����KWL��)R>Te���],L7�2����h�}B�}�s�R�Y��/�5�����;a#�F�r��W�~�ϑ|��y��+��n�?U؆�]|�?��A�&�\�S֕�~������TA�vY�p�W��)e[+9� �s&j� @D��{L$�/i�����κ��	*��k���'��w6�8W�|�K&��3#�AW�k!q �^���9a
@�L�ik�r�`� B���|��\�w�߸��k�R.�Tӳ����7+��d�Ғߞ����A���Zr;9�h���#K?��y�L�W9�����t�H[隭��'����Ӑt�,`������tE�&��r	g>�ml,ᆜ�����������ʖԽV��r�n���DO���K��e?���i����}RmF�Ҟ�K'�F���CP?�Ey�h-n��1!�?D��?9�������f񎯉�P$��{r���@�[� �#z�e3q�#$^.�H%��qO=mPWy��O�ِq��7�,z#�s���L�� }7��6.�O��);����'V��g��ʫ�� �Q_�M� ��퀚k�b���E.���)�?P!�gQ%H٫$Ο ���=��Ņ� |����3�+��`2�`@����nv7����?泻{�-ٗ� �9�ɘ'e�*�O�!5��ds1#R�T܆�`X�X�\0-eP�!�z�v㌩��'�����T��i�(�i��4]i�H�LdN`{DTs�I`�Q#��<�H1@�O.�X�o�6�:$�i��4} b$&�~����K�G��e+:��̐G˴U'O,���"ѓ�-�%�bc���������BfQ?�@�-]��f�1��zljP��Y��!�^���:��'2T:�x=���|J��� <�n0�̷͵���c���b:���ݭ���ͭ2�4D��P��O)��"e�Q�2����8]>��m����fúZ�[6�-����=Gˈh�9��O=r�"��(��K̟g�	���( �^'m|%]�D���q�H&�~�̾�l�r���Xn���z�R|�������4��>6�}��*i�J�!���ƚ��D-3i�1]�Ly��d�X����:�<.=��ke�`Hk	�\�������z��+߮L��4j0�/���D�Kb��"�0�>��������a:����F��|�v���$�8�s�Q5���
r[K?ǌ����#(���Iۻ���s����gi��Ǌd%��Qe��
�ie:Q����L���D���e��dA�i״�����f�� ��f�k�N�_�~�>�5K�޺m`O�D����w��6�� N6W9P �&�sT�Q	�-�_���9�M�1�(��\�NTF0<{�c ��&RN���Zǟ�P�� ��.��b~O]����O�:fz��s´�t��Nf�� u�g�5(�� ���%�6�* 'T��1�.���{z��%�x�B���۬�*߱(�.դ�Ia��[�QwWf�q�}�O^�C#�u<���	w���+N9�Y��>���'jy��$�4��\��x��}.IOˇF��m@5%�FI2�[��(��"�5F����=U�z�0t�14,�á!}x�Fi������y�?Pa�]������l�����E�(I�z4/�񗎳���I�侜v�f��]Zl�OЫ%#)����r>�P�HXd�
823�������_~@��!XX��#Bҧ�s�:B �t�u�٠�li:6i|C�j �BD^��G�y�\��w���&�ɯo�i�V�j`��$+th�;���5Oi^]����GiCT���}�}�T�(���[�|^<'k\��7��7"OQ�G=��p����Kj��Բ����d��P������b\�x��D�q9�%���<������/}>(�NJ��8ß?�>���]�R���d-�.=h�V�dCP��L��X�>J<�֕Oo߾���rʌ���	��/���T��fʠ	�������s�����+b�a5�j%���SN�~vm8���yx�+j� 0�<?
%��&���\	_ݒ��/ �Y��Ӹ[���.~��������W��@PdD��"�Tζ�4o:��S���oQ����-x~��y�+��XU?�or�6��G:<I
��'�Kˀ�s�J�� jZ@�[��2����y'�vY����6�˄�1�cя��iN�j�l��[;av X�-�F��zo�p�8�c���$'��o߼�)�΋+��hb����={�̷zL6�I�j�h�:K�;�뽥#���� 9��p���}/� �;N�fϤ��0̶�'�f��:�,q�Ci��+�5��l,~2p�� �D!��}-5uX��[�ꮝ,�b��,���K0>�M��&Y�w�A|�%��vc:�4璔��nH@c��^������؋��F�{�=�̇�)��J͛��
��D��tu8+o=e��������ǏO�����r�S-,�`'�]7��y�V�m{�PY��G-Aͯ�����8o�1&0�$N�?���D���S�zޏQ���T�ZB�����z�����>pdmy3�s�[��"|	 ����	,�`[�D����Q�p�XSZ�k�I�=U]�ⷼo��1^���I� 0�<,磦d,�e%�՟5����43t����q�?@������ۖ/�S_��9�o��#�/��`�l���"�3��z,F�.g��Ey�}^<>L��޳͑Y2I�i�[-3ұ�ew���ؽs�<�̌F-��wUE2�x�!���"�� ��L�D^��J���l�L:�q�_�✮:�b�ȓ���$��"8gbg  ��=�'�E� ���<��>w������������ᄵ��#'~QΕ�}3�ɻ��5��
(�2w�=)��A$Gv]�̚.j�@��*I�U��w,!��Z�w��s�-�Uﾞ�L�o����q�u�?��Y#Q½�ſ�&u�m� �t��̂%?�ڀt�6l��QL�Kb�닚V,�w6®i����f�-��\��ȋ^v]�����W�U�������[�k��>�]�����?���]�K�G�\���8�D��s�e ��ǥ��f/���HX%�O�
����-$���&G�A)���e�R��ԇ���D��h$*]\8��+N3$�L��'�7�N��H6�E�]%v�.u��x�;��n�[P�~��B �/�N�e�ҿ��V�ڕuV�O�d/;�[��֠��X����=pܾ�:u�⅍��j��q��q�>��`��Vt�׳�[��zz�Jm?�,V�K;:��%8�;�� �������]����S@-��ۘFX�3ڸ�_��X���q1Jm֯ў����!�\�ջD�z��G�T�<����:�Z�iT�&1��-4���%��ZJ	g�+,.K�yU�?��E���G�E�:���&�7/����5CN"FQ��܉vq�if|o���>/
�p�~dR�q��Vz��DK�?�zgl�� /:Y_�[���������/�t�z\������ҋα�?��	�L��Qv�>�۔���i�������Ƌ$�7��m�i�K��Ns!h)J�c�Q�p�������q
���_ �PL$y����&-��G#i���W��-�F�j{?��J%��%jKh�[OW��g��*�E��1�W=��Y^Ċ�I�/Z_W�S?����z_�zY|��MTc�-��.ʨca�vD��4բ�}������}�~r�a��;�Kj����(h>E�"��l�zS'��<����P�rM8���]�b��M�d�*U�\�D�*qS�ʥ`��a*r�e,z��_�
���� `���j�(y��S�C,�~V���!V�-�B�\�1��'si������z_w΀U��X[O��\my6���>йsF�a�U��w��@exA)�3m�R��g�/��rS���.e���0���V۽��ۦ"o%��ߪSu�J9,��s�������i�ZOt��;ʭ��u�'�R8Eٳ�>��5�T"��}���ߜ(�D�$ǝP���� }8����p�ݟ��[�Oo%�fx�-��9 ��흹M�a� ��yi���7�C���h�1����u���Rur����z&�X�Y"򤠴���"V8���)w���z%�����G�k�)Z����H|�V�}�0D�\{�Y�r��6�Bm4&~ѿ9՚:3&8e��l�`�3x�4S�ip�XK#��������p�~���K�W���_r���&� �:kgƭz]���xB��A4�Ȫ����U�N��p3���	E�rS�$=��~�C��ȸ�q�t�
�����_�o� ʡ�s�h��R4O�ў{�:p��T/�:�LP��V�<�z�Z��uJ��_G��K�c�0ձ�Eu���1Pm�G���M����ZZ�͋����=�?��~~3jE�:W�z_O��8��(3zy�+W���6
���	��h �sp�s	�d���DeM\&J����<$�|g�d(�>�FX��<�Ӊ%�N]o�w�m��f s��:�Ps�)H)�Tq�|���nLT'2f�w��Ond"q!����n��͸��ӳ��V`n
\zlR&��Ts��gi��+���VM@���uۖ�Z�Mp�Z��Ӊ�5|=�{k���jYNwv������"��r�_�+��U�➰Sn���wܙc�9��<ƙ�59� ��Lq8���KE�ѿf���b�4��^D����'����
.O�b�\V,�>�t����@R0h�����i����6ս<�"+���[������J�eMhb�":U�T��"doL��hA����@+<z@u҆�[lwIeT��S��[o���J0���/OM��?�#�"u��(\�tT��t�oM�7���_�E�^++��;mQ�� �s=�;��>'�mb$3cA�m����D�+q�Π4d3�/�0�h��0�>4T�nT��.�I�'�:(@��iP)	H�q����b@F���N�����њPK<���ɽ('�,W(�z�=O��u��nME�E�?v���*P�s��U�����DI��!�h�Aoam(���؊�1����Ƥ{�ܻ/G�@
��Sq�aw��M���)b�r&�	���K�'0����|�5�D��r�JP'v�&�'ɍʾ�|����oI�V&8�Q�S������Mp�Y��8��{0���b�n��(D'���,���C_*˾�J�(`�8�)�q)I��=}\��$�	:QB~�W�a�����u��c}�@��?����-:'��z/�T���N�o��~5<��Ӎ+Cڗ֔��K�޽2� k���LԸq;m�V��6ʗ����i�!}A�-�+���$�L�_"j*�ᷖ�hE�F5�����0iZ��x�z.�����e7�h�smk�G%"%���DMB��X�P�zhxQ=()%P��-.:�yQ.��S�#�	�:��*o�g��U�n�X�t����a|QA$HZ�f3� �"h���X4��Z����9��U���T$Ne�_T�K!�������Չ�&�s�ٽCu�V uпX�D{�U��X�ݤ ��D^JvD�MS	(�8D��w���;7����m0��+��I�o�&��Q;��Q!��DܥZ�䯓���$���"���4$Q�%a�#y�s�8M�K�!�Mg��	dLyB���O��HyF�+���u�<Ȟ1�1�k�~�g��4��g�"��m�]A>��:��^��q�~�7��n7�� �w}eѾ3���vY��;\ >2,��'U�� �_hfuA�k;å=��zC>���S_�Z�V6ǉ�c���
=��&��F*0Ÿ��;h[T��������_�!�"o�P�_���JD�]��BpǺN@'�}��
�ׯ���n��DW��/�X���B#q"�B3�}��?G�ڵ��9��T�e�R�T"�d����u�yQ(����N��Lf�D��M�[P�Go9�Ǯ�,��y��z�t^�ό)=F�Q��x_u��w�sc��E���r̀C�k7�L�~=G��Eْ�m�y ���|��]%e4�w_UHm*ѫ/5O����_�2�9���s\1H���4��|>%Z<e���ʸ�wk'�иN5���<�4"Q���[ؘ�ݺ�o�W�ǝm�rV�}z-�n�U���+[�s>�>����:Z��x���n1B�<��'�8�9�\"���
��&��V1@�����H����U��fl�EU���GV�c�(k�?$ջ���|=X
���B�p��q]$�kt\��r����\��9�
!6�X���<���N�r�|Ba4�++�Ή�'%
J&�iBK��%�
��\/��\
�k�Sq�#��ƁXgpE�n��h��c�]*����z�7�y��#�h�7P;��[�So�Ͼ�_�ѻen?����a�x*��~�ƺ'#t�oԘ���[�{}"�aQޥx����ʠ-׈�6S�X����}�f��>圱���>n��0녥�o�xT�����Bsծ�������|yR������~z}�X���X=h%�����VI,�>�y�t��uy�xޛn�m߱_���5w9¬z��y�q�	56����'h0���)���Aa�C�bs�j�e�l���Z�]H"�&�b\�ߏE����?
#+|ӏV�~9�;�D�(�4u�y �(���>8(���cܮ\IQ_��.�'F��N�U-
�׫A_�jI_�UY:y2�49P�g�ݴ�t����q��(�Z��B�[l���=�3`��dȡ�}��@0�l��C�?���*���g@)�`;�a���y�FN���C1)��I���Kt��H�Ro�0�S�U��+���)=p���{,�g�\]�~�
h��9����2���{�_���c��\h�d�L�\��v��<YsA�����M�Q��:_��x�P��ʝ����{�ש�C�����(x�?=��bR��	��}����z���>�~0E��P�Ϳt�fzbԕ����Qm�$��[]�ĭr_}ł{ZG�<󹨻̉j�$�����H�7�3��� 5�R#,�{V#�i����J�^�6�����W�icE�z�� 1�!q�o�B�^$֖<��I){��V�PD�N��"\�-ѾxP�3��To�i�%zXyVG������x˻�r��w^�wᐼ���'�6�>
���獄���b��T�aS1	qp�O�>[����a�U�:���X^ZF���ڇPQ_�[���j�&挋<g?�&'8�
0nR]���ל��x,�CUˮ��װ��� 1����µ�oiI�7��j��⣣*�q�3�ܵu����`�?��;���2���W�S���|��,�o�8����&��=X���sDs��#���{��\�?�QsǺ�"V(2��PD���q�ol��c�r6��=��:��Y_:�G<P�\�n���cl�*��)v�q�2Tв�)���nK���Ձ�X��~�w�U�vܔs��v�=i�����&&�^�1�_jϳ���:��E~�w1:y]���/nb6�(\M�5�f!9ໜ��e0P��5v\�;_#���\�x�ۦ,>�->ɭ�Q��ɺ��No����8�z��_�x��ED]�F�R:�=\5q��SZ�ܫ'�@4w�W}_%!Uꌾ�?�g�@�cǈ�5@â�]��}��a"vD.���K>R�wYO��~��\����2��=6�M�fJĝs�F+�ôfQg�7��֡�R�$moM�s���{�RFn:��l����ܘڭ�����{�����q;n���I�]�ʥ�d��]W���=�����~Vå-�3ʵ!��yu�>[5��0�	v�[}_�mu��s�x�:�/�C׺V�(J�ߏ1�[��7<@e1���k��F�;j���m��LK"�Ƞ�-Ke�{��f����S��'\�����z���ޙ^X�L5NA\E�z�5�}lJ�6Od��r(��@������+8!�{ml�8c�(H��8����_ O;vd[��,)Lk�;�rO��]�7U�v�g�y��S�=��*ef���5��
�j��,�I�RF�F����.����>���`��uG�|@ã�s7��[j
��=�O(�H9�d�(���LF�lb�Q-\n��ZVޗ�("`�~i�Ȋ~��9qi�N��r��HPcq�n�K	dK�"�����i�lJn�Vg�^�R%�W�N=qL��\����J$-�}��T���+�@�^��6�
��g��~�A�Qш�����n�x�^ߓ#��� ��62N~��CV�K��$\�hW��1��O]��O���Cd���G���?W۝��)��c£�+G�^�����!ۃ3nU��>�pD�k�oĤ�ͬ�:a5щ��:�a�i���'�f�׺O��[T�v+�Sݩ����g�K����g�!/�WV+<�ܟ{V�w�I�^��1��\��>8���q���]�k��9W@\_�䡭�N�n$5��B���.^����Nr �A	e�g*}���F�J��]����$ب�0b�҇�Q�^�;��0u(y}^E���gLWm�E�*�V�7#�#�d���wд$0ׅj�� ����kq�M�POp�	ݜV���1^����-���fQ�$�8��z:;#"����9BӃ��=,��(c�ǡj�޹d�tPW���s��JU��$�6N5j�¥֎���E�MR�M�����WO�����W)-����6w]c��T+�[����|M?'B�Y���ÍYo��`C�5�Y�Tʋ��]L�0P�����wb%0�J�[��s��E��L�}���>����W���@�h[K�i
b+���x����	�g�	��K�;
f��8���t����m�(مl�4����"WO�Qܘ8��a�d�v�B�1��+�!CD�L��} <������τ�x-�>�d���R�����{Ml�W��ӡ�g1=�{w�mS�t?�e�Ux|���V$'87Y.4�m�6�a�����z���"Z`�>��S �R��R�ґ�LTeP'?Arm�^��,�v(!t����*s���=K�0���Đ�MJ�%
`�Z%a�u3V�k�S�{s%\���]=�Ym;���R�59DF��/�B0��T���&�M:�t�^'���^J]����&��R�_�O�
 .�iee��K%�q(�G�=?��)�y8��'�Ƨ��ކ��^�w�X3(���C�Gm$M_�XAUK{p�o\�ܫ�O���!�M�n ^��F떄��2��-[6�Q߱���<����2Imژv����y���7�}�Ǹ�Ҕ\l EY�C�P�"�Ƴ����쯡��ٲ)��Dّ�R�vږ 5Y�G4�"��_l�q��p�DG{'�_d1��}���}�b�P���8m�|4ݿ�~�:�]�0[z8�6��݄�y��Mx��yx�����ٔt�L�黯moc�j)��JvPu%���J����)��)�6Nʪ���9�}hT8�{�Wذm��q�x�҉�v���0dc�\S=f*�8q�c�X���a??��4l�l*��ծ�PO�|\kۗض���W�X�vPrd$N�k�)u�)��� ��P�b�D3p�	��+��c)Is��T�^���$z˻���E��4V�^��/���tvp��{������ɓp������c�Pg�=�J����.RK���r���j{���Kq�%,t�Q�u�k�6&��-`귝P��j���z7�aj#�[�S/�6E��/<Ź]�C����a�o~ʴ��mz[Á���i�ѡ�D�.A]� �Zܹr��$�-�]K��DK��Gp~r\���N�X�@&1,��B���4�r,r�"g��&���L�	N�DS��'>A�����w�����>Ϟ=#МH)5<�=+@5(PV�����	�U#N�.ba�L���u�d�{�3���f*���|J�|��uZ_?Z�xA�EPF��1@�wN��ΥT���')��n"�[?F~��VO�s���Y��LT���
� �tR��O~5L��&%�y�((-�.�l����r17��Jd�L݇*rr�{�y])1lr/�{1��||�rI��0 � �s�&�2�x�X�g[p��H�K���,��tt�^�f0($3��S��WN���-7�r1�� ��~���K���c��`"�f7ٌ�-�����n
��O��w��HZ���{DK�S�0�/��ө"N�.��Ż�Ho���m�.է��:0��P>g۲��P�@��7o�Pyߣ����[�{�9�Y�~d� �/ `��O,�(�a��T1�?�s��	D���\v��ŀ����P�@ݢ��s�|MO��e ^Ȣ�����/��W����}�ƥ˗��T�?�T��fL��|Oť:��8[��<��Mu�i�N�F<�d,���6}>~}�6F���>��:)P(��Ѹ40ũ�Ե�~�c�gj�?}�Xۮc
�%�!�-��f@=��������ի�>o��{�><��|���'�C�N��?����9��* V{��uˮ�P�oh�,�ͪ�;�cݵH�V��Vr�p��KZ��6���H�D�|�F�_�N}�޽s'\�v��O�U9oT�i$�2P�(I��J����6k�quzJ����,mد��s肴ɳ]�f�p#�Y%)���w����w�~���-�z!���<"�h����q�4�T�����})\��c���L� l1�0��\��,�{�.���?���>��dN�$s� �y�����h<g��A���|S�#�d۬���tF}�cُT�9��9L<��o4��0��c��$���0�!�Sz��S�����xx���1V_�u�v���[��J �V���"��N�2��e�z�Ę6���Ʒ�,M��!���q��҆����Z������sz5m�V[�.U���D~mc��9D�3[L-k�_�n�ʯ��J��? 'X��"uppnݾC�I-����(�������l5��@k�Ne%b`N��Z����q���RUjıP6)�@g����q�網��@�ntJ`�J+��^�.]�k��V�$-�>밚.XU�t��O�d<Ne��m��]����:��m5n3�e���Q���T��71sݦ�H��@��t���1;�b����ߟ|��o�mPe��U��p�3�v��Eڅ�0�t}&�%��/&��s���Ws�W���v��k(w��}�Κ;�{����T�!�S� LM���{G�c������%�B�~���\�?'Q���DU��Y���S�sV��V7�69�\{6�O�����6c��S��O�vw�=b`�T�F�o_��]�F5���b�&7�I�g�����m/j��Z����.\�@���ǧ'=)�V�:[�= ���NA�sM!)��+��@f�|�#�t�$)�8��Փ׫�hsÃqˢ�ŧ�`�w���\�����Xv�RW,��� �����sp��e*�gN/�L�fT]��(?]뜳���[�Ul�8'����2I�D<�f>�6�v,(tɬ���er��Yѥ�<�ꜵX~W�wr{7V���c�S��|�������8Ԩ�9�X2�g����U5�)����u��Q�_�8���2X8����-�$pSK�.���U�>U+ n�&���K�x}��4��.���-:S]��$-�1H��} ���$'ꮅ+�ϰ&��� &��z�֣,U[��
�����M������*P� �I����Q�6�G�x�QF����5�g�E��������t�u�G�qSN|��0m�AtX*LR(>�^"-N2�`�����\7����(o�(%��θd����������]	'��Lw������Rr<��{�]~�N|�i� 4�����c�(P�P8pS7d�_\��X����425��F�0
��V�K�Vw�g=S�W��e���~��o:4�	�C<�n ���H�u��5�W�_DGƤo�?�%�!�]�W(������s�>@A�mt夵�$96��f��Rn�cy��E@MC�WiMW�S+�#���a-/���������J�ш]W�MIl��k�=X���җ}��
��c���ݘ��تs�1��r^r��'l�=S���v���e���>�{f��1�4��L�1��%�2i_C�%�n�mJ�� ��^5�|D3�g����,�B_�t�Nű˾���mYAП�U�^
uI�?�Λ�zQ�������ǥ���4z���/��Y�}1�V��G�e�/"w��Oa`)���ʦ�j4�Y�~	�)��a.�/��De+�;�W�mZs� 4�����7y�}P�M`�&}��U�+
w��f�D׻�Y{
AT��cPk��48��mk�J"�H�ʡ�I��"�cZ	�&'ڦ1�U�������l�=���m�����ݣ�S=R��
F㌶���B���1Nu�~��c��O�=on`���2�=�Y�k��f�Z��	�j4�ax�3g��}�l]�O}�߶�(:0�3I}�����"3xP��8
��D5�z�zc��~.@'�
�t����B��ڧ����ԸV��(�Z�_��͋�!xZ����FO��l�
&����n��έ��2����ǵ���`j�iϿ�EU=s�<�T7_D?Y[���j���V�����|��m����(l`*�j�h�7�Z���*ZL=w7v�9�q�A��m�������yUK�㪃6jt�f�/�i����1 5"O,;m�����W/G:�jSoУ�!�*��۴�kL�3OX5�[M��B�6�J"�����뺱�?r���Ʈ�y�7��z��h�s?c5���_�M1o �$�_�_VO���ډQ��K�a��B�t�n*�9n?9�s���h�Z�\i���9�Յ���K��0z�x�o&Jo1�w�#�ڞ�Zmc��U\�*Q�wz��D�I��]��Zf�G�5����v�M߇q��ES%�(�b5�}j"��e���	���5^��U�]��	쁭�M8��OY���ȯ��cpˉ^!��F�����0��-��W�-��e5���>��U7�!�-:V�-�=��?��h��]�R�5*X�Ł�Yȹ�;h[T߬��Gx�l��$�U]_�n��=��G1����U���0`c�� Z�r����\������~Ζ��j�����]�9Z�GsT������]۾�_��y��������&W �G�w7�O��+B<>\��JN
�(ɺl���������vnE�J�̭vvm}N�r��+�0�X�Y��� ���eA��\%-���q��r�����x�Z=���%ɰ��-M�O��#-�X��izڱ]��V@�)��v�b3����N��x�j_O�.�������|ڍ�}e�rA������Lʕ�3��p�a���S��g��z~�r$Ϊ����0K��
#/���JT����yH�xF*��?�ǔJ�����˔�٣�$dኪR�-%y��ݿE������Y��˷L�g���:V������lY����#ъ����ci�T�H��u������s��c;�V�I�	�я%���m�t��pr�����/�����N:�a��Q�sxy�0*�ڢR35���g7��^��Y��U��j.�m�����(�b�{S�O�[���d&�&��'��&^g��\]Y|���S��L�=����s��|��y1bɶֹ�\S�����''�ou�$h��]�.˸����t�k��}=����
���M����뢽����Ϩ��1p^����U�ۖBx�G`�D�\��Q��ɫyAHV�Z'/ˢ�e�פ۩J��V��\g�	���~�H�@���v�Dw!�d�"��G�i�&���Ⱐ}
�>/,g�~j�C4M�=[H�W��E(���?�:g�{���^�>�z#����zlx�ݹd>��t��R��q�7^H�����k��~G�NQ��T�HѤ��9X$!�8���N��� g`��Upu�ȑ��i
W�!�q�a�uێBO�mi�����Db�*�8 їǃ&^���(�����S��P	���ϱ��`%�K�6��Z�f��<�^tbN!Vb�Of��X%�}�I������U�p$L���L�)k]ƴ[��'��g�H�1��&�V�_R]V9aMTC���i�|m������^���;G��ݗ�QV�"	�-v�1��At�9ްt@���PB�	ԙ/1u�r�E� �ܴ�~����D�Ui��4��Z�3�|��_�>3�*6��PH�+""����Bx��
j���x:�<֔�Z�V �;}���h͗s�����c�I􍭉�ZVş�D�Mǃ	�c�Z���K�l�����â��=3�Ef�^bL�g*p�A_���
��O4��F[�ȶ`�EG���Z�?T����ߌ3M�oC+:�@���]��/j�;{g�y�;[%&NK��U-��.\����+&��B�`	�K�O�O�Z��+.G\�|څ�'
\�����(y��U6�g���˩��4�K����y ձ��ɿt��k4�/��o��rp�S�Qi�ϵ�WRT��"��9@b�	�)Q��z. ��Jb[���DD&��YT�05��,�*^uxғ��#�0_��Z��!G�M7 э1q�2�t��I++?��/
��O� ��3�D㡞���^[L��Ts�]�E��=�}�6��O�`&�k�	���PR��{zW��|���NU@�H��UZo�E+uږ�*�	�
e�`�E��nى����a��A��Y�X�ߎh�q�cJx+"`Dl���5�P�խ��_�6Q�5�9�*i�+�e wܢ>
ㄈ��+)/ &RA.C�K�qJ��8i;�S�l�W-��i[�P��n$�]*G�6v/oDS���M"	ՠA���>��r�:>8��`??��kj���h�>pTin��ڊ񸨓����óg�������Ix��u��̍����Ҏ���Y�x�R���'ݥ�ẁ��fl �d���Z�ՃA'�$/Jҟ��h�f$�`�/D�H]:�U��[Qm��};�t8k�:TncR���	6���h��X0�ɨ���k��^���
��������3Q�Ė%����$ �ϵ�_��Z8U�T����8��G�е��OĄ��^�)��:]M�.���&��{]�~����ӣc.��r� }\%�����CA-�P&@j�g��|��J��|���z?�&d��|>s��|�I>�M~�c)�rd�*�b���жS�:w;�~�m�a�m���;�65;�6��^�
��^�w{��C�V�e�[���� Q�:�@�y�ƍp���pxpH�ڋ�T,��<�`��~�,�����X-���E_^�z>dp�	�~TS���/^�Hۦ2��V�{b�N��;���^�\�C�@P\2�te��Bx�C�L*v |3�J:��0����R�O��<��G�.T �)�P:�i~������T.�s���>d����Ho�8�^��gb!����Ȓ��y�o߅��A�d�~!�a�����{z��TA|�._
7oޤ��\��+U\cd�A~�w�އ����丘��f�tg�%���I ��ǏIt<��߽G�{�}�v~�k����t?<����j�����"����KVټ�4�(��g�.>��@`�ğ8�㓻F��jb�� /����y�Ύ��T�@oO2�\̴��A:�ٌʭ�C~��Mx��q� օTV�~f.����$\�r�\�̠��͌]����g��H��(��֣���Gl�Qu��0u��ZtcW�8w3j�'d@y~��?������H���PEx��(d ;<��"8̼
_�p%�# z&l'�P�{� a���������߻w�t�� f��DtTV]�NJEs���ׯ�O��>ND�z��"F)��ɓ'4y �Ws�p=��2h��&W0����E����������<_�u����N�\�0���<N�3����Z��p}�V�T%c2�k��?���Tei|ߘ�u����
}%
G>}�� ���q�׼ 7��֠�"Ť��� n�KUmb&�MK �?�Jt����[�*�z����_���<���ǔ\���|��޿���^�v��c΄���0�C	Z�r�"D~4{������gy�j�D��Y&#	�ݍ�Kw���U�Ko���%m[�n�T��&�P�t�Tu�Wc�=�bO'��f�p^d���?o!����Z\A�Ġg�|/"�q���]ȠN��H�Mqo	Q��os_�xAAXX�nD�0"�}ޓj���K����%�>�\������_~����_a�y�9��1��ϟ�>�/]�d�8\�d�\��zԏk1���DǩɆ�w4�����!���7���Vu�#h��Z���a�j�/�-^�~�>�U�:>|Dt���!1]�v��	��a
��T���+�a xE:$�lhL5��P����;"���m��畊,�XR^C�7˓T���Ҿ�}b�zM���I|� �w4 K�5���؄+.D���\2Zk�`n �_�5�: V�@,�eD�s�=B���F4p��tP��/(�{J�"���5�t�Y��q��V8<<�F�}�;���_~!.���؎k���h�^����S��ܽn߾MtsX����~M�\�����Z��6o�8�{
����,t�cH�Y,L�Cq�B�j�][֧+���
�n@�y�L�X��k��,�p�U��mЕ>{�T�vn޺�}u���G	hsj��Y�z��%-��2�N���*�yAӢ�ҭ��D�rS�/
H�=�%�NCU�ٛ<�<��:����`��@ \����%pwy�O2�%���oџX�MR?5���~h���J���+�y&"��W._! Ұ�N,� 7��!X
������N��
���}�V3�B$S�< ,�^'��_�sA� )��m%r���^��d �J��@1�ײ�?�Zb�'�|��5�MI$�T_��*��i_�;��-Ĥ�sab���G���o�y~����?�b��I�;s���f>�=iM��KX`5d\ã��t�m��Y6śFRK� ��nJ�c}��L#Б6���;�L�1�͘IY�ÛL�/�"_�v%���K����L�٦���W�3W����l0(�g 
��,�迿�!���j�i�2	�xD~�K�����IbjTev���/�[��y�z�?�3���l��;�3�<_$�$����e��r�z��'���!��|������&�������#epM��h�CW�U`�s��e�O������;$�R�C?�-f1`�&�,o߾	<����a"�p�Ѓ�#iE�S�����Qg�<)�dB1>]�+���^t/���T���Gp�X��5���ac#�Y>��sߡ����$.���3�~}�^�z�*����L����>�ܹK y�/���@�����?���+����l/�*g�j�y�7�bq�F������G�@[m8��� C1?�ă��B:�{��S�1�Hs�LCqMd#p>R���~�4�a3-�̏Y���^!K	 X�}JX�H�3't�9�� A�翳)/�)�L'���>�P��IK�ӝz���������fJ]d�~<�&I�-r�#��.��_)n���;cHCWJ������U�J���ɍm�L)3� >>��M�b߽�|ٽi/�.b���� �:�a�?�{Z?�j�z?T��O�H��jN��o�������$#��8�|� "yAXЊ�&<����}7�� �}��ع>�b�G� @ �k�3������I	o>�'$�-����-����	~�ӿu��(�NX`�ڿ���t���)��Wl0x��I#>7�����߶8T_͋�
���	M<"G��U<�A��(h*�m#G���$����c�C�=����sV��Aq0���C23��V��!�d�@�ǔ� [�FB�Z%���$@�Q8ݥ���:8�Բ[p�[T���rN� ��}��r�X��HtCEFѶ���ԉf��{��ۉlG��!��I��. ƍ�y�h;�: (��F�$�G�8!�b ɂm��N�@�}��ӷ�\FX&��,���)o!�������y�n�W�.*�M����AU��)�-�)���A3��O��фO��\�[����A����'��A~���T�����2��B��ɋp��
�V�Ebiv[I���c�͒��� :���3���Yl� Q`�}����B% ��ɓ��ehoܸN\(�8jLU.ĩ�*�x��ex���j�?���U}3��h�M�$�АX����^�I�m����J��G�|Q�ߦ#�E@U�:Ъ�eC��h����@۰������3��G�,����M��fW?1��3�Ry�T�X̡�j�`� �tט��[��Q�>k��0a�@V���������ﬕ$����x�����U���j-�P�I^�4l%��b�EW	�����D���@�D^r�tX.l�P�Jr��u�C2�l5`��$Kgo(���	]*|�<6���I�]"��x0w̺�VR�a��Gs�3����}>И���֘R/^�?�t��q�[�n��_}���2C�}EՁW�E���	1����W�R@�� Tp礯������⨙V�6��icnO>��N�X!�IM2o�0�Ӣ�Ԁ`F��?K47��$�h� ��_d:&���`��A��˗.S�'G���YR���_IZ#ϑ,eMg��X��g�&� ��n��|>?T����ѿ�� SpZS	�$����>�9p�'DnU�J�����?�s-2��I�7�4�b<�Ħ%w�X�Y����_&\@�����`t��I�K	$��������W��#��kWIQO��D��*���]2Q���`IG �S�o������ŋ��x�W	"�c�_��͛�X����f�cDN�֘��q�G��u�ac����W�P�����VI�=��;��J�:iu����*�x"���	T��oM����r�1S]�.^�Hn�� �~E�	�=�CsMt�<�yo���	Cm��|���|).�C���| ��--h�(8eo7�#_��Ԙ2=�"�k틚���#��"�Z=��+�jS8�*�_XLO��V�׫�-�2�t�T�X쑸 �C�pP��0�@QEY8���J8_n�%�bפ4&�h�����?�"��X�[
gј[���gU#b .+=\T�s>&b��?�B�?L�|���!\vZ��(�A��I
���ϘxSϟ=���5�ql�cd����8�J��s�y5�I'\g���?Q,��&�y6�
�,e�<�h:7�^�s��s||��Q��<�S$"�
�ɠ94���� !��ܥ��(-��H-yu�J ��TՕ�[�q��6�lvj}�S�7ש!J�����ޖ�5�˪�D�o�.+z
�f�$+y`NS���ZNE�ٶ��L�%�&���=|D k��C��_���޾��*0weLl�p����x���q. N���q����G�����}���'h�;8�j"�3Y|�O�����&������ha/S��d�p�]_�7WC�/
CRl(�0�/���%Y5�p,��T�>+>K�|[M79ɏ�A4���k�|N��.:TNn��b�B��&�~�+���u	��s�Y��]iѮ+�L����P,�
ܩ���|\G;�b�U�_[���ѷ�Yl���y'����F� ���� 0M<@��=������ �R���[���c	��ʄҡ�����y���(�lP�����ݯ���|K�xGǒ�Dߩ�����Z^XR��U��p��?+E�<e?�K����9{�/���L穡�唢å%;�26�v�� ��;�a�9ՑB]��E,���	d3Mr`��I��e7�߸>����D)�,A�fc�)Z�l�}V@5}�nW���o*bG�7"�,���T�yr�(ⷲ��=�C������8<0�6��f*��c���Մ`�0�#4�:C�/�L OP���<���x
�Q��>��D���W���'O��u6�g&j.������8�VBi%e ��p��z��a�HA����~��3���`�~����	O�F�� R?���n'.�ێ���D�?�J�wl2b.ڐKR��*q�/~�D�����C����m��p�����'"uQb�'O(�|�����WwI�C )`��r,O��E�B�5ʎ
'�6����M2����mʚr��"��L�K̰z�d̡�m�'�wɉ�;�(�+�Ke���F(���e�㨅(E��k0G�}d :��i5h��uP �8j2Pe���h&XB�G �' Ap���u�V�m#\�eZ,i2�mc�r֖�-:O���~��O9kD��Ȅ�{�=�,�#S�f�{%1���?��� D2 ���O��AD􊜋t/,���Ç<5|�~(���_2���u�����k3=f��� ��e����C�7�����a6�,�U��}K�`M�\��������^S�����{ugrǨ�в���{����I�|���[�q0���� *���eՇAW;�,hp�T��J���lU�$s]L��fUG�At��mJ�P��(@:%D-!�� _T%��J
�MY�����\o��HE9[�����\z�t��6&e�!�=}����+|
�y%w.	�����?A3`u.M���2����c^<�.�ER��/u���9U.������pO���/X����B���p�WH7z)\�z���@�a�(�)�}-])�	d��~*���f�8Tm�=w*�6�2�6�-I���E�����B�ĭ]��?b1��j�E���ͺ-ٮ� �z�  W�n�4����2��Jy �z}���;���8�1�SE��O_������f��Di�:��)bKt��O]`ba�G�R�y���P����^��O)�_b���U��Yp#P`���ỷ^� *�&~��S�G�J����U�V=�&?7ݽ��V�~�ꍽU �h�'b$@��ר?�\ɋ+\���`�k���n	u�4h_\��Mk��Zi�<&zR�Nr��٢�����GM9�J�P.-�5��{�pw�(J��$��8	H`�J*J[�B��T��{������8SuM�Q����󂸞��zO����	/]S���ϣ%�U'�\,e����[�|?~B�>��_}F�����Im�d%��$�ل�ƨ'�Z�.�s�HZ4�+�A� FJӖ9U��Y��q?�wd�� w��*
�}Q5@� ��y�P��eo�ri���^����2�A?Z��
�,P	8�����m�Qۀ�Gu�RN�}��3Ƃ���f�\�H9���M	υN�H��b�e�IA����#�k]@Ճm�.�6$)�G��e@u��Dyo�ID�g_Α��D �bi.7VA�ďNqI+��A�R�,궤uċ.�s>
 K�iߩϧD%�����K,=��9X�5'��}Ho,���G�4E����."�!�g$����Tj����V����=Қ�yA�0`��k�χ�)"Z��l�H%(5�U�>�W���~��|�·n�����RA�ЉB�  ���N�-PB��r�Gj�7���?�L��:
��0�a��4�~%�a���g�����-�O��H���q��m�٫o:Ozc��8��@eB$)��J�=h�������9�:�VTF�"��%N�T�d�~�S3����m¸��w� =��V$�hQ���΋���D�)������Z%�'~%OpҤLI��{[��k�r��$��5����t�<N�V��P9ߏ��+F���u��_��$�`�g4F-ł�L�^�R�7mf���:I���@I�ˠ���)�������� ��W.!���T��T�R ��
����o�o���R�a�=z�J���G)�+�����0����T�<^剢b&r �W_��	���\�����%D��%�0���8v�c��~��a����.�Vq�P)S�M^��cB���ف��˜��a?jɣ*ю�AW�"�4AϚ��И#�?��GK��R^ P�:)�s��kpj�R�y��t�����t��[EE{��r���&����6g�������UZt�Q!Jl����K)9��gX������Hp#b֟s�Z�@���� h�38�7���)% y$�J�b$��}����"��<����wT3����?�~��{��T�p��W�M	��>$�0M��u��ăWqx�˭dQτ(�����-A��Y�w��i&�u���$�-8����I$��>�F+A#��M�O�Z�����k1�k�^�~�C�odp�z
����Ph����ܧ�t�4��ᓭ	R��U.)�~��5����<7m�>�K4W$cWKp��La[����q��\�[D���(�a�/lL4Yƅ�c� ���W�������NY�N��4�H�R�uDB谊~�ݷ�Mp��GE��8���Wh\R(I
�mT[�������E�����O�]�ʩ
3�� �9b*c�+&�Y��B�I�s9x \&	&,�$�e��>�-�x�2{����+E�m���b��QM��׵��Z�q�1�ۀ�8�rC+��ds��J�Sw�d�@�5���+2]�>5E+��r���@�VC�Պ.ׂo����$�4�tþ��}^$�?�i(���r��N�^q��ߪ7u��ؗ�V
ߏl�nR��(�뛨�۝�@iNu{�D0�w�㤜��ߵ�m+��=��S���$�(��1�(����a�9��!�<�``G�p� �?}�}���o��e�x�.Y`����0A)�+W_��"d؅L�!G���D�5�aq���m%�~>0U�"�8�U�/��M���Gދ���*��Ze1���zo�9���y���H�ʘEaZڙHV����<�,�2�%�0�� �]l�v�ND~�<[�k�����ʁ��Dܨ�o'5>�c��NW0�w�׵A�}�)��C��ѥ��S����}EYv@d�� �d����>��	D��@��Du���k����D\�"��D�D�ą���W�]���}���0��\����?SF)��p��k\��	)P/��Zo���_��F%1q!g����+;<�q� up� ~$�=��΍�f�+���Vj�INt��&��Y���]�u�$���)��[�b)!ԇ$�PJJ���Y���m�;�X�t�j�0�y��K�� �cb����-��E��C=��[D;s�PMU����
��'d�'�(�ۦR�s��c�x*5"r[���9�/)���D���yX8!j�>�����mJ����	˵��ˇC�t� �� ���L��`�W�5ĈX}2BeМJ�Q��(�B�Ir�gR�D"��op��,��h��)�D������O4/�7��,aKb��&#��4���/葔�P�`l�po>�"�Ph���ϥ�u&���U"��0�a��?��@{�O"��D{�v��c��qց��7Z��~7�^K��8P.ָ��mg����ۢ[��X���>�/�uΒ��j�	1a���=�(��)��Ը�$vqJt^����=% "��;�I_y F�jW0ItB�H�϶%��)������K��Ԉ���(�/T/}
УDذ�Cω}|m6&�p�B@�{I�lW�T��1��ip�s� .^�㔨f���
+�\Z2����/���<�>kSfäJ��?�^�T;�k8�J�2m?{p����t�h?R�}��ʦO�mq�fI�*e�	�HtZ�H�z�(/T��
!�i�d�T��(�˾|������h��%J�+"�Y�V��#�Y�W�q���xX ��787#m��R�=�rʜS��F�������4r�H�j��<�S���H�ʼ�r*���ω�8�,��ZvB�@P��_�J��p,D}��������Jɇ���u�&jb���"�:U��p�Wҥ6��T�8���Je7{��F�S���nc��V��D�X�����ӏ�2��D=���	�������jw�T*<����r�kN��@CK���̽K���uN�!��(��.����:r0Ew���1��~��;�B-����(\�r�is��Q�D�� 4 �v/^���/SkL�o�9j�C��d�w$�E�\G~`	���Z����S��DP�#6nH_���\� ��͋���jRe�z\��'��w{� �Cb5�_�^� �Уb1�7�}��.�(�8������*���BC)�br�_ ���7�~NPX�h�� �1U�X3�R��KT�H2O�gJ
�RДh�A΢�����^9hQo�)}�B�"����]9V�ay�纋!ߩUCG�  ��x.��W�.�+-nTu֛��e�K�(VO�9�E�ZXXq�%��I�Of�o߾�?�Hw�"���3�ׂ8�g�=��z��l%�n��Nh՞͘�}�6��"�	��huH1�7�|R6�ٌ�^������I��suע�������1е@a��}Y�%��%�C�@-�A
6�b��(�d���ϝZT��>w)�����"T���ӵ<_
�C��H�8��Ą�����xu���k��Ƭu�S8*�}�&��rC��ݮ^�Ծ����e�sw�����*�=�_Ǻw���Ƣ�Q]e1h�j�B:�ӹ�8�l��c
յ��\�4;�����RJ��O�"-��'�(�E"���rQ	+������	*� ��8#YPs��$#E�@|��E9�����uQ�P�.�믿���)%:�����ұo(��$���x(t�l��+�Q! �8W�o��`q��	�#��%1��R�q.g61CY\��ҩ{�#��~��2���ۖzÊ�#g&�K�R�Q8T����!���4q�f�ЀlgR�ɬ~BY�iޖ���.��DA��d����	�}rV 1K&q;�轶=j��͍�1+�dW6����I �Pt���T�����%O�P52C.F~��[R.*�r��er%��Z̜��5�������+��1�7���ʤد����Y_ ��ף��%Nެ�����D��ǵv�b��.P�;�K�����tf*v�?wnߥm��Zb��!Yt$�#'jp�y_'o�,�a�9}a�$�V}�ơ�I�P�K�
�M?zRԍ`�a��j�������⾃�S�8#�m��CN�����pbg��md��6E���"R�8�}�t�z���a�@g�Y���Gq�O"U5�&S(���r�
��Ld{���@L_�I�=Uj!7�}�B脩P�V)8E��I>���t|�@E2y�Њ�6���0t�X:?f���R]*���E�_�@�=i�xӨL��%��bj���~x�0�.;N5G���).R�+��RJ'wjo�2h(\G/��(J�\P��ɩ�x6�T?,:K�ń��n3:�ǃ���r�h��I2��1-�3W �C�ir-�r�
�T	��ƞhE	P;�`�F����<�9�ⶲ'�ۆ#(��� g�-%K����PC�R�/)�0�ri���X�p|�o��� ��w�Wtj�U҄�R*9�^p�CM�5 ��@&��W����m¡����$�Y�LJ7A��h�6�V
:쪪�Ez��E;A����� ;��\�ٯ\��̅h{����%Q�vn�<��|Ga���|�>g�~㕊���A�5F~K�:.����?��[��	5�X��B�/Ǔ3�8���ىN�Nլ��8qv��Vs�$K}q��'iP�(�î����?+�XO�LbIe5�Db�<�apb��RU#&6նp�@���Z�(�TC�-��r	-/��T��ઞ+J��7��>��*z�>�&�V�T�Ē�@��0.�0�}�/��~��9=�e$����1ZXW��T0:h��$�����?op�mf>J�|����1E�>"��G��b���ytrL�!=$�&����{�:ʡ�-)�s�y!Db����<�y�$��uA�Q�Ч7)��b{M��3;�ǵ��Y����GU(�hAߵ��]�cR�l%�u%t��B��-�ގWZ]m��g%(AB1��S�N�Vj8Q*5�9��2a���jYH'�A���IXo֌+�C@t����5]�����2���E�p�8��v��'�z���4�{��i�����M����e�H␜�E�)�.nB�X��4x��,�,�r�t$���O������U1�j��@]fM,��T��Xh�i/p1ᬛX��6�gT��7;��Z������@��`\,sjC�h8���x����r���S��FVЇF-���T]��":��R��%��w�| �� D�7�x�s"���5c��^�ܰd���=s��"bUn�<�:~���<�X�$�+`�	����t��{'z8�z���c���K4�-%>X9��q�;,Q�A���D�`�L�MU���h���­�����C�G��Z�:��Ad5C "_<{N%�o����W�`��iE�2�]{2�#Y���t815���gTav�mX-U�(�U|�D�SR���
�)���]'��{0I֐�R9�"��k��H˹A,�K��p��VR�� M��u/b(�a>���8��Œ�Kx@���A��bT؊`���7+lb��kD�B��Dʘ����8.�ol�#�"f`��8}u��\x�犱)\QƕV�$E�"p��_o_�~)'��"!�`�>�T?� �Zo�Ҫ���:]�%7���BQ}pˋ��%�5Wf�I��b�3�b����<|� \�t�\
�A2�N�j,X��I�J_K���:�0f���q���������PT3]W"���B�����U�`�[q�B
NG��S�zTNH�2���9.��׉�M�f�e��h'&����L�в���t�HO'L��,��Ju3������=���@�l�I ,!�I��;�O�X�V.:5 v�0V#+zm����+��4�M�`�/V�R���\P�r��j��m��Dy�j�;{z9���"��^��Z�)D��Z����W_ݶv�ќM�	Ҙ~�'z��
"A�>�N�O��?'��˗�eP���$ę�1�1�y�8	E].w%q|"Z���
�CJy�0:��L������c�ӪA]n�$V�Ӣy�#g�'�g�>r�� 8���-��.����� 7�E�N�G��n��1ȭ�u��fǱ&����v$�u�z�E��.h���4��ou��1`�f`f#���$�x�+���]%K�
r�f�I�Ul7G󶔳F�-E�:ӥ|X�+U����P��tq��,��v���R!��7�1S]z6?-�*�P5j?E֪��b���oI*{�����"�L�V���������|��K�\���?�{Vs���,A���N��@ߗ�m*��n*J-)R��Dy���4R$�4�fd~6�]z,�*0M���x��3j��@y�F(�ĝ���T�>��̉D
Gݑ�с���Dm$u�4JF'���LM,N!T���������+'����3�/:U�$R-̦�8���Fǅ*pgqg-��X����IX*��w���ʴ�:��FE�t�薡�&�r��0VT����ǚ�	�� VUq90�@1�w5�:���"90��d�T$��ܙ�Yw��d����:��>\
�Q�w.�h�	�)8Vp�0h���yQ]@�x,��~F@-����aV���W�薽������1V/�D�X������&(�1���v��
uĽ#�
�x�2�{󆲏/]-%��#W�<�2����	�Fj �(�3��S�6k{`@%"_�)�4�q���DY�2��0����px���Bb���}�D0�E��iEV���7|��i���(쇬Wȫ������_�,Ɖ��DNH�o��I�)�k���J��S�jL��C��Q/���M������-�hl&�c���7�����KT�pt����D�Z�K����eࠐ���ܢ �W�^���*eg�
 ��
�`H�s���⅋���(�Vm���-��]�/�(%<E�*x{`����!(C�/��m��^}5���g��Z�{OG�R\���!� �����r�+x�8�Ku�3� D��i&��E�y�)�j�dj�n�N'J:6�dc��)?P��^�krgy���~�;�4l�ʧ )���/�
���%��n�D|�a\j2�@9my�ՋTH&C��>�`� ���}�PO��5��΄3�a!�� ��a���Dn6�V����Q�C"F}��JW7��L7dj'Jԣ�NhWY��T�cE��N�*N=������TLm)���J_t�x���<!�鈀��:�J�E\ʤkM+Uɉ���v�N?�QjŮ8�U������9�������YS]D7����`u�V�J�����u��sr��N�g�@�|H?p�\���m2��9N2p���D 1�	tMHf�lU3��T���gQ�܋J#�z*���x�D���1e�G�^��t\k:劓 ���iJ�5��vBݡ�'s~^<#R�������B���
��^T]��3���G�c =�EYk�@O���%�IA�e�����w�q�⨊�6R[A��{�;W'zS�ƒ,��+4���($,�T�4/����}W=ӣ�̌B�8�Lf�����t<� 		��f��%ȶ��J��&�T{d�?F�0�9ǋ��u��b}&�ڱű?��ױ������%����}������d�x������Pf0{G`�(��.C�A��G�*㐹4ҽqJ>*A���n��d���	�V�`�����	�(�����C�v��G�U�h��?�z �;�)b%�;W8�Z��Ľ��6������N޿dP�����jU.�.R)y���i��9��T����AG��6i��޸�M�X]O�>-��XQ���``�S<�qn*��7o��\ �,%ݧw�a�¡6���!� "�n\�A�!�p���.��·�����3T� ��:���^3���D�4����jl?��P��f��r�>k�R[O�TSs�}Db�#e�Ղ�~����Q��P�9���B���xL%�) Ȝ�;q�	� +џ������~�'qs ��t.��3+Q�ϰ4gf�y��ɦ%�Ŷ���N�h}�^��ƇI��ꝉ�Y-ۻ�o�+����U}�cZ�
`���H��B_.^�j�G����3��~H�}+�ddbF�N�	�Zp����?¯~%5��?q�F��K���M����!���u�Ë�	j��|ɺ��s�`4q��3�(=��S���l�Q.j2U��R\���K�����$�4�q�;b�cc4_��D��Y#"�T����۲$����΀۾��3x�[ݔl-�X璠�5����"��HD���3�NJ6�̫�s.{J���_�I8TY�N!�8$��ҡ���w�۷H��=�C��Z�a�ވj�}�T/��Պ�}������ ?�uo6���?�B�����3I{F���)�������ЗH��2w7τr�^_)ɬ\�Z���de]���o#���0��ء/l-�L�N[q{��:���1q��8���d@��'���Ts&f���A�
��5 ���g�u󖉄���A������O��
c��/G�N\��+-�a��Vl+$�F@u��s�3�]�U�����U7��۸�U��W?��L��A�]�p �s�������p4�����S#ゼ�d��
,AZcΖ+b@�\h�X��fK��޲>�}nSk4�v����a�ߨ�%�FV]?Z)}̺��O���)ZI��"|��4�u�~��>��Y�锤P�>鄮4W�Äo�V�;Ҍ9V� �_~&�< �{���������q&�I&���o�E��G<nZO
��ݿ?�����N�	YT?�> c���wI'��U�NP�VW*��ͭ	τ� aH�*K���TǊ~�\"a�֒.�`�Y�������O�������_�9?���|.'��{��ܔ�0�8�R�͹�vJ�F%o�>7��h���W�I�­�b�IUCEE�)9M/ߥJ�W���&���
�$A�Hb���^�|It��û��6��%��	�!�@]#$��(/ ��]�O�������g M��l��A	�����ȟJ�F.7��Qϥ
���O�������&
��e�=?��)<��bȠ���gfd�a	��MXu��4�|N�Q}בh�� !p��|���H&qY���^<�9���`�d�J��"�i1���@�ʍ�R~+��{�(c?�� � �h]�Ɔ�G�н�en�`Q~Ic���K�.�kD�	D@��o�q/�{Ρ���0���L����-���T�������0�EK�;ƂT'R���ӫ��pxȺ3)_m��(>O��t� �F�4m]k'�PMV<#�Q��d�k���2Q@���k*^+A�o�"�jp�>��0ׯ^���&q�P1A��~x�`WO,���8|qH ���_�9�RMctB6H�MM�Vsj���F��X����<��K�"�]�����D�%�D �x � �J����DR�!94� y��p3�%�,��{b�gC�}���3�u+���4�?��%D����[C�=�<2Xv��Ŀ,��e<Gt�b8��������T�Oݴ@�t�Ŝ~�m$�N�J���/�d K`t}+H}+}/X���@|�� փzVp&�}�]���L\&8x/��X��Zd���*�����ne R�4=Y�1+l��Ɍ�����ǨN8So[��:w[��`0�X�c�Jx�I"��0*H/D"�$�lP�]c���$�<~�<:`�W���Y�Z
4)
�'h��;J��8�p߿#�b=�ܼ��#����"�v�� �X3E?+B�Z�v�L�9���}ōf���X�E�E��1�?~BD�;�3A,s_�A��D�K�1_�8�`���b��{eq�����  d���A%NP���ݯXG�Ŝ��  �1a�#�z�d�ӟ��~u�V2op$]��b��� n/�� 0��������	�}������P���5�Xd~����:QZ�Q$#^�3������������Z!�k�`���P�,�-W�]�7�9�_��1��Gp�cb��6�"ƕ�a�ſ4��I��]�=�X�(y4K-32��c
l9��� ��0������;w)��8�,����cq�ӟ�#��|�[2��[���'�����V/�z��T��[�]���jrNhјxM��Ǉw�6FUٌ�bT�9<�[px�TS��T�LA\�^���#���Q9�Fyb���2����_�
`y,�s�;��2� O�2�{�����[�'�<P! �>�cp���|����@-���=��5�4��D|sBqSB���3B��q'd 8�q稥�\[��TJ_���)~�1b^M�H�ء.@ZW.���[�I��%�`M�RAdW�Z2�a���E 
]�0�c�!Xq�8�ܴ�T�eM�Eq!�8m�r}1���7Q�)[�S%��~5$���i(Z��N�;�շN���,p��NA�; '	���3�����W����X����b�5��Ot�D�?�J��/JT=����S���(OF�yyw�~3��+hIxbnSd���P\��$Nz��M�'�+B����Շ����'R����J�VR�ㅼ���)|�.KI�9����V�_�!�f�)�a�{a�s�6)tO��#h��譄�B�@M\c�-`�3�QT��O���q���I_q)��Cu�:(�o������\L����ܦT�"_o��*s��NR4P|W=%�n%�����S �;��� %��й�<�mx+@���T�HD?u:or��_��NݕF���I�
�)E�-?bq�bn���V�V(ã>��Dq���h�%�����J��\+�K�td�w�y��L ��v�����/�鳧��Y���!�tG��䜒�Y�7���)/�����2��\��Y�/�MZ-`�l�Z
:DX"1�A��nߺ���Lhz�p` 'r��ۏ)V�D�qa�8������:��^$q[6 :D�����{rB�D��� I\`����lA�^+�ҋ'���'����WA�G�c��I�!Vc�8q?�`��vp�j`ڧlAd�SR��>���J�pe��"�>���'.��m$ �����{����%����
|��i��
ԍ"����L�����}�s����Rӈ��K"�P�w�K*�WjO��mHpI¡6��|Fa�"]g^��aR�<id��{�zh�.�Z-	
��W�FU�F����Ę/��Xh�L�a��~C�j�l�����K�cK퇻��:V�x���c0B!&�T}e�ۧ��*��\Vz��SB��/I�F*�!��M-�:X�R\�����U�i�@��\R�U �
�%�I˓d)�����?�՛Z,9 �S�Mh�87Rl�8U	p�_JZ���	���9rI�%l
xoF|00���F�,q ��Cc����صʪ.TM�H2����97��J�XX:IC��Qj�}�#x�1jo{ٖ����0�S<�Hs��&EQ��X���To�fҹ���dqo�;b��B�����_�xBRc��B��o�rN�w0��n��� �42����o8{���+��E�S���0��6Ki&�A<X-?yL�������r]�8��=�D7GJ�N&8�tM��Du��9a��/�C�D�/�gb�R� �|�	e���"���S�|�B�:��Z����R�&��*Rb&�j�3��j�1 sJh"!�b����alR�b���\�z��"��\ ��g�Rғ��Z;�~�~Sq��{c2�0&!��+>�N�A:kxQL�`�3���?uL�y):�3N��0�|ڒʈ�ԺQI��ʤ�K� �D+� ����C-�)����_��
���oo�0�KjK� I䊇œ��_� �;�O0	`0�ozFz�%��L
�oaWm{���YjH�׬��>Q�R�P�&����H$Vkl�-|��[��`0�$4'%;>/_<'Q�&��X�|�-qa ���٭�L�~T����U�ZJE�?\�2v"� t�~Š2�1�*�����Mp��u�Y}�~���\����"BG3��oݾE�DAOW����.�g��R%����{G�%�UER��ڼ��~��������~߸۶lI���Y��� 8DV�VѤdϝt�EV�8 ,���.%��>!g��uSx�V��~zc)�s�oq6:F��׬���q�g�x60�BV4W];4�b5Wg0[<g��^�a��&��|'���1�����ߣaɴQ#���j$��f�|��C����xt�R6�A7b��{ɹ?r�ݻ���+$���+�����Y0q��#��3=\��e|�n
�1�r��=��+�Cv�X6�U+�tV���j���Cl*3�I� �մ���z�'�����ʘ�3���ZV�T�Ȯ5�IB5�Yu ,z���X���'�;����_9[`�p)F�������%)���}dt�A�f��3_v��RB�h�����w0��U|,��*� ���F(�sI�u�����[wn'%_Qs�aW)�Yd [Ӿr�P5���H��*��h �}�7.hU���M��
gYi^eh>�j�M?����:Pڿ���2�PQ�����8����%�����J(�32^&w���;|�u"7i���ϛ>ϵP���
�?-{I?�6r�*6R>��=��_w>���0K	c;����*�)z�=�QG$���/�ڂV
͒I's�mFE}���E�.Dp�������ü�
�=��n�am������M��{�����GN;[5�2���B����-���S����0X�vS�I�V�\�f:
�β�+H�cQ��i̍�a1W,p�deϡ[%���+g�S/�x�L�J�����O�j�Z������0��Y��M����Lo�G�� ���t�R�^whs�88<��4�1��_�k��@���tx4��i�Õoz��)��O' 0\8��ДwD���ǳ �i �E�QG��!�A��5�?0��k��+&67*����k��;��$qh��x�Y=g�9x+���n����9>4ݔ���>F��M�n����6�e�9�3*�߁�k�8�fF�Cj�*ʘ#�;Λ er,L�?B�#x����\���/]Lׯ\MW����/_KYih��P�t<,w´SD��/�a�
9���v�1�p�,�Β�cm���㐣����P�y������N��%z�nɅa8Ii��쿇�wZ�N:�i�Z�U˙�~�RL�s�*�N����h�E���>���߯UPU�nY��������/丠-Փ�T�LM���$���g2�5�5{A<�?�Q��BWxL��7�l8Y�Z�N���P�E�u�%DM���ʊ�i���8(��G�}f�%��sR�x+��X{F�b�*(F�j��1O�
ܨ�u�模w��{�x������l����̴e�@w���eg�#皒��R���?}��\�>N���:.[��(g��Y ����Xh��R��g���5�2! �1�z���=[*�8ą��"jB�zX4�����@��"��ϟ�&(�	n��F�h�2%�����-à�-u�/Y��R�׬x�H-�a��i�e�x����Oq����yY-m��^\pRY�"{Y-=�7���Z��<�#4r ܚ�=�"����c�Pɯ�(Q�2��g�8��#R������V>�6%��R,�i�����2�I�M�R��RcJ�r^mbi�dO~o�R�ǰI�&���uu��$H�q��������-:�����fpQX��y�Vb?AM���sq��Y��Fl�=%�^J�:2J���'H`a��IJ�'���5�aӮ��čB��<K�ǉT��	��x��	�P��ug|0�� ��F����wn��-�Q�%������������Z(�؀����J�}�␠���>�� TA��#�0}�����-�M����Qw����/�m3�X�;7<��|cwe�t����Z�F٢�2e"ĶiצsS��N��i[��ʎ?vx)��f
���G�l
��x�#�	�3
�{d�c���g+[��-dl/7�~������^�MG�7�U�;����z�X������gJ�Io@'d��ci�^9��n:��6s����cx�NA-K�k����Ɔj`f���h�G�+)�H�U�U���˗U�J/��r��& �]�"�YbU*,�����8�7}5�?쀣�%�5g�c0��B�������f���)oǘ�g�Q��Ń�W�$i*�9	-dF4��0M��+�A%�	�wz�����*U�sJ�S���搚9�f��{��1�`:� L�ǔw�@5�ʸj��fsvJ�r�®���!T�3��۴	!th�:R�ws�-���N.n���b�@�.Wi<�
J��fc�i���C�P�q�ڍt��5	��ֹk�T�4!C�{�z��+E0�a�7o��y�Ze_�3�������<ix�Dll�Iǘ�ĈN@���MY��l�BH$?�IIR1m�@��G�M�^<%�F�Q��2�r�zX �	|���M�eҼ�]����j8�T0lM�m:m��>dW�e>/lA�#��M�Ks(��i:������؁�!) ����Q�9���F8g��C#^f���Z)➇ٞfޥ��Bl$��������5�?��?�ݻ�$��t6�������.�K��D
�?���<~,d8Hxx虊�H�X�����F��`��v�$~5���>p���n�-�����"P��D�D����q�t����)��������2O�q�i�� sRja>�u"������S+��	n�o��N���w��D� ��5g&Ou���q��z�'-�WMK�2H�G�����m��
I���/��/��N���y�2h΢觠#��,�,sy,��ת��˔�n����?+#�.�ijh�T@�zE9pE3U�#��)�\	�q��RA��B��@�B[ݱJ��O9�����MB��(�����Y��vQR�KV�t*�}�$� I�R��3[���<��-�y�A/�C׼�(
_�#���K�(�TC3����)��c���rjp�"�U�
G+�$Yk��B�����~+�������sp�B��!Z���2I-����#[Li68#��M��Z6	��[����Ѧ<p�����[K�H굇��M�7')��h�� �<4�)]b�j1��=+ H�������ο�����g}�m�;��V�c�B�	S�u\�ٵ��j�� ��B��*(4=�Q�)��]k��l�0�7	�s�T�<A���7K6#�	���'O�� ,@��޸Nq>���VS_�.Ꝗ�~�>l#�Eg�$��+3K��!<y�&������F�ϖ\h]�������a8⚈	 ��T������2��0	rp+!�I�����i�m���5�k�����G�
9��+���0YU���+Z�zy(�R���%P��Z�6jETٰg�͝R]���G����ݟTVd�[%Mɲ�"�S�$�3�&�Q=�	��UԢi�FC6D|p�N�2������Ҁ���?�xc/x$!-G�I"q|�(�w��myo�M�}�i.�kK4)�G��dcY@�%��A�-+ьg9cb�zK�{Jۄ��;2G���M���X.��_[�w��S!�r���_���j�9y�
��P%�H�gn1���.em�q��W_K���'τn��۱��]%g��7d<���:,'���}�k�0*@�������(P���ݫQk�k��KP�~N|F�Ӛ�8i�㌛[�ڱ��
�$�`�.�QR��G��ɽ�t����4�\��(_�&Ę�.d+��L�_`�Õ�QC;}Z�(�ZPl�L^����U���o�I���R΅D)������_�@$�f��H^Ѵ��	)|���̞U�f�CŴ�iO����}����[�'�������{�;�fI̪+��xz)�Gpȸ��L�.:�4Fl�����j�R~_I�0�ף���L~�u�
ԯD�.��r���g�8h�X�FQ��/�G�M`r�u���]�v]1�2���z��
�3��p��ɓ�I�'�7��&4�4TmD�g�z ���Q�@Ǭ%�gVMс�`�g/�[�փ�𚉖�o3~��~�2nr	�����lae���1�II!;�c��8��,���&l����]MPʻle�w-�d�"R��*Ʃ��\,���Ke��&|q��Χ����R�	��Q4��pU�=�>���H�i��}��Lˑ�s7�̬� ��P �F�6����p':P۽�Vx�tF�����)J�!�[�Cn$'!++�5����-���m���):��)��O�0+�>� ��`i���~#5���@jp�v?\����%�/��*X��ѝ:�ׯ]���}�>��@�Ii#4H@9q%�?%�I���~������y�UC}o�$nײ)�����s���P)l��9O7%����&�z�<=ML�j����<���M��M��K��!�WE?�X��It�m�;/�{�MRzKSXP
Ǚ�9�~!�{������g�vH�j?f�3�e��;��4�z ЊY!���=���Xn�� ԌGL����i���Nb�`�G�^�_W�����d�c��8�XZ�pc,3��]lr� d4�H�Ki=�s#Qa�8	�����G0Q��r�Cˀ��B�'n��ɿ��m�FKheT�S���K��a�t�n�U�p��M0㑉�zh��@�	�+ -��@�Ar�B%.0�Y ����]�|�wp,����KWd��$C�Fc�b	*:3��k��T��!��:��OJ�g�Y�`���g�O����9����O�}�	�p	#A��m�M!{��^�Y꭫�Y��Ġ�״Cm�z�?\T���bĕZd���$�j�9���@N3SD[�U�0�p��L<2�w��:�ciB;>_J2[(�(8	=x(%~���	\Lrh�0�P$�)0+)�b�>��!%�M�Xh9���p2��;ڦP�0���*P�K��A�炀Ƌ�k��c0bk�pB�g�>�z���1�_>���W:\�&�G�$��fO�:��pn����F�|��WŁ�7"،��� \Q��ʪX�X���7��J�H׮^������:,m^�.\�|XS0���s~�XY,2���"Gf��R�iD��s�����L&X����`Z�n��g��&Z
[�-v���q��h"Ɗkn�K���W�?�1� E9FY�Hj8���N�Ѵ'j�q�nm_�<b�8�V	�!%�W�'U� �2�'�=��P�yӆq����B�)5S��E\߮�Ok���o�J���?E�"#
�
5�K.Zg)Zd�,��f������Ŗ�)����i�\�r4G�hCGK��j��~f��c�k����ګ.�?������ڦ���,8b�tnъ��VJ?�tW�Ik�鹘��s�źcm+Nr�U� ��~	����K���`QLh��{������6�M@׉>kfZ�����SO'3g����q�m>o2��㹆*��7�g�p�mX�{~��0?���F�X.���^/�p�V-�,�ì=�5٨-Z"�Ԍ�0��@E�Lt8 X._ޗ�;��(p��;E(��<��W�D;�B�h���IB� L�;kC£����ߊ'f��@��BJ�=m����0�#b׫a��2hy���(�L��ʰ�x�h����!PǕs��v��H�y�n�5�a���bS!�?*�r��N�oq��lo�x�ŦNO'$]�{�A�Gxu1~�?͚�P�*��eK�s0�A��]��a���7c,0�p,��8884%jaT}:wD0�
��>E�ߔ�����"�/^�:R�Y��>��M��ٔ��Qu��B��?�5z�Q h�KR���V�O��gr��`�A��]'l^A20$	�Gk�3�����Q�*�I�>i�X�x-�#��{�@RB�%�_Y�o����tD'�i1���H)}�~��*�)�X�0y���;��v������l�3Yd���`״I�C!�u�޹9�Tƕ��]��Ls��ll�;����±f�s��TE�s^�B���e����v�.�+:}'�G)������2�Q
�mx�`ަ�K*砖���ٯ�`:w���G�� @�"u�6u$��whP�6�g����Q�3u�
Q8��܏:UדV��1��΋����Tn����f�3��-��y׍i_�y�-3���üs�Jw�x����26��Tɴ���-ޚ�d����	��N�b�0؎w E]n�:�"nJ�K�哛���D�ZQ��ǿ���yIqO�>�m':�p�������>x��<y"�?��,�?K���B��p�]+�&aO��Mj�d�j�4ŵ$���Ę�D60P�C_OM ��el�T
Osč�pĒ~��S�;��%��A	�!��k���P��O�Ov���`��C[��+��s���,js��/�l|��%`�h��!�Wu�~f�$4+�������h�0/����(P�86�A���Y1H�j��w>��L5�|�]�z3�Ï�&� 8Ҳ�D ���U�:C)�y	:'��"���-.��4��s��)��[��:�(P/J)�]��vqI�{���=#�V!ي�y\j0O�MW5�G����bE�K.�+�l(%]'#��K�S�ٲ��"�ӏ?���	
MA���{@�a�7_�nߺ-Z�6�cc(��,����V�<�cmʘ����%<[�er��9�~�CK7�+��\ʹ�U�6�%5�S�㦉ϳ���X�t����P�㜃PaC���_[걯�:�ÿ�MZ)�BXb�'�P�?�8u3���9ax�`��MR
O�0ƸA@jl7B���.5^B^�e6w�VF�0����G�M��Cg��~�1��cZar�h9%LX��M�,�%��Uc�_u���_M9m��"t�x�
�\R3���>�`w�\�i������v}�[� �ϒ�ࡘ`(��ة��/��9w�3̙[��Ջ�|������$4E����D3ŏP�	�E�Ф����0��KMW�dh.�x��f�<� @��j���4dj��"�,f{}4�)5|h��I�
�Yg���H�@t���18�'l���~�-��@�]cN͜���y��h�k�{{��ˌ������}`e�A�[�N��@�H"h��&��P6\\]�G6��ӯ�~����k,1�G�s����g�d�*ԑ��?�QM�����0Eh�i���t.4�_���tW������{�fr�����+H=R�U��5�df!oM\�O��5�'z�Lg�����oH <���QwTh���$��۵2�1�<��0�f.7�d�$�ڠ�C��j����&&��.^��+��l5w�����4B�`!@��A�~�}��=%��ZC`V�19'�K2(�6Dj3��Ա��S������Ov�W��`l����\�����<��˞V��4p�'�PF�g��fs���~,|�HsrB���,�`?���ƼA�n	���#�fjZY��h�$����}]l���X��r\�@�c`�`sݳJ�d��=4��gq�Bb�޸~��~U�%�b�x8����gqd�
���;w��cOxs�)�q4�q���Y75j�n�R�� �P�p_����)�B#��>��?f�8�k�H�gv,j���Y�s��{��Z�b�?���H�����)�^��.rgT5�_�	�����)��!��ф�C��Z�__��u�
SU�NX4��������W[f��W��3�97'd1�G̈�j�^&�8\VM� �|�.΋�/�%�~r��2Ύ����;&�:,	��b���d��a��Ӑ�К괿�N�t\�Թ� �l���p�j޽e赥���J���:� `��` >cq�#)e�^�Ï8�����+���#e����?�J	�C�/ugw!a{3ې1���bӼz�����6�l���\_����æ�9J��i)�P5���u֧U��=Y��UQb!���Ԗ_�q�E͘�^���{�{��5�N=�X�Y��ʸW,�em����]ٿ���L��4�<�
�#�H�{F�=ާgϟWa�D����3��Ki��7��, z��zk��O�>�f�C�`���ʑ�����!������
d�'�VFlb���ciy߸�0�l+uvH���0�U�&3�G_"����.&?��&�d��y�M�Ñ�%ơ=�M��ʐ�|�&��u�m��d�EPt�i���8��8��M�U��l�"r%�n�����k�G��{���טgBJt��GÝ���&kۈi�{/>�b��S�[��!h��_<7V�ך@b0Zm�UHh8G,��6P%J��~�Yg*P����b�`~�:h)r��Z� ��s0�$&'���311F�
+���\VV"8�"�Lv��;!���&����L�	Zu���1P�^<V�e>����uǼ��g"�`�H��W� L�g�����`U��['���(�1z��dNd�'N�U��V��G�ՋWR�g�8_�h6�P�
��
S�.�r��`�/�?�l���=Gk*f~�&��;w��ݬ��H��h������GKR�Y�s��Lܚ�L<sR�Y����{���>|eq��0�/]�)z�,��^}���s�K?�ZB�9�7j��;�B=i$iIbcK��;7��̏�S���ͺ4�}�C~|BԆ7�]�������m�0�2�:_ذ�Sv��j-\���F̜�X��V١��q��{H�:�,�ml��a-@5�Z����H�.��z&���woe����z�M��`6߂B<&X�2�?�`��z��(����N�ח�6 �.�U�HL�&��� �l1,4h~0&!xP���	)Z���UbEp,�uGf��]��]=O�3\�5���s�Q�N׮_K������￯�Ӂh�R޸NV@���]���b7]�T5�K��e^N�z���dY�%"Ӄ_���ߗ�Q���;�L��C�`�~V�	�c�`G�AdA��5��� ~�*�͠%B�ޫf>��nߺ����z$��Hj���n���E�H�r�Zk�3etF���oG2�TCD�6pց�zy�5��Y � ����Bɶ��X.EP���o�ԫ��o�/x�nf_|�U5��9Ɯsɕ)I��z���hu5�|'��9qf�X���|�����7��3��	��>
4QS�y�gY��t Yt�*ԮݸZ��-I�x+!yi̮!ʼ�:�l�����`�-ϾX�1e�|V�zb����.��]q<=��?�0� x��V��RB��@(}Avє�Aփ��I���[�nF�Ow|�T�pB�S�i���}�d����]1eׄ��X���r�؄6Y�A�OZ{rg������Q0c� <�Y�<�o޽�Ҹ��D`���䙤v޹}'ݹ{G�|�_B8b��N,]�$8���˃RC�D��>�x��^��n߹%B�Β=b������+�;����#�0�!� d���>cB�dӲ�[Y6��C����y3��� 4�s!�Z%	�E���?�����.w�M�\�0tq����0�|�gYhR��PY�`�"�k���+���a�5ee����Kt8�כ��Mן~y��? /�Q(Mk4�{aJ+�8g�3OW���q^J?~��W2�Dq��G�il\�3�j��Ν;:�H��%��T��)�*a�0-]-F�XKu=$%>�p=�H�mIy��5�1�=u���)��z�'"�&^Xl �'D3��v0�[m�B�lp���E���xA��oAb�ih���\A ����b>�v"���I.&0ǥ�������|�B�W�Tv�-���%���e��eK%�� ��UP��Y&pX���,�^C��=�Ak�E���:L{�}�
���U�W�A�)8����XL~��`�V�W�"���[|������Ǝ>$�
���"9bh�FY\�X�r���qh!B'ǟ�x�?3C�����dEZJf!lb�q@ bIrG�����j�����@�{����y�g���]��0.�U$⤮�K9������3q�NTn�����G�9��3�����M�ib���r��j�����$�+K�-�c�Dsڤ�d�ɍ�X��^�~��
�גƉ���A�"c�ƅ��(f�M�U�@��Ź�$���������O��k��c� ����~������Cqj7=�����b�"���]3�c�Z
��Q�GHk�o^�y-׃��{sY ��|��	95��PA����������/h�O��8� p��n�N�}����4X⊍s`��"����x�Դ�d����Қ��"�7ٟ�ҟؤ�uW�{d*�>Zj����GI#.�s!D�8GEt:�!� �N��\��t�����!u��l�W�W9���?�@����n�)$'���V{o� zG��h��Ip����eؐ�K[l�+WA���%=��az\M�w��o8L8��zY�E����y%��+����E��[������7��;����?D# D�WZI/��IrAV*h�0���8�ќc�$Rb�Y��J�F=��Z	�ܱ0p���&�I1���D�����|��1 ��p����qcZJy�#u�9ś`��}�o\Ow놂�ܓ�\dy_�������3��&��ZHU�X��'[�/Oj�ʹ}v
�ln,
3�~�^����L�͎7�D�ږ D=�DA�yr-NC
=	�$}�x;��0
�i��,�2��V�'w�e6�3>>�@uAy�ˎs�I�F�i�v��E��kY�'B�����s6(|ɒ%��2u��/�ᚈ �=4�*T��y�N���Y]�Y-&MQV{`�z����5�;9�Q��?��?��><+�gox�����d����V;}%��UH.Ŭ��й8�>�\iv� B�L?y�Q1k+,zPR�I��`6XM�Ɖ	m,ڍ��Ç*�DM�  @�����kt�w��M_~񥰷C��!����5���o�����k1�S�z*a�9��Lk<m8��=��J���p��]R�T¨Bi�(�M�.X��/-�1�1�����(a���lU9���x�!�ֳ�pd�����F��8-��i4Ԭq��O�)l��05��&��(P��S`��&�����5�m���X�衱�C�I&�k{`Z߸v#��_ߋ)�4Th�B��z; �w��L@l/_�pHB&᪚�R���ś7�7�~#���
�m�vBAB_@�W�!�,1���0�!� �!pᜒ8NI�\y����0��|E[�z�YcM���^� }	��u3�^ūo�7 �[����sq��7*�r3ea�R���-&���u�	�����:����ֶ�t�M�h�V��xl�V���E5�1���in�jՊ�)s?)�|`�l���>_"�;��h>�X�������j6���0��j��i���
��{�_.lj�c3vZ&���߽�
���i��N0&W艹f^�;&N՟���W�RGf	;	7U`}!���Ѕ�A�pX��G�2�`2-y]*i��52�eެ��� �}��i��VE��ƥ�_�!y0��K1�/]�SzoG��W��shaVKK?ݱ4�,���LP-ĉ��]q04Sx��6���9�9 ����17ě�1����ژ�L�2��ʰ@��p��X��1*�&��U-uF4�q������Ι8��=Ne�����F	���aR��J�D�q�Z�|Y��O
/
.
�lغ?WM;f6N��<�ب��l��s�!�5����2+r�-C߳
�S���П9>�S*�������=]�_��[-�����~7�x�i:��c@C��ʌ	j�Bh�/�x���~�(�ǟ&�ޏ�1ߓ<�V��,�"�l3
�ݻ{OIF,f�0� �/��)�V�vBcE,b�s@1Ghtv-����D�gi�AԿ���g3�Z�>� S[��>'��.>���G*"���
H0�Z�@t�l��pH�E���}.x)��X6��^�K-�(�Hh$�bT�T5��ZY�a>����ƹ����s����q&����"��'*p�Iǐ���H��(��2�r�=�\*4@�H�|$1��L`���������+��]���0J�fˮ���:�>(#�*y�e,��Z�=��m&�WJ��NC��=ۛt�/���l��wr��b��̴Q�]�|Qr�>C��+��I�X���͛��)j��C3�W�(����X�'���Ȭ��\ 6{�\Ⴐ"�:�)g�2�q�ʃQ�����z�����X��:蚩>rg�\����S�%_�6����0*@`��;��i���B�Ҝ�Z2�_�� �.U�����$MS]߯}������':�����:�m�N,��g0�KgD�}���f}jk���)���:�~��$׎�
P۬�a�]c�z�w�4�by�hm�;���N�~�:i2�8�(�rZ����:QX3�u�Z,�� ���M^�61ΰS�d(�����k�fx@�b�\`�����,�N@kՌ��A�4��'�J�j���p-J Y��*�3i^q�:>mݕ]d�"�F��X�
'���0����hP1��jƇ��?Z����N�"�m\�D����8�~;:�eMi��f�fFm�lme?u
C���$���V���"��M�M�I�W�27�VR�41OAE��m͊]�Vݹ;���`Bx��a�	PMi������w�8M���Ͳf��Q���Zdw�$TsnZjbg6�+.~�V���'2 ��P��2x��CR��"HYK��Aj1)����Q�,D��b�?�|�J�W�+�)����,������;���#�y�@��$�$�Soּ��0"`
/�<(��(��ʲ_f!dep�#��24[�:�,��"�-���`��Q�hԁ�UPc0Lve�nE����n���� � ޵n]�!��CU�pF��W������IT�6�-�M��i�y�"d��_L�侊��u��&iO���t��5��N�Lp^ͨ����?#F��*iNNFT�'� %��ʨgu�]	�J#SU�)<��-�$-���N��A��Z���*V���.n�����t����8$�a��h(�v;�,څ���k�I��$eP�ՑYnbΈY�4)j�Z�~��9��z�	%vg��7��L$Nŀ�<1Yv�V�,7L���LۭM�#�S?'�DP��a�ʘ�Zx����k>���~@}3�>-�G�z՗�f)�S=�����5<l`��(���}�w���IװƱ��2����i;aɟM�y�N��8��g85*-L�RZ�/[o3ü��H��'��b�U�Q�A�i^L0.,�~4\4^3�K���  S�k+S���{m��v��L!�g�&�3j����t�ٖ@�R��h����D�����ꔝ(�y�m}R#Ӆ�va�NS/�����z�wơ��=#�2?qB{G�K�y�ڔ�(��
6�*�X\�!e�`6׀
!h�M��q��^����_ � �f�����6�-wPLfr0�p�Z
�?%Ιql��F�O����o�P�Q�{h�c�&��&`�s͕�T4a�]��z0�O�3�s����w֮a*&�-�L��1���y�:ޅkf5j0b��e���_�­/���{&�4%��E�&P��J�{t��1O���2��=���^:��`��?��V�'�Pه[M��Bj��nM�� $��pSϝ���q�Hr�kKa�ۯ����$�H�K#w���-y�"j�]�&ro�f���V��I�e����'r�	�_��p�I�Y6ez~�m���g��X��ht��.Ϝ5�q,��{v���X�h�ك�R�c,rL,YZ�����>���fz�ƾTI�N��.����K�`�D��f51d�ֈnP���X�K5X�i�_�:���E*�Z����������s�';�;Wj����N�(����S:�1�`c�;�6�G�{�F�f�&j��1�⚑�N5���F6�ډ��/�����&�*:$U�Δ'��-��0�8�~Ӧѷ���L
�:ng�WN>b��`UsW��)|0�8]�f=��.�fOꈖJܼ��͖sQ�,cM[���6���K�������w(��1�=���16�=��1�I0����!�1�7xP#�>K�\)�Bu0���x|B�:�NrX�&ͣx�F��Vj�&��v��5g�����;J6Am/�����ő����,��|g�G�m�6JQ�3���R�>Sش�������k����2{>��~/�+��Z\6�M>�Q���Q���U��|b!���~]鼢�q׶|�f� ���ZC2�� �ti�C ���M�vs����{���J	�dC��,7���*������55�lʫ��\o~L!0b��ߦ�#�2C���w|2�J荇�R�IᜢN�o6;�/}�C���k�ײL��w��co
�	�S[��^�{���L-l]�C�Ѳj�N���Ԏ����0��̜�3͜}~uh���D�}7�I������i�8���־؞ܵ��H����:.Tد)!��"*�%�	22A�!�&��y����%�۸d�ćB\���9(1M�M�Yo���q`�J��䊙���l�sd�ny�f<̊����{���m�m�v	N�.�>Z���;���7�9YQ^R�[ω'�ߍ�����l�8M�Eۅ��}J���\jl:)�v�V��ǣJ*S/g��g��qǚf9�EY�(HHG��2+��w�[K�0��@�l�,XWE;�c���J����l��߈�*�"	�����C��;剛2U�A޳궹W2���&<c�����`��dLV+KT�2ވqf�b�b~��ϛ�4$����J/KR�S������&Ȥ��)���������&?��������;�:F���)/�}�QC��K}�tS��&��ѡa�E�`ݔ��4%3hg�T�.���b�l�pL���~'[�b^cK俓LՍ�RG��]cg��)�Ԅhg��!L;K~V;��+�����$���3b��Z&�>l�QR�N���LB�+�d�!�q��#��P�9%i�$Fؼ�y�ɴQ�� �Ӿ����kZ�b�Bzs�^cw�~������f;M�7���~j�!������2�	Tj5퓍&wIs�nz��4���&n=�_�m�ꎟܻ��"�lh.�f��*��5�7.�Ιb}�ߏ�4,�=v!X�SN�����ф�.�4��'2��Uq���k^v��@�������w�peXAg����~����5V���l^�8�M˒�YV���ۿ����py_��f�'��埕�L��/��l�N�\.�)���f<!�h!\�3���К�,Hǡ��Y�o�.���m������Ã���U������'bC�A�RgN-C�������f��"e�Q(g�����&�\t���TM�5��ؕ`b�1
��1v�6s�K���ʉ0bN��%vy�G�k<��P�4mś�~��{�_:�`f���%��Ǽ���k'P����o�H5���������*��W����l��,��O�c�p�F����К]`��q���ܨ?��l5��IL�a����<-�����Tq@�X��B�1����8 �}p�*��zdｨ����G��/���P�m�]�� G���
�5)�^�8va�W<�RU�T�IL0�^eh�L�T Bc�e�S���'&�0����9��~�-�;��w�(Z�RV^�q03M��qB<�<�:$(z��qC�[銈m���Z�h3�ᴻ�����Yk+n�ӑ@KG=�v�0BÛ�%{��*b:�Q�W�g����ɿ�$i�d� �f��S�����+R�z�TV��Uo��U�L�����62��&!H����I�=X-�	�h�S�C�{�>`�����ϟ�H?��c���ߥ(��؂6��E�">���P<�M!���&����y�(v^���υ8�j-��t95r�'��X �A8�&��{{{��w6��q�5j�����SmF4��o�9(������w����qV�s��aG�)&(آ ,���lLAӶ�pO�0ul�4��`��CLA{r�����xm�7��Eq+b��F6"�S�u�W0�Y̧��m �[�������1e6����٠R�M�y���w�m�Y���C){�
�/��J� ��_]���bv*-����9��&���I
�`#Y��n��H�δ1@?Hs�\.�m��؟�]��+#���~����ÿ�]W�2R��ϟɜ|�����v�:g�g�q��
��2�����m�N���v�"/�)�_XoR:��?��H<O6��C�L���8�V�JOv�L���$�YH��3�UUU2+Ⱦ0�9C�|��ڑ�þ(�,Fi�O�p>-����~<���u��˚���(+u������Fw$_>� aP��/z��N�Tt ��i��;���uA:����q1��j )�"YI$7��*b��B+�t���ى~�ju��2%
��[���<pv��Eud� h$-�>���.�s���+#��B����a5c�	o,�U�	BKE�&�i�=��%<!������|���ψ3#�_�z�x�G>t��?6Z��fV�Ok���R��ѣ*��X|�XV�Łs�5C�ីӅ��B��U��:WQN\�SU�ʤ�v�D)�a`��-"�qS�6�9�	[�������M ?P>Ƌ���B�Z�b�}���ˮ���3ժ>n ���H��W���m�ݳ�����Q�oi	Q��b�Z���&�H�V�iw�+��3A�3��MH��&�iO�4�&({���b���ga2jg֓'Zh&���1&����[�{!}��w�̺��J�͙kd��[�5_T6�v��������`��sF�#��A�ᅛ�0くA�٫�p��D!<�s����(d$4Ch-tj3��ʨG&tD��+�:����#���L_5�GL�"��Iۄ��~ϺP�Z�.#&����X�+�hj4�"�a��(�\�<���y��*�]`[U5O!  `6���]}�����=��ϒM�΁K ���Ȯ��d�n
��y�K/Hd��^�CÄ6�yۦ�b�?߿_��j�ߦ�>�%�`P� ss���'���G���m���[�"xv�VVkhge�Y����Ê�q�γ��c���H"�UC8::�~��<�\�gl>x�r��0��ԱAM��H�l\��cw
NUխl!!,M���)l�vN��8C��Q˜���	��?k��b��hL8yV����d�"8L��/��nE�i�1�;���b�� ����^�v#ݸ~S�l�!0�I�9��ɭ�U�R�-�PZ��`|�♘�X��H.�]jAؘFub����,�������LG�8�Դ��s��u^\�����ݢ/_<�&$�O��͛7���:ai�ϴ"j6B�2Hi践��xR;�#�� �J@k=��܇ڐ���Lnct
�4S*�q�>t��@����s ��g�L�5�f\-�}�c=^V3  ��IDAT!C�`�d�k���я��qГNn/�R�CC����m�"�/��&}�ͷR%�1�q�S,���~+N���f�3S��F6N�V�h����Aύ}�t�����V�֠W���F)�K���?~R��t�
Z��.2�χ���kL8D8�[�y�	�ꔊ���c�S��bh_��頶���{6'�&[*�S�f;���lԌ���pX�EB"��������٠A�#+1���I"��g;?L=hy��,m�%��;�ơ�B�������h�h��-��}��1��}���Â�V��ѯ��_�Q��i��d��h]�W�^��f�WGJ�Xt��9pN<x��am�sߘ �@N�5n�?߯u�	eйἛ�O�T�9tf(�) h�9��j{���d�駟�K�J�hl)Ê �Y)V�Ǵ�%������R�y�	o	6YR%R����s BUo���˪�~��.�����>{�X*�P�6'\��%�d�Ȼh��n]�����@-6l�Z/MQ��.@��K��m��u������V�9�������P'�r��99���GJ�%�& G��pk�Ү�c���:l�b����
ݖ�T�)�٩	Aw %E_��b�-#K,7�K�Sjg��>��k��4����*�~/���`\,�G<��N����_b"�{�X��Aͧ��oR�ߡ�43�;>������W�㵇�P�a���"���o�ݻ��s��fgWk:�C[p/��k�E����%���[�����pk��ls��8gm�.dmb��Cn*̱�Ѧ����w�z)j|��j���l\׮^K{Y��$�&y��;�i�U���kR�ϊQ�&���B��!��ի��!��1>�[��z���?cr�Fl8aUh�+���R�����k�D
���ul�^��@�X�FAI8
J��s��>��bs¦;�_OW����R^x��Ku˴��9�,���m�w(��SJ����YT��}��*�Ys��;}&U��w` v�p�R�!�v�����4Tmnl��pbL��Cٍ�ѺI
�EH��ʄ*���6͜:51�0iQ[���R��!9�i�f������j�%��w����@5Qh0��B�T?۱�kj�8"y0��'�l|V5Shh_~�����dTa���˪��*�N��:x���x)� ��/�H7� Z˓��Od!�=���\�$�e�5j�dG�z���}͉gK}��T�-�x>�0�ꫯ�!�xh�^pܠ/��J�Yj�6o[ll�w)��R��ʬ�tj��v�A�g��A��7�y���^7�Cl���;�Ox'l��X������ăE���b�B`�mb쟿x�~��C��W~����!�;��846a�_���5O� ��~�}��+4v:�R��VdLnq+?����8��%S�N�������l�m<��5�������i��Bi�U�#�3���"t0����SN�����Ζ+ ��gx6c|��w�>�(o!�R��]��R2a��A�(��}(<�3GM�{@��q�
@:�o���UJ����b(���&������{ᜯ��*]�rUڠN&5C��Θ	�ʨ�3�&4Q����ݷ�	f�k4�Pq���X��wK��Һ�C�(�k�_ntZW��R	1A��8���#�c���P(I|HI�D�*�Fh����|�^hN���w�eĄX`b��U�� m�)�sf�{���s�E��|�����nb��n,��2��IE�ӷu#~R�����_����6�բ�PV��Łv�,:�$@_�[l�h'�SD`��~�p����N�R6�����A��4�?�(����f�S+u��7�uZj%N�L�5�^�R���MQC��i�m;���-Mܛ&���d�J��#1�TL���3bk���^%{h����/D�@˔r�A��ϚiM���h�gp՟K����Έ�{� �K2-Z%2j�-�"A(���z]�/��P�GՐ �	\�����B��`Zu��ćb�e3���,�Bh ����#��� �$w�H�ZJ����Ii�ݘH@�����*��ܾ]��KҮ[�o���e}'3�I��C#H8>�%nҩ�.��-���9�#�y��I�}���0��"��+�l�[M4h��,4�	s���Ï?ԍ�7qV"��*~8���^D;��ע� ��`ΠO�Rmm l�؀����V�e��ք���G:��˿n��Ǆ�����n�7���薾�4��̻�ACQ��~~9��hj#�ϴ�S��I�*��L�����'�b�I<��˄Ƥ�{ﮘ�X4R~�$�tZ��ɉN���>g���X/C�b�(&>4��z��.�h��D//5k�7�y0'a��D�v���8���Bx�T����kMj¬�	�w،I2����u� ���w���" �e�z�m��+�?�͍@ &+�!H�R6;-4��۵Z���U �+��e���.�o��V��P�=��Y�5����ܮ�ĝj�3E��82�~!�G�;̿������`� �M�RsJ�YU��	��_<sE�P�u�M�1 h���֍�V��B5]x��8��V�l��Al�a8������N����&7������2�Nʮ�L=��1�O<e�l�n��4G���<��:k:&&����{	�A<߷�~+&<�`��1��0��&F���3h�4��C��d�BkQl��f#$G��f-[�e�!1a������a�B�� ���OC;^%DBŗ��`VZ��ﱄ%{:m2S64�tfI>���3���7p;���Z������X9T��"*v*|f���������|�����q�`)-�z*\�SB����9�����mVX��,��#�	�Z�)k&�
Tu`a�={*��6���~�{髯�V�{���wfC`�0�/4��JC�a#����[���Y�+'�kG���c\�l���[�G�~:���0G�7�.�6��0*ӝ~
�8�Fa;يE�I�&�Į���n����J�NYv�&��CXv��	�)�(��^���\h	�ijb I2px���LC���Th��Ы�u�P��u�`1|��g�A(9�
Ly'���5������l����0!̰�mp�$�:�����nH��s���U�ͣ%�|	�12%f^C��6�0���2�Dê}�_��_�Շ%��jGpH&�vz�[�{V��w��5�l�)�-&O�B� {��XJ���J���s��쩻w�v9��ٕ�����G|0``�/���>�����w��G���o$&�m���M��גz��魪�b����^�sBW��L4��W�ӶG��hU��|$��|N������g����S��.�o������)O(�m����z�b\�:#�A	��Ǭ'w����B���|?h������qw���J�f7�:Z�����3���U�4�Is��6�X����@�pюy(F�2���粏�5��H�x�:�5�g}����M^��&��3�f��.vH������"�]d��6��8�'K���K�I�-��06h�B������@mN�v���w�/�<f���`Fs\b<�
��0]ٿZ�-��I��y�+h��T�'���/�fe*6�;a|'�!7�����Z�}h�b	��cS��aZ1�d�(�
 "8���؝˽p=���k��s����-[�C��1?�̝}�o~g|��@m����uN�m������9�JUIi*���?ٻξm��Z�h�	^Z|�R0/��0o������G������vp\��h��T���"�V�5b����6��gfAC�f+���^�D�3	m�� Li
�am��@�a���)·�L6P�a�}�l�0���B�����G^�Y��H�i�Ԝ�9t����
iE�m���FK�AA��u,l2�ú�R�7�e�xg��6d酥՜b%jJ=�i��o8�[���Q7���|(��_|�e���?��>F	�x������	bLp_D0@�II��ʆo�#
�=�TX/p�}��w�p��U�<e�f3�{]x0?��@�%�W�HKqo	˫�DS�q��f�3���xS��� X�O���Nq��@�	��Cj�lX=�X�G�f�x�C��L�Ri&>��3ĺ��G}�p!3���yhG+�"�A���]�/��DF���M�)�[T0�����X��!%A@D����N�_L�b�"�	YDX�G�
!��/Ne��[f��.\C��oē�E �?��3#���o���.��
:���H�ڪj�*�,�o�:��x��i������߅�ͥ#mE�y�&���#�sF�؜ -޸��ԲП4�GR����	9�"4R&馶�C�`�AJ'"$!��}�^�p�0������R��/.�(t���Mep�?��,��U��y�x��{A��/�@U���r� ݼ�΅+�Ly`���8gO���w�w#�PC���4�Z�3l4���P.j�p,"��]=�w#_��$m�!h���7u
�La��r橷6�b-���c�}7��h�Q��n�N+v�F��v�)��3��V-s��7��떡5rڑ��d�0��Z̦�6����*�{�E����9*D %�!5Ar��m_�ZOJκ��D�9�BegxF�J�P��B�L;Rh�����+���K3M��"f�O���z�/���>���8���2��@��.2a���}�q�{FG�^� ���Jd�����tW�������ٔ�yД�	��eUF7�hV7J=�V��T�
h^um�q��?��� A<���B��zdRI�R��<�Q1�d�,Fx�9a�,0�7���_@�J�_nߺ�>��s^{ڭ����k׮�@E��C�!�y����hd
��(�&�g�R��2*F����Z$柰H�ł��"�&>6a��������'X#
 �1��ي�  �gB1�Ïyr�;��v��?�>��"��"��L�KM'W��f���~��)��V�COk����p���ܞ��뜭q	�V3G�i	�wL�D�%�~>��"2LF1���T��S[��=���.*,<h�8���DB�V0S�a���V�-&U8v�܂Z��&MuZ{��}Q�nf���9�dYv���*�H��-}T�M~��ר�I���P���+����L/}&/B���2�v,|��R�i��oA�4'��Y_L>%��(ϤO�p:6�lۊ12-��N��k؞�������@ӆ�!LY�YW�cX���N5�٥˦�&~�E)p��5�+�I��V`R�!;X3�:@��������L���[�|�Q�e�c�aRqImN(d��!��T�d�o<�2���A7��$&滑_՟��a��^|HLe��|ؑ��Ǥ�1��3Ϝ'-�(��I�L���g��9jՅL�&�f��?w,@�T�KjZ}d����Ex�^�cq�$"��W�h�a�v!��/3��V��-�kV�H-D�Cw�L�Qkh�E)ˡ�j�a�{Sc���+cjYSaC����6��J#�^��J~�Q.Rj%{�>��o�	�Y6�$�����P���/��3���	��s��lz�g)-��E���>�Ӯ���d0�����3��!����D����v~YL}�7��� ~����+�}'B_b�_�w)��eD)�I�4�@j]-v���}�x�� �p��t��U�"����#*\_짍���.
��L�F!X��i�i��ύ��^k�gߑ.ܬ�6#��~{�SIC�79ޚ�NɤE�D�)��_д��XwGL%�������鄠{[8��a���.w� |o�bH������4X#���
�eP���*LI\��ba�Z��)G*AѢo�O����C9�W�U�Ь���e�mf�]�<c:�����t�39����^N#Vy)����D��^A��o5�t�x/�A҇��K�ϒ���I�<�^�Z��B�lLsj�"(�F��f,��3% ��h;zn�1�����M:]%؜L���?��E ��~����<�{l��x5�X��L����/���pĵ�O�ޠ��}�N�/����ŝ���_X�=��y��O���A��.4�F7��N,c�J����`�-*a۵]W�#���o�Ҷ�q4�P9>��aMJ�A�xV�GA`B;`J�
͔�|eτ7�}`�ǂ�)���;qF�x�B�c8.�,�]'�{%��R@�l,B4��W�"ƹ�%W�C�D k�8�A�T*@教���I�+IMT�kɮ������!��u�~�/�q�1�E"�Ԣp,��~#��FR.%��Z�����SM����cO�	���B0|��vZA6#��Cv�m����m�Z8�>c�>�Wh�Z�s��`���P�0�U���S�\x6��_�5�y�Z6Qh���1����RH1�����%��Ν;�/pU���0��V�u5"�^j��z���i��/���3�s���Og�c�N��D��1��&e�*a�������h����¼�⠘����L����ґ�c�
Ќ#|�q>�y >ɔ���^�o�"��W��»:����K/�(T�Ґ��k�Xp~�|�R�\��R%��
�V�6��(>x���~4Ȩ�=�|��Q�j�,Q��%�g�p�j3��)he�G��X\����
:���e�ءO%u:>{_�M5��iR̴b�0'	6�����m��~z^;TTæ��~��\�h4�gCt�$&Yl����S��4�e%�=7�V��x.0�+���\X8�^���Ҩ�X��%uWRl�r_�����@�H��ۺ��m�-�/)A
�MA3��K
i��_~�p5@@3\ߡ/R�w@��G{=�Y�g�N�����<�*t�2>�)�CBF+�q�?�\"͚����(�y�����F���L�UT�������� af��ӄ�a6�gf�)0��1iR���h�/�-$������������ ?ĳ5���W��bq�AB��������Vq �x�=@@�M�`�e�0�+�
-�Wq��F	�m��x�����o:��	� t�6E�$hs+�(K�g1�-�"��ˆ�MЦ 5�M(��M���Ԇ]bL `���ƥ����R���:�^̌b��ԣ�/�@�	T����7�ފ�g��U� /�>L�	����Il�!W{l寵P�:��`�@��x�L+6�=�{:u�p�E5Ә�k����Q��fa/�1�bI�Ɏ�Gc.�z�*]}wU�%��-�Mq�щ���`��wpJ����1ԖO��/Wͧ���Q�X�=��w)�؁��d3�����zM$�+�9Gg��[�M�#g$��\�Q8.M�V/6&>Bb�!񄻻���ZQ@����M��܈(�y�l �%����˖,@���xBI �S��c�k�"��(8����(+I4�i��3��@#$�� -��o���ǒ_oV�J�0�L2�`��KR�!���	IS��ߋ��m�[]�ёnn"`j; nߺ-LK��4{I5^a�s��ȱi�fj`���+"�IƲ�G�(�$����3Z��z�j!6��	샿5�t�bUJ����Ԍ0����]K�_�L=T���,��B�r��p2

�K6��J7Ø�y�1\�vU|�I}�60�=&4%�֨��9�2Y�':��OS�$������
F��s�."���Qn2U��D�	6������i���/9�Z$P?T�7�"��ݛ8�Y�L�������\�}_0֥NV/ng&"�g��W����ԯ%����Q +оV̤'�L9;3�
�U3�M�#��>_����x�j�W��]���U[��x��eYL0�h��z#!ipP�R����jv�K&,4|�4���|���A4pFC�w�h���,�_���RJm�� S��YLjw��|�&MW&L+�27v,��E��P��&(-��A��ٷ��W�^�[7nҍ�p��]e�ߕq=x��8�`M ������*�d0�|67��xB��k6� �A��N�_-�"�%��0�̪c9ouB��r�bs�s~�M�'�P�9�wq�ell�A����k���Y��M�mtٜ�d��R��K�㦅3�=%��T3���,7�v�v.��D��)�NuQ@�B�3.5�i`�^��K��p����G%�5l��炠��/�t�����L���k���$%�n	�a��-^Z�dh5���xЪ��V�;`h:��Z����㫑%h�]�|���� �f�"��|!i���o!�^u��ņs$0�a7��k�8��*a����'7JGl`o�HM,8�0���K*��J�!D��;6Dh�S<,�*�:Y:+ݾ���9�FP���߅}
07Zh�p&�v�/s���|6�HV+f�$��BK�HYȧ
���gZ�!:{mM�&a��)B��#�)�iGn�ױ�5�})���f��������\X6�����\T���P����GpvqQض,��͋�Q
�[�d�̈5^��B�7{�s�E{*�+PRt�$���l4aK� ��څ���)�ͬX�Y�Ҵ���/ O�f�Ɗ z�´�&���'���zd�ȁ�_R�;�B���٣f��#����6jL� <�1�/s��fie��?H�Ms6tYP�1����h��2߼Ѫ��+:��ǦY�Moq.�8�T��A0��~�@=88�L7� '���g��ŘôVrh��	ݰ����G�>�'�Z\���+�� ���%!���/{X�B�*�u�Ю����
!��'����E�_�=A�~���gE����sgW��הAa���aS���ϸ��h��(CcY�l`G�r�u���OzC�s�q�g�4E<D��7u�h&o��Q� @:ݻ��29q�h�+�3�0����@'�΅XE�=~���aV:�������eq�INm��SY���;��<�/p�jUQC�?q�(&��Ѩ�wr��H�������e1Q�	G$�f�X\tR/�����K#5a�?=���U�hR+�[�\;�֊�9�qҨ	}�H��)��,p�LwU���O�1ycsd��+�ߠ�b�D{ȧ`[���2_�OYa"`�G ĩ� �o�j�ڃ }� 7n"��N���aݗ|�CT�,��s���+��|Ŧ�kT%�iO��#q����Q��j�W[������0���bp�(C�枾{����[��Ķ��o~�=�XC��R;�Ƕ�C +��~t��㵋��RD�Z�ѫ�N\���&3���Ke��ef��;�X=V����T�v�q=Z�/,�03���Z�J��	�Tr�x+ON�s �X�� IP`M3rZ��gE٬�K7.�,�>��g���ދ q�3[�Q��9�$�2�"�.�	Bءb�C�~g��<�0g_D�g6S���뉡��/�e�b����?Xj6�Ss� ��=�y����~�$Q��ZT��}���B����[��Q����H�K�\ZRQ���E	���3�qh��:%۬��e�M�W���^h��N������?���~I��ۑ�Nط��I���ݽ#�'�⾸wO��f��l�#nH���&}O%_��>��Y}���f6ؚ!I5Iv�)�p����?v���~_eFݱh�ĩy�q&U:i�����Sn��]�� ��ގأ9��o�	HU�"�Ò��`�_%�j?l^jm�C��m�mj��), �@��{�v%ڥih�4
=;���HNΥ�'���q5I�Ӊ�λ�s��������]%Q(lQL�x�	0�B��p4><�7f�pz�vZ)�|��4uϟb�à!cوy�o�ێ��p�i����{:Ϥ���jM���l�b�x	e��zn}m<��4A��ߦ
K�V������mr#F'��������ŵw��Y>�pA=�L"��h���%qd�w�j�RP6ɢ��bG�'�|n�����9%��6���n�O����{YC�Ȝ$�9��%��fLa�i�ݩ��9�����t�S !����p� FH��&���rK�l
BX��x	��*L�^8Z7M"� �g�<s��	���&5;}���u��P X~�9���6X����)'&��ɹ8���mLܭfo�ȁ�vP 3��� sW�1~t�h̩�c���վ*���e��ډ��8ęA�J�A&8�e���B��-$b:4�`�c�)9���Jؿ��-��fCs��}DhY��j�U\qD�lBs�	b�L{�J��|�`qs����w�HF3��-��W,x������t5j%����m�XHr�W���^?���f1�j=�i��䁲��7S���F���f�PjJ��t�����Եk]��v���L�ܞ�YJa�e�j�����T���3�u�{�M��'߳)�*�����'y2��b�p��쇕�^qG,��lV�e �=�װ,ӛ������<�&�)PY?$��}�V�XK���,�����Hy��dS(�f
�����K�n��i�А[z/����SbR�ʲ��h�E���H�ɛ��� �6ȨO�Ώ}!)o�[�w|����D�(F�T�L�G���&Ƹ�|ԓT��n%H�y�y&A��V|�	n����}��ŸZ*���
������Cԛ��E��ޙBe݄�X�_3�L�i�)�G�N��{���:v��%�������u���f��F�L��m�9�a��������x/�k�3������X��8b�N�[��ĭ���'�wd���|
fIl�unk7��A��6�:����iz�d������e�HKioE����v?�u[�t�:��Z��C���@��M�e� .S��߮i��G��:Y|��͆\�f����x�a��ͥh�;����ǳ�	�%��$ǐ���Q�1γm Mȑj-j�Qh�g��4)j��6;��a�'����Ip��������ۻ~��bM�YkYx���\YRs��yύSK��zD�<�9~�{Nӥ�Ԣv7�3��0ju�-�t��v A����M�����VY`i�U��侦�T0,4b�y4��6o
KZ1z�
�&���ݜMВ�"Z���mN�U�m�+��S:q���/}�3M&��|�r����^g@J�ݞ�2<���	K:S�`{G
�ɋ��;�������ɍ�]�G��ǹ������i�y��i�p����"�]�E�i�A�F���/JX��� ��*�K#R/��{�&cW4f��E|xs��V�[	�Af~��Za@
��36���y��So�SG��o/Lo9�����Ni:"�bN�a�c�6����Yl�>��Ij>��& M����-9k$�
v������km���|S|�9<9��`��b�Dੱ���P U�@�����4u ��s� ���VN\�y㯛�ik��(���K�N/%��?�M9�.�~��ߡ�>�ot�����ޫR��Q��{���hK��� m~f��-��J��YBp6�f@+u>�StP���fq\X2�F�yܛQf`�V��)��
B�Ǿ�A#�&��q8��8�R�=� ��`��x}����H }wM��z����SH�����Vp����G����2Tb���gO�5Î5�tTGˤ����c���8Ͱi��ҧ�t\,CCv���a��柷�i���M�(������O���kMs��D��M*���Qyg�fk�o�e��
�4i�n)!{���GIA����lRI��*-���k�z�:���Dܿ��h��Ў��֤i�blEh�Vdq,5Zz����%�Gl1�-�:��u�ǧ�)忘~D-��A4=\30�r��5�?�ny0������-'p$�m�˔�4��oN�a�L��Z�e�-b�x}{.ئA�]M��p�?m�s��n�����:w���]�<��%#v�n�f�/\����ڢ�\{�<}-$I^�!����i������ڙ����78ַ��Á�Y�,�Kٸ�t�U^H&Dyt�0td�"fE���	7���17Sj��1�z��߾�y�ֵ�c���F��;co����
����ݺ]�ػ�U�g�L�}�5[���C�E�%.Dy_�Q�	+�1�g	��ĸ�>�3�7����$���]�	���Ɖ��t�W]�Wo.��Y3�8�7	��,�=h=�ݓ�Mp�Er�'�#^gZ���(e��̭�<��׀�������m�@m���VG|�b�m�dn=�i��8�Iؤsn���;'Js@5K"���s�����ùM�H��~�3m�LEjp�DY��:ǧ���0q0�/�bB�q��Ʀ�1Gؑ�;�+p�0��"���@#
T���e��uc����&�\3B����u~��^4�z�z��l
k�����ЛY���֎Nk����5޽Yw����R/4ܒ	בe�sL�-���[ zj��!�������Y�W��C��$�f&j�����w�K���8�4L�����z�i�zQ������*'�L��a��hJ�`��n������>,�2X��_�8�V��g�qߧ�V01ݹcE�T�+\`0+c4�0Y�U(ʦ�SA 5U4�0("R���N��)R���wg���r�B�8?֏��?T7s�m1�Ȧ�B���%S�ܹbfX��ڂ{ʽ������r�Cq��4{�8Y�����9�	_ �o��B�O((��*�r���!�=��V�>��Ӷwq��a��S�O�a��{ns��-�c�{�'ZBܬK�*eΛ��M��v4�ʻ��qL���������>�x5[��L�ԝ֜�\�Qk�Mܩ�$z�����2����q.u}:��]c�/�&֏Ql�P2�w:�\3���	�'�L��eZ��f�M�Q��VNoui� I?�^N�:�Y��ƣ���M��?������z��֤�l��c���	̊���?{���ȍmA2��Lɴ�6�u��y�o���'s��9ݭ�7%�MCk;l @&�����e%3���E�8�9n��[:��5�����w����y�I��ԁ��n}G�_�2@�uٌ"N�����b'�^t���cqV� ��_�-d^:
�w=��d��G�b`Oo�T����P��$w���=*r�B�ĩ�)��B��\Xft����w���=cO��,/�*��?��}���)��j*I��8F�)�.ʶ.WޘRZ0��:g�~C�r�T�:J�.c���e���%	��/P�t(bț�yNc�������Nl�&:������Q~Չx�k�mT��z�""�p]S~g�6"�m!��Z�C��Y�c0w;Nl�0@UI�'�E]���޷b�W\.P�^_���zƶ���'��H��D���c��zc��[@�	В��ri
yv�2u��}��$>��3f�qڲH�Nl��W�`�hoi�q^����r��Uw�aٲ('��i�P��B!�H�e���k ��c����S�F��ω[�2�E�jz,�� �٪���*����f�՚��&U�Cq��͔��m8O� 2�Y3b�'�ύ�����r[���|^_�欚�y�:[�s@�\�p5����z�d#���,c,�n���h��;r +/ɑ��/����N�2���&�hJ�b����P��>�Nf�K�x��������Ь:�	�k�3$�>sOj����o�]rnL���X��YO�g#[�@��埵%��j�#�{���E�}Q�^�?��<���%�K�sM
�F�ѾX'����������駟Y6��|�}�5[�Ю�`��A�)��o_���)�$N���_Qc]��V��E��B1J�X�ӝ�o7Gu"}sA񕕿�T�c]B俤F��B{.����g lF,<��`V�0��:? \�Vi�ЉrU�R��.���ӧ��~�!���/�/	P�������<c�-lӭ��E%���Ъ:�E���-������������A����n�lr���^���=Ǩ�!�m/6�k7�CZ�'O>歉��f��M�i!��\��3s�ظf^�:q+�,GS4�ܽ��}�����a��g(�θR���yx�����Y�ٷ�����8��/ip 굔�+C��}��^��}`�V�T(�iذ��5�+֡��q��}L��V@�i�e%�7��a}�	`�Su؆�t� L�=�#|��7�Q���і(�g���3�Ruk�A�����i��� 1٫�fy�0�/���YW=V�f]���4z:�=�ݧT*�@̋�yx��%�'0U��;"�)n���so�ͺ�Q��2WG]K�{��¶ �Z��|�1�WQ�-^�	f'j��x���>4q�����4�`��3hb���ǳ���?���E>a���b{�'O>	O>���Š��H6�H���=��ڻ�׵�e�^�vs�a��JUD���4& �c;�3�1R�B�Á���slۗw�4�y����#&��߬WR.��7g��q*���׫H����_cekq��|X\�uC}�YC�H�Q��m�yK�{[��qB{ů��.,s��Zė���[.C��y��M������a	�C�! �M깴���z�;rL�`��W���:Z�xpbH<@m������̊pe��m�K�o=g���oq�RN�c�I�"�LY�V�����he�-�� o�T��y����-(�o{sК����� ��4ȑ u���������n�����a��Q��H�6�m��\�����u�%S��닂[�po���ǫ|e�ͤ��8��S��Q��.�Ey�h�!������B�^�s��&|A\���֣���zM�CFU׭qڪ[��v�㮄6���lDd�8�#q��P��~﮷��ߤ ���*M4¾�QS8�U��\�p �=~/�AŘ�ԌHN��2�-�m}'H�U��UDW�Y�aT��^�����U��n�GB�U�h(�0����FITB�' ���_�-�
���J�� �m!;%b���f7c,�V��K��>��5ZcXR�pԴN2�b�u8=;��QX��!�;� ����0<|��H̑K�>�q0�0���~nQ*��F�Q���
G�iW��ːN7���Q��I1̕�
�>H��4MwԤ��$�	$�6��O �&��ld[�D��,BCf�粋��ZS���)T6O���huLz�A�N3�C�c�G�Ċ4�6�f���&���xI�:y}��6���|���ܛ�m�X�O~[�s7vO@�8x����D���\K�zD���^v|O��^1w"�e�@m�������>_�ϰ�0��CY�TʡEdaϨ�tky��ryL�8��o�?���NQv�]нy�1�Q2���.V�54���/h.�䶾wt���UN����az��n����-sQPjjŕT*i�KdΛ���'�QJ_	*���+���wEXA�B�4�	�(&k�懗Kf�u�*�*G�+�� �� 5��,V��� ��L �<�h@�Z)I߂l�k�'��<	V� <�	��3�i��X��o�BI6Nj$�Cbf��D]�s�<G�´0ᏗGR(g��<؋��zx7,��� B�9����(�7�%��8��cX P�	ȱ��h���k�]:u;_0���ek��M�y�@j�Űb�9��<>e���gd�BcnL?��V�9,%�P�:� U6gS���q��+����+���!��դL6�!��脋�7�+ԡ��n����%]�9Kg�+�t���u�h/e�)��mla�D5�Hm����u�:d��`A����s�a�R�ֽ�)G{A�B*����d:m�J���m=�:�gOq���BT�U�R*��3�H���^��Jq%`�ŉ�gHw*.���6�ӿy�ִ�N�`Yb+h�eJv��6K'P�H����s��P���i����1�И<�e�9O����4�Me��uCAa`�����S��|�	�e��!�^f��dp8=���qJ�fU�ނ�Σ�H�Č&�h�I�π�����-E"�ԁy� 񘪍q��)n(y,��Ld��e�Q���&�&w :�LC:��2���(�G������KuDi
�I�?ZbxI�d�-O3�~}���C��z��&�&Κ�PKh�3[����s�\I����Ҽm���X��~�~�34���7d_zZ����˱rmW�)��L���̓�S:�)��Iv8�{�=h+sgeLz���4EY�R�NK�{���
-m�a�{��`�7Ib��]�Fe+��2���X���X�v4
���#�����a��E3�Ϻ@���XV֒�Q{'�:�uuy0!G�ZS�-�I�n4@iYg����rq
4��
i�%��P�TV-��,�v5�jN)�Ny�g�:����,,2Є�PݯN��NVe;kL&�����2�s���P����[&s�&`p�P��u��@ܧ�����3������A�Z]��yzr�N������x�����cѧ��e�y���������g�4!�$ q��=���L�m�_�z^�|��U��'��G������=�������� �\�l ����\\s?�be�yK�ٳ�ؾ����ً�<��z�*�I~�M��>]��G�=p�˗/�N��6�}wt|D����yx.�'�&��7E�	���f��P��K`J��U:�9���}���!'K_�b�2z��u9��ǹ��Y-#S���.����d���qU˚m�cd�gꉠz`���w�Ők�e/�{�@�4�A4�х�����3��7���o���dKvf�݃�j�� ��NJ�؛?w������O&��uL$]E��ցl?�/�N!=dR�I"���2k�=H��P2u�3�(���R��z��c� ���a�Y�@�,��
��5a"���\��PY��fz�.3�^�IG1��&��< ��% ��D��e�H?J��E�Fshl����P��,&:��9OP��	��Й�gy�Cܼ���'@-��\���/��?�~���*�{ƅ�����f�{�� �a�{`�G��h�y @?��s���o������D�F�?��#
����Y`d �P�������_��Wx��%-"h �|���!oǝ�_z��ze�nLO3���0|�6���;TV�������_)���X��P���ۯ|_��T6��x��b��\I/2�L&p�":W��t�:/��lx,�z6'���ws�S�����>��ʔ|U�T&�}�k	<�$b�z"�O�MݿX��*��v����k9 �U��T�R� ��	���A�Gz7Z��/�O3��#9�y�� �¹u�r%��4���t��H~���(CjU��k��m�RE� �?��GT+����ϟ=Oό�_hR��K�5�����O?�4|��gP ��d�_�o,&(O�d�S�/D����	��ӏ�Yf�p�"�xW�- �����_�X�J%�ڣ\�����"� �,�ϟ���>����d�����΢u�w�.L4�s���d���느^���?�`l ���q%��>f0����O>���Ԙ%�
��������#���s��ˌ�_#����(ba�h�*��+�����ȁ��WT�'�Ë\�?r�������ᗟ&VN�23,����o�E�7�ɚ�m���������Lv�(LR�2Ii�`{���X��� �֞i�y�̫d$<��}��h3̙(���A��P~/T�ǪaR��X9�O�* 
��窚��[R�V�OoP�B�$	A�B;�ty�?zp/������$f/�X��n�%Wlg�휼zV�ð̬".�h�}	��d*��Q�բ����3�^
zP���{�߫�o5�	
�!��8
=�	�7�������w�}�Y���b0A�nWK�_AO|F�	��}�E�?���n�(i�bq�"=m��`h�e������(�?~'�ƹ�E/�攐c��w����s;��x�����/%�d|���6�G�UddR��m��� �W��e:�5'�QP&������>����<�5�{W�%���[`���;��a����@�s��Ԟ/:X0y<� {�y���9����o�E$���ӧ� K��E��D?<��)1֔�M��6��0����9Rc���^L���KO�����	r9��S���ms�Kv������-=�UpC�P�^D����D�N-90�m�r�xu��oPKs��"�#��r �yB�5����pz�!}*��2$��1��>���1B�	�y��%ۊtO+�`1J����4�N��Z�-E�$����e�������B>�}-��A��#�x�>��?��A�{b1���1MնR}a�p��H�����}���ٟ>'VQw%��^W�vҷ���=���g�>�7��wXO�����69y/]֤r`}�fŢ�!���ܸԊ�����u�>3��E�*n4y2��t���YE��K�68��mS�����("6����n�|���PųB@��b��ږ5�2�g��?����u;�~�w_���`����:T�Gfu�N�i\�[�5�V~5@����x*�I���So� ��\
峛��I=Txw�p��b�����M��~��H܎��CM�!�]Y���o���CF}O58�;^�p�eRr�ץ�gN@��<���*�CĂXy��UXg6���l�V�db�3=1�<hO3;Zf� vx��A	`�N��QI�Ʌ���)�C�`u�	���w�*����U+�Z�5�%>� ������w�~Gb8�k�|ad%_��%��,�`� E��102 *�@��-* �^���G~���,��8��t]�=C�g� I4]��$0S���w'�QX���O���s�;��32�A��g�ŒM��-وcTXh Bx�(�#Ó��#aC̙h֋A�f*�����b��Kx��_��\� ԏ�r=�=<�,�ۇ���~�#�w�� i�;�~�{�)xweܐ0NN�߿w_�\�]ISuRHl�:�����*��NĮP#�H���Ѡ~��LU
��U�l|�L�5Tתz�GO�\>�'��ĭ��yZ虑I+{�d@8��QV�%���jM��4�s��͑��E�wu-
�o�q�ߗmЊ2��z�E����<���v�T�|�y!�|�� >y��C8�$CƢt�l8'd+z0��&d���PGT_vb���`#p�I�Q�)�-�����4��e��&��MDLcf2���F�?���M�L����q�e�����R[�� LD~\W���	������(��1�,�S��rE�Nݤh��]
C���
m��MF���1酿����y���t`q`��^�2�|��j ?  ��	��f����xb��1P��»��w�``��t�A��,	K �/WˠN�`�P@����C_r�,!m���_`w4�k�,$'��8y[����w��s��@Is�(A�+���d��ҁl谁�	c	Z��8��n�8h�T��Q�}�NEwځ&5~)0[���4�y$�]��0KN�f p�EB�͂e/�l�V��JMt������T�%+�s�<ȃ���GF�!�C�����Eƽ< 2��fѕ({ �ҩ1��8@�%�8�ݢt!�ډFF���F��g�"
��������瑷��X
ۯ���>e�/3��(ޣ4m�Ly�'�-z*���o���xQVhnb~	LpL�� �O��za� �6I��}'��;b��lIb���	-�+J�XdT��$��``�A[X��q U��+|����/�_~�e���O��}HV|��y���t��	��$����z�nq�:X�Y\�A�ܚ��$"��O@4���@Gz[�*����ft*,{-lXT�� ?�� �ot;��W�ﾥ��E���5��>~��H�Ņ�ƻb�Ӕ��e�B*#��Y��#�"�"R$�hH���R$*2bnJ�_������H�&���YI����*��t�;@e�l��I�J�e�ѐ�wX�H*���{|�E��=rM]����ZÂB,����PQ�QCŴ���Hs?b��E��0�h��FdP�`YFV��i�9YE� �y`�����H�b���D�ď�As�;2��"��*8�1Fdف6%3>cR�`q��B��D��b��_�����_@�8�z����T�NEQA�IaB�'YDV�ƀ�d�B�W s���3�h���믿�1�ַ�:�`��XT P d(����&-.X<�`ȁ*�qf�����_��ȿ>|@�$��~��G2����O�f�z&����(��e^��3��#̏ ���y�����f��^����q? �~�X@��UYQFq�WR�o12����t8��ի�t�G������S2�)�ճ�oP�@�/��m�"^ ib-FD�x @�����Sx��3$�u �&6�I�}Jcߒ�Ś�;�:Ό���BP�U��G��dzޖ	Z���?�~qa�>A'k��X��~���`(�Ev��~x���Q^�@��}>y��^��.9��r��j"C,�!�P(�8�x"�8��XjDF�2Ơ����iH���w���I��$]C�g�����X��yp塚W���K2r��>��R��6e4P��Z�,9+�dD�1{��R��1[��
v�V⨿��Ւ]�4���,���S�T��>��qDbj���x�c-u�&]�Z��������W�3=��T�����j�PQ'��}>�@�ş�D���}���߅!��؛��1��=�=K�IEE0I�3����%�V_Vb���x޿���q��*T���2�A<�H����;�
@�&��F}9�}���`:���G�O�����9`� v�45-�G��d��ܢӰ����ޕ� �@��:��>�`7�����D}�'�6��y��=O�5U�# ���Ə,jþ�<?������uGK-#�pS�*TQ��Q�O�;�y;p � &dW�рiZ,"�9�U/�{���&t���(it^8�Q�S�w?��a��,/^����B�^7��-w��b�����\9C�ΐ���Q�dV�?�u�D�(�Q����.8����GyUBƩ����~�b�m��:�N�,T��AtN�ٚ�9Ƀ�E��z=|�(��,>������ zV�q�z�!�Wpp�Pj"�#tlQT��7`t� �D�R��a����5D]���O' RH���'�Yd |FL����ڳ�uK��q/ 41�?O�[�3ƍ=��	�������z`P�;�1%速�9�xWf�P��9:d�/�:�(A��C&������$ �AW��CL<��?��?����2� M�H�-�[}��"1��?7���:F�Z�9�{�9#w-���\�`���iႤsĉh���[ڄ��kQ5��T&Kƴ|?��g�}�%��P�+ s�U��ǟ��K��(����^ 5QۓKj`���ʿ��c8��- ����"�i�A1���g�Zl� -X�i��"��|���Acn3Ʋ���ċ�B��>�PQ�	T�w�� �X&��E�x=��ȓ!3�\׳L~���瀨�G��'u,�yp�FD~29Ex�Y�BL(-��`/=Ϋxe��p2f�V���=(��V]�0��Fu��M��YXg�|��3���9
0����5�%�c`� �$X�3j(�����J����力]�T��%�F0����������s��|A�X�� �+�_�,yE,8SX@Y��t�`�؈��\r��a�%$� �<Z?$Ƌ���ً��u�����e������0�ί�rcZ--�V]_ V��7l@�D�
����0� �^�+ꖍ�c�I+�(Ɏ �Ѩ��V�f��+X���<��}�ДUm�&�j}�`�^�J �v���ɓ'�P�3���dĂ4 �q���b�J<1x؍����4�GN.��3�b7�Y�[
�_��ڮFWU�RZ�["ŨٙDX6����6_KQI`�B��֡2��T'*7�azO}NCs��1��������d���(�QV��H��	�Y�p���t��s���-���(Lh���^��h:f &�f�yp̆
1��41>�_g0���D���G����V�3����<�n@d%y�x���,�VL�����H���(jf0;���8���
5��Hb�1i9��1���ù�F�7�3
��a�J���0h���L:gU_H+MZ�<�9����Sz��(��*H$�ȣ�������-1bMF�F��:$B?�0��h��2֦"��GH����mX9���!�F��g��Ң��H)�,�F����Z^����I��?m�'��f��R��fѲD+�U.An������ʈt�>��"?T$5�Q5��_��������ŝ�U���1��0U�Łk`f��5�EKy��c�$����RY����xǅ 0�Ml,WQn���>c��ʋN�-y�t5;Γ�񇜾���,<?G��(]��X�`G}9�y�,�'�B�E2(-��Γ_��%"gp-�h��N�슒��TwU��_���i�F��M4M�K.�,��Ơ�Q9�tN)�ǚ&�J���(�2�X�R �E�	a�d�5� cU'���G�̆��[���	R��$Yuq41*��fX0�o%���e	�\2�I�R�W�O�R@��&��L����������D�X�L��ɔ/��R��m�@��ho�����>�XNn;�,����#D�8T��3و��|Syw5��v�����hL���uBe3�?�̾���פO����b���Om��ς$�1���X>������wNT���A3}Q@���1H��h�J~,����Bq�R��Ƞ�C�4:���r���H�u����(I<ƴ&��WV��+��Cz���,���S�7� �4�7"�Ujm�	��L1��
��r>Er'�˂|U�S�a^��CQ6�T�Re}:�����sb�Hp�J �D�������4�i��u�n<xPG�Rg�VlX�1�e�1�ġNYp�+��d`�!�?��y|ϡ�`�e��<dRJ}!����^�Fp!�(�,(k��u��p��'��E�����J@f
0F�=I��ekoU��b(��i�aZ@5�Fb)J���={�P?
j�䲖 Օ���;)���Ȯ\P������'�_�{�{�����^PV7?�mf�ߗ�/x<���x%ޟ�Vs�O3�ܠ������w�Q,��LN��ƍ�g����n��a:D������M��D� �h�9�4��sƲ��эǅ��Q��U�T/"�飼}f� �I�@�,��{,A�E���`�j}FII�SA۶�����R��>|�E��$7�\�C��fm�.�B�ۢ�1yCWR�&P������}_&��Tjm�0Q1��peO��]���
��xr?�����|99�ǆ7{��T�_���rLR�~���0��,� ,x@��M� ��Mـ�DE�u��E~�x���J�|Y�MEeʒ%�](�^/�m2hB,Д�=ܕ5�Jj?S]�����<�H�1n�n�HZR�^����$?��\��0$�J�(., p�A�ls�]
� w� 5@��@l�U �u�Aq�U���.k�X��j�	c�*n���e��t�`b
�݋�� ,�Q�s���*�"g��d�C�#"�`�Ԩ>���4�~G�]ӡ�T�pRxu�
|h,4J%Η'�*�ԇ���������WY�Mj�r+�.NI%�E4b?�5=�:r`���q�h�>�Ě(�G�qh�V�Z)�r���5���b���B��G����c��x����x�W)<ً^��Ǚ�|��禗��`��D&������A��C7&7�)cC�T�-_�K6�b��$�ą�v���A �թ�(G	�u�D
�_)��I�6��0�T(zRMy7:�����R��,(+X0ݤzN(i#=��ǓS�yo�w�l�$����W�YL���+���V���ʍ�Tp��XP�Ht����xhF�(��,?g%?d���8���Ye��R^���(X0�,Be�;pL�=tbTsđ�:^E�[[~��^$Iu��0��'�|�>��BiWz����@Vd�����W��q��ӅU�"��G��+7��hT$�]
hp�XS꼳<H��@]�8���4���+ʛ��D��u_뉳�����nD�"�z�FT��-���:�p$�TqEg����${QLam>w�3	G%��#bG��34�.dP@��r0O���Nп>�����X�Ŀ�2�AIca�Fq���L�Q����)��UaN�(��i�8ⴟ���QR��{��E���W<��NSu���['n�}���[�-���t��.4s��}R�����/���$��R��Ou#۟�	���RG)f]� �Oϖ|��&4�aL�����*jS�睧$���L�M2�36
������;U����ֽ�m��y�Kц M�(�z@���K*r�1�y��,��X���#�&I��4�_n4۔�F�ʉa�$�Q0�Qc� �ny�ْ��#����E>~���e�I���"G7ɺ�*��a ���gu��5��4Vz%3������Y����\�w�"$F	�����'��	C���	 �+C�(�
�S0¼��E �3�t��o�����G�e5�/�l����SJ=2�p�8L��S��)m#3V�0�՜�3١�㨝(Y�hRl6��HZGuvq,q��܏��E��Q70R�꟒�<�R�>�/�Qi���:�$�je�:T ����~��(}I�s��S�,��-��_~���&�����/�z"�h
��h%G�(�{Z���$Y�x;��l�#Xd�
Mz�>����X4p��.2�"@�y�SF_��P�g������:��hG��vzm�F�w�8�N�d�Ň�5/z�٦��|�~��4�8�|��e�Kɨ��e���S*�J7Pe]K�tZ�b�^'5�Wd��������>���0"?'�,�ؐ�^��X��>;)��"�F�v�ӃA#Wr�P�!c��A]�6
��Ⱥ.�U+o>�D�Jh)tjH��Te��D�v͝J�P��JnL��! �(��)2 	��*�	�ԐW�!ļK A�R�d��������Sm���4����Ň}<GۢE�m��X�*�0��,/$�L:P��EHQ;=�q�}�7X$(���I�B�%j	�"�lL��D�1�F�:�%a}b$d�H�X����pO�%B������N}Y�\�E�¼+�.8}�
�h���K@�:�E{s�|�G�(�`'����s;�"f~�fd��X�E�Q�G�K	���Q����'{?�.���u�H���Cs]�unk�R�Hz盁����bu̞+ N,����k��7�V�ݖ�S�)j���,��RfƧ��F�[g��$�ʋ�`y�8<>zB~��Xv�������73�;σ��ޗ"��7�D�VЋ���ف���Eu]b�`+�m����O9��(�P1�G��B���a��/�D��R�K�K�3�iF��P5IE�P}��"7!t$>�+�jL�Ȏ��T�3Bz9Up�MfwdHf�a��$g.J3�8���-���B�3�2�B�p���(j<��������� d!b9�7E�eвJ����ͬxc"��t|�xB`Խ�ث`(�[�@Y5V��/ʢ���C��.X��8�R.�~F�b�+�.eAձk~���l�҅��i�����>~HI���,�:��X��dҮT6�H��0
Cg>@���w���
��� +����j?Y����Ư,���!_����#�I������V>�������$Q	\�
�j u�`l!�����;(ڐQ�*O���v)ڏ��#���4$΀�|r���Ӏ���`b���q�����-K�3dB
�~����xvt̫$Y2�V�'u�^Ȩ�	C���i���%��~L���>e����ҧ�`B8-9z��o��	It�Q6Oc1鈶$yD�
H�pġ����~���9iL��bQ>C���'��E��oQŅ�,L�P_?sm_��~��%+����Wf����_�=��ӏ���&���i_�Ȫ��Y�F�̚���܄.yiM�(�Ӷ�⣸��Q��i�3�\�V��";S<���A���-�E�����x.�W��ҬO�%� "�l>ಏm?�MIm��8������a��셅�M#��2G� ��DJ�����`���*{��:�������C�K�=�yPT�7�:��j�/%�9}|đB�����щ�8��n5G�=���.*W �Řd��52'��l�nUo,�ڈ����4�
|=�R� ��ºA�X8<
���������S8]�)�	T�>��l&?:@��ê}��q8z�0����p���o�H�'0evA�āqi����jE1�eP�DĨ��5�������o�ὤ�>%u����0 ���)^�w}>�����W_RRҡ恴L�����>����!�o�����ݷ�&}�H���N��#2�I��l�ےR)JT��,���p&G�֍l���D&8>b0��aM	W�
 ���������Gg�_���������\�u,9B��Cc����&#�
���(�������A���&zM��Y 9���Y.���2_�zj���d����>���~����ܿ��>���ꑤM$ϋsk��qm�<A2�s�FzM�A�z ���T�?�����
���R<��$��"�o7���ϛ�iS���0Mm��U��z�@:�)m��Lj7�9/���SA�H6m���J'Z����R�T}���ʥ��O��3��]4��Ģ��MY�v"[�+w0 ��r_�B<����p��i>��SނDҟ��|�lQQD|�|5���ۃGI|��]#�p0K�VK _�T
c[:�R~(�; $~�ظ�a�Y#�c��ybS�)��$��,�5��\L,JG�(�\�O2�~�����O Qh��Ĳ�~��aaQ�� wv���d��/[c2����Y:ʒ$��u��f��c8���>���y �.�]��N��ɀ�\��O�D rUGp���8��%��2$@}�	�b�6�Ÿ ��%���Ph+j��"t�������]�<���>����{�d��?Gs�?�Q	���p]{���&�L� �s�4f��
-���=��p����69e�4<A(0l*���ȳ;�\$��B��;��<I����ѕ*$t�5?V{�`�b�|����
D�"3�J�^���>��..�+��}�
�uF���(D]��9�\���Z�?���AD=Z��q;Ĳ�B���V�̪��AD�Ɖ�1�$&���K����X���DY�(��&�) "b�a�03�jz-����"]q�!m���T�|�)��[�(�R��ǒ�6�Hj�$����XD��dF��g�_�=�`��W/i�#�tx�*�y4�R���B�)��f�gk{1�Q{�* 8�0���e���ʜ��X��e��,է��B��e)�>]�{�5�Z|������{7�)�����4���C���<�,�ȃ
w��(��I|��myV��)8#�;�oІ����``:$�������g������:�B��j���\���T�L�AvU�Qp������j�-���b���T���P��*p�����ù97�߅���]�J�L�0C$���r
��>,0k��W�)|�w][8��&���Q�2a���&�N��5+q����EĤX�P0�('bݧ�=F��/H|G|;t�p�Q�
K�<�����9�J���T ��8��(1�%b��}�p��d�G2�ӳ&8��[�������	����_���H!^�|pݲ���jit��u�E�W�c�����:ޙ||s�f���\T��	F�$����l�
V$���G���]���J sV�)��օ�r���n%�X�������ص�}�(��X���T�C�R����J�|�|��^�B��`��R��������*�q@����&�905]�����F��u{��[�=Ь���R�=ǯ�^�}��|L �E#]5��p�F���
+�$��/��p�6�px�O>&�vOE��81��9>��q����1&/�����>'1@����/oЍ�$������o�{�X�,c!�'����0b��uf�����CD��h�l�K�$돲̠��!���?��Yp��PC,��i�ح���d6��\����g��"|(����4G9��	j�hw��&��PPR�[����ԿV�y��,Us�
�������4����@�
pl36#u�����s�����!���9�9�b	�g:Á�N�h���Z����[��f=� �y�h�g*.T�ۣ����]��ۍT�6��)g��Ki=��b�M�F��3Q 5HP���  �u�x���L���爔�`���!�T�Ȟ��i8��ڌ
��(���i\�$R�(E?E��k
=��)[��QR�X�3�ń$�}���w������_�?��?����E���$ʮ��m;�\w��H�c�'/{ ��������(�0,:w��$-U�d`OD��fxD!�N=������h�3�;t�
�z� `�lQ�F�Eie�F�O"3	�e��^f�7M����E�Fc�9L�HRu�t(�8
2^e[�q��]� ��Ds�ڨ��w3�B痛8��ͩ+�'7u�p�i�:�{�(IV�L��4��D�@M����0���%?@����z�y@yk ���0!��������^rnx����"�}�*��y���!2C)�pvec��?G+��a?�$�Zδ�:Z���A[q��#=�qY�L���]4���
S"&E�,I�A�MI=tPN}wB�I�y�"���yXhw ٱ��Q��8��	q
��ZP�G��f])'_Ѿb�����Jˊ���IK���&]!&����>rޅ�L�(]C�T��$[HN3�������"����"t,҆�ܨ;����
��������'�e�����a��a���t��x�`yv
%�@-����,QEzU��w[A2&�.fR�喷
P����q�4�΍�����b��.�N.������jwh�Zk$�5��j,Q=�r��?���g�g�X�녊��/W T���]�M�8�rFF����� ���R����ğ����dː��_�O�#.�N:L��6[Pw��F�z�f�T%�o�6�-(���N��Y�&yO/
�3
S��3iT�M���E �Gf�2N���y!��d�O1������a
=WA�j4�ݔ�&�OW;yWהe�s����Ws�������
���j���lXltc�nh��frt_\Ry{ U�{'�l/��zKS:�R��(zid��� g7��I ����j$��%����D�$B�@Q+���'z� �v�'e\�(�7t2�	���@�nVPA��~�p�����g��NeK��=5o-R�N�sU�wAl�b6h0�}���b�:�M�p��fM�K[�(�S�*pv�w=��V=N��6ʅ�&b�Co�A祠*�X���6X�#N�wߗ�̀>�
�[�+=��alIK�2*'���<��)�3%:21�<�䕬2_5����'o� �a١+��\�g�9��:D��C!Q��8���� j�1	�ǽv*�ys>;n�0Π+�S%�ߡuT�N3(�I�Dw5�(�"w ����B�a$����)�冩/]
�)[y/�'�̀�X�4:����C�I�ȅ-�)w����b����lw��-��($O½!�#xV�G����9�A��D$�Pq9�������X���`�[��k����(8�+�#����c���Ƚ�&��(� R3�Ҿu[7��!k�.�%L7u�q"�] �~Kba_
��'����ˡ��̸_�~7��e����4y6�"� �毎7}����LY4w������ �/���z�|SYC�@U6���IBB4�Irh�L0�O�~��ȥ$_@Q��:0��C���J��P����qK�-=؄7�� 78�q�w"7(2�q�z�� P�M!�_�^��Sث�<(��gl�����7r��VӜ���O:d�e��ʾ�uH"/�eK��Ce]�>W��T*$u{�Uo,Lu#nt�W3�9�Q�5)l���)���׫Y��~U�X�'t �C�c����z�%�Yno���ԑ~��O��5����o�5NR�����c^uW}[P7D��c��;Vj�S0-5/m�n���}�j��R��m�QDΦ�bTv��*��d>26\�1���Ì-�	��"�D�aЭ/`5?'B.M��ſPҜ)�x�EXϠZCEI�z�����"��>c6�M�� [�˿��or�W��)E��3��4����u6���'���K��������S�V<>�a�sI&��V��JU�,/E蜳RM%7�W֦C��W/��B@������S�j=ϒ�S��s��T`���"�=��4M�@�+�G{5�H�U��@�Mw(��TE����z+������%�$wu[�
(�Em;�mj:�n�q����"��Յ�3�mצb�{����hN���z����*P���ԈQ<�T�cO��[�V5�*�+[��2�WX��6���ӳ���8�jl�d����:{{�B�~REAU�6 Z���8R��*������A�� ~`wQ����"�+����2�b�A��W_�����cTI�� %^>q䘶ud����dɧ���+��N{�(�:eA��d�ɬ�6h{9uPP�+�Jr��� nR�]J�bM�.["�:���ܩ�m����4d�s�.3��ɵ�EW����<#�����>��-��I�l�R������/=����\5�?ۉx�Yd�0�n��I�I�WzD�`+������b�2�ur�OKǗj�ʽu����( ���qJ���B������,�1�S�T�s�V�G��F�@���E%.�(
�?H�]F��������g�hP"��{�d����-�iK���Zr;Au�w���I6}f�Z�\���.��($v
��6	�����K
P��}C[�I=��m'��ල���������u9�v�8eX]��rk�yn�Z,ˮ#^���AљN���˷�&�v��v����u�_-R���(�«��]뙢��&����4�_��p񺟺���*>����^��$E�����`�R`_JX�&D�mP�"��� x-�wG�VT&���7b�oa���zYqU�m��8U)I%O/��˾�Vj�}2�5M����Kq�z�$M�y�+H�K�2Q�:H$5��h��[�Z�����Uo��+�k�)���Fm�@��G���CK���^X�%H0��T��1��� �f�����x-(�f�1��� �͟뵩�{���}Tg5U�*wMl�T��O�n���Q��� ꔃ)0y�>�[��]�N�K�����-������N٪z�b��1���y��P����^�g��H��_U��̯WǶ1�r��1
����o��'��s�ҵ2��#N�������y�	�_��~���^����1���L���ggＭ�_�d���p)�Jt��\�8`Q 0PI!Գ^�qt�	�q��>��gr7;���_j&�7��:���wQP�q�ȏw�.ft������H�ff/��3`����M板lz��&W_b�I���a��Ŷ�Ü���?�f���y���y�y����09�㝥+�2��N�/��N@��^&f��4�R#'J���T�|�R�[Q�������N뮫:��׻� ���V�ru�'�F;?5��?=�B*�dLTۥ�&m���~������g�TU=�b8��Ec(��j�ھ�Xxqu��r����������XO!%��4U����9^���c�A�iH��d�P���$�d7'ש)ی�5�APV7��T�+Ы 0��hD�N�Aag�]d��<�hT������$N�0����	��&rMEC���tǛ���@ʟ!��F����5��ޥ����zm�U���W��ߡ�a��WnP� j`5|I3N�7�2�Q�[��� ��r!U�LX�"�^���º�%!�c��jߢ��[4�R��U,��&o���z�#c�U����u���?}�'���CWY�����W�c���3��Y5�}�$��uI��g�oo�k#�������K��g�MS�t)�`���tu3�?;�[M�T}�R? t�ڤ,��j�C��.��}�GեvX 1�����jyZ=�g�Y�ŉ�*�kJ:JhKa�>�@^�A�Hu]l���m���U��F)�絈�3�k����p��s��Bx.�C���?�L1��xb!��.��8�ZQ��؃�<��U7�}cF����b/��T?�nR�k��ϩ1�^XCp����*� ږZ���z�34�Ԅ�5���إ�2B�{Q������}(�W1CY=nN��+�U*�ep����!�p�����Gh�IUF��Q�I���?[l
:���ň%!���4��Vn�
�*-����2g*>*V�Y�j��d%�{vӀ�dm5��{�vP� �X>2㖔}�p*c�]|�݂Η�N��h$�X�V-c�jðoK�W�j&zťK�nW;OK�ͫ��e"��bsY*B�z���\���ġ�|v����z���_��i`ks]��N�w7_�:>_� M�0�ϱ̦U]�u��m��u��(��U��\Ԓ�)�ɹ�<�ع�D����D&�Fa�a,Y�ld�e�e���[�i�^����N:����������*��?Y��0������A�:?g����R�Q�K;�P�"�܈�Yu�1t�f�ѐ.T������꒩p7)�����=�u�&��Yҫ����k8�^"2��UG����{������q��ƶ�����i�kGC�l���Ӫ������1T<c��ܞ&��e��x�YC�������$���n�4��>�By�&�ְk��i�f�qb��c��l�lY��3�R�&�g^����")��fR\�s�J��:����.���gR0��d� �@i��y��R#g�J�	b��7�m*U�(WB��<OZ�TU5�%�Si,�g���r�5徾.z��53���ô����V �H	5S�7A��բ�@��J&�R���+�jU������l�^����Ǣ����-s75��;�g�I�2�m�u��J`�E��F���Rg�a:Dh�k�VQ�� }4��z,N_@w�����dI��%�HP����rjS���D�'[�ͻ^���M|��������!U �?O%o�:[�J�R��u�طx��m�Zܚ���2�N��wi�ʉ^�������9��MYh�n�G�6��J`��zB%��0��sj���I��g��H�JHR������?�l�sկҎ�d�]JNc˄��ɽ�+ﻡ_�,@U��M=�T�{M;�{b�~J�Mc(ɢC5���6g�{w�F
o>��+������Oг��c��q�M��܌��`�e(6s �{�����0����B۶ȶ1ڗSUQ�V�!^�N�Z
#�)ex�`�����2�Ԁ�'yT��ʾr��<$�1Qv��5ZE6!07�Ռr%V��
R1������
�{m`��T@՟�I}륭�[��������K�~]Q��iJ�q���s/��~�ֻ�*����t��.��������?���0��,�y����� ���f�n� ��;��l�k���׺����F��
�m��U�u��j�d���-t����.�U��Q�{@$I�Ѯ��BhZ�(4\�k}1�_��]%0e���a�2{b]�&���<���@5^<@��wh��t���x �\��nז�-}7	X��%)�YCQ��T����һ7�H���Uf|���JNe������X��r��!V.P�Ê� q���@[� L��fկ�S����Ӷ﷨R�����x@��\ݤ,�3�c~z&�G��/Xۯm2�^�S�NΊ���<��.��{G�q�S������S1�N�~�m�:t�Jj�-�gG}���/s��;���W�h��)*��mL�0��%e�s�j�8��-��������,�S�C�("��ɕ���N͠6Pl��C�3������f8�TS�c���7Ӆ�sϦ���攋����k��|,�mt�,Ց��Ew�\�b�mc�,�H������4��m��w���(�����CR*�kRI���\��;.}K_�U��	"�r+W���Kd��*��t41/�����UXmx[��sU�eR�E�F\�)kU�5@�_��4�UQ7��.��n�������X��WQ��y����]O�7v�Y�"E�93��ۇAk�:�����zJ\� T���6h�]���[]�y]�F��R�F���������m7Q�`96V W�F�MgZ=���,���1v�c�rd�b�}�4�1��K�����K���X	U*>bv��)�_�|ޘWl�F�6�B�n�m���C�W�V�vk�N����=�U�?.�t�g��:��v���7h9�[�����jV_߰e�}p���2���?|�Hҙ���ae���ۦ�N�E���'�'�__[8���}
�J�u
�|���L�M�ɛC�Z�	P�GT�B�WG�����{�ݢެ_/P���'�s2�5Ҟ�=�ju/�i�����\G�f���d���h?k��,���8s��^O�,�kU�R$�H0����|au���͕2@�����^���ٵ:^|s�t�|�Ǹ�dWTUȸg�P5�ް8�z̗]�B�1�Y�5��4��n8��T��.���FSF��d�$ �s����{�Gw�֬����Ϟ �G+��w���ύN�X�|n��V$��8Z�"E,����<�K���R:��cRݫ�*��tNyKV�5��"��{,Jo7��5u0�؞o��ȼAf�f�TM����X�S6���B��8��E���&[�Z�߽����+	3�2�鸞T�{|�cB�U{�-�mc��8;L70ٟs���͏���
�+�l���)�����2W|>�ν�?��y� �3� L7���7`���<K� i\�[tk]������� jG!�V%n��+�1��z�	g�g���<@Aš׈��Cnit�G���T���)j �MY�[��.�;�Eɉ5�w�"�i�궝�t ���ݶ�����ˬ�	�'�e���q\���mEo��ں�(犱��s/�_ד|W{�q�e�Ʈj����]ؿL]zZvX�M�Ϙ��ֶ�w����&�x���*����2��]��rv���Ç��G�	[��,�o�q�lƌ'љBp��\/�M�5��.��*��]�]�.�X���A�t?ϫƫׯëW�MT�K��<�M1�Ta���1�%s*�̌�mb�-�e�i�k(+��Fub�<�O,���V��:vX����I.(Q��0�z:QO����:oCYI�Ju,t؟�6��vxQ��m_ұ9��� !���a�@l�V���ܹϸZL��D�(��|fkzO�Nq�HwX�qQcr�&7���R>��p����L?|�0FU+0�\�q��W���1�+�1��k���u[��[��qa�Gg�����Śi����8�2�}*�}[�_�� �Et��;��-u�*"�4�T<�-*��)�𮃵N�0X���u2�[��=]PT��_S6����\�� 8�7A!�eBy�ej�M��.�}(=�k�+����ӴF5�U\=����Gt'ϥ�x���+��5��|㪢�{kq�`�[���;�s�4�W���^w'�U�䤫�1@��`�V��,O�8�	�Ș��֟PO�<ۡ7��N}���+p����nxZ��R���/�!Ȁ*�����P�3��GrM��1X�_�YZ�b���i�Z-��`oY��ܾ{<`»�-�|x6�:{мھ�N�?�d�V]\W������Ť�Z�VL�߱�W�V=�'�j�����Lq��oϹ�r=���Cڕ����}� 0笌n ՘$�SMT+b[�X�M��j���v�ݘ�g}n)Pw�R,)��\n�T��!�rM
�U��͞��f����������|�6W��nFւp�֨���D��P�z'�ϡx+�ya���k?5�^�Њ�- �D��:�:��ĵ�Gkox�([�Uu�������_([ ׄҡ�K+W�ؐ�Ы�a�F^FJj^R�9�$b[;w���gd��U�a�n�7�8�� p���ϊ�P����ir�]�"���+��Q�:�y�H�m��)�E_�Y�� �9������j���{hK��x��V�"�x��By��o)n�{�����P��s�D�W�-�'�{f�+�	��x����k�Sʿ� 9	u}��06�c��&���^ R��d`rƞP�.n�ru�Lk�Ɩ���'�C[�JVB{��H� ������0Pݢs1#��L*�*��}&��N�Q&e�MK�����[*6��b��[�_Ltj��fC9����uW_��s�$�g�3���\����Jv��)���QyX5���ݣ4�U�P��n��r�r����@o���I�܁j���"N��ګ�_�v����E��mפ Ã����|>D�6?�Ut��̒Z����P��&��r���p7qJ74+������*`��S��R2ޒ�-:T�r���ɑCQ��M���������Wr@Z�ğ�>�v
�����y��֗\.P/�cjȇ^�j��֨��DA�Jd�Z�T������$����ؤ�A����щ�vw��5hb��To���Q-T�L����&�-�=w.��Y�h$
��:�- ����2�(����C8���{�f8��[�v(k�r,iN��������$� �;��WT����&�a��Ƽ�7q8��4l�ϸ~t����~���a2	ZQ���m�7�}ω�w~_|cs�>�vP�1�CY�z��ae�S��I�@����Ŷ�.�s������� �}k���T����b������>xW�2��lR��$i?i�++����`���#�z�GdE��!v�X����J˒q�X��j�,P�
o=���;늘J���[!C��e�~,/�Q�����\���oN�n�GLv��QbT1�����e�W��ڭ:���V�+%�^�QNq�[�hĵ3�-� ��k�{T�S@�-�
������qwU�}�5X���ƅ���P�v��+��[KahU<�^<ӥ��bT��0iͪ.�0YU5��!H��Վ��b�'���-��[��_�U���e��{�J���qQ��XH�c���+�մ�:|1' ���r��TQ��y3i�	�"՜���7���2������e=)Np�]��tѩ���z�%�K�C�WD�ڥ��y,���\O�&'�n�N1`t��X�3T*����Pg�D�9�u+l-bLU���-w�a@4�Gb��[O��"ǵi�M��(UTھU�-�7���������g�.���ݦ�1уF����5��N1k!���Zx��_B�~D6�}h�=ѹ��HS(���	��qw�9�ڞk�%^%Cu�r��0э�DJVʋ���;�"���
nn�4Z`���
�Mʪ�Q|�^����bl�oE���CS��M��|Ҭ�᥀��Z�Tk[��Z��E��� 9�]�]��Y*��}O��P7D��?�~�zВ�f�v(��|ة�a������8W@�t�2ed'Lu����j=��K�ޠ\����R���25(��T�2��&��C-�FÔ*�էBzb�o����mk��I�2�I��#d_����ϊ�V���}�53H��/<pq�{������^���+�`/��nQ�h����(`��j�Bɡj�|~�r��v����k{q��e���]��8t�h�׷+<��g�W_'��=鯣vs��m��5�m�~]M����-(H�|�����]�+w�)7
�*�V��� ],�L���8���x+�+(�{�m���U�������}w�_n��v��f����@񚦡Z��]��ޕP��n[�������P\mM��x7�w��ͬ<�^�z�1��ݘ��������ٖ�7x�m]M�ʥ��b��>ʼ��E��[�w�10�����6���Q����(W��x�͋��c�7QD�p7�.���"f�&8������נ#Hs���,ݕ^�"��r�"�������2����z'ʵ�@� ��j�[WnN俍�$�I�_A�p�D�;��]�+w�)7Tl�KC��]�+w宼�� ��J�K�Q�p��/1JXj��R��{ڳ�jxj�,�t�~f~��dr��'^��y
J���ͧ��1k�*O��$pns����#,�09c�zd�����w[�����+�Ҿ�wir:�6�2�&�4[nWyS�߬��&�I�:�����7��/1��Ų�+D���4e�lT�7�68��+�q0
 ؖ�5*ڦ�!@�s�O�u�.|^�Ua�CR�83�������ҹ�;�+�������~�ٙ��n�T�N�:M�A3��)����k��I�'I�^��(R���k� �%e;$~�&R�}�m�ٌ���L��M�+B�[)��&�����:7�Q��)ny��5|�\��k��N7L�1��J$U�sћ�Ɩ%���gܖyr�:�9E�Q.íb_�;]��[T�?Wt#ȫ.=:I�޿R�w1�U����=�nv�@mD��.� 0�ģ����=-��swD��0�d�Nt]�pc}v�]_��������h�E�e(ٞl�͐�Yg��)��u}�m�j���c��>sǝ�.����X�`��޿���@��ǀWTV�� Ce��&��oy��e�4��)�*��I���ӡ]���+�zJC�+��ݏo3Y}� ���	魘o� S˧fv��|w�v�x#��	�`8W`�M������:�!I��[�e�2Ӊ����Y3����ci�Y��3��Ԥ��:H���R;� �쀶�;���x<l��E���-`�R��z��F�
��W@	��U��C�v�i������pn�׾�۾��ޅ����~�Y�*��]��]�ߕw��B?���{r~�Q6�t�Xu���o ��]_o��0��{����+�Z��̻�Eu���� L�w��o����`�r+ u"v�A���1��R�������{��u�9����Tu����<������jEKk��1� f�;����'�=�u���8�?�����Qj��T�TU�G�u2��� �=;+n#f�u�׳�1��:�7)�A7�~pMni�܅�%61�%}�1$��:�@$O�~�}Ռ��[?u�R�T��Ck�D&���H-�-1Z�YΟ�{��'N�~]���%V߫��7)ǠA>%A
����pq��F��Ň��H�B�Z�dǉ��43L&�՘Uu~�èC䙤�a�g���x5U��lذ�� ��乽�t۳��y��2��7߭��_�i���Y��n9�in��$���L��\x�do�<y���75'x�摛o�)��涕@��ܢ"c(�������]9�D�);�%���8�(�X�P�>�N��"�s+]����O{�ls��ˀ�uu�m��g���s��2� _��v;��)9�.��ͩ�?w�ui�ׅ�%��
)h��k-7�5��l�`�����%*�Tn�2�]�� ��Md��vn+pW��;^T��TM�قjU��S�W��[v�L�`�r�ϋ�ܱ~�]<մ�Pv��������������c���(�S�O���,'�$R�>B*ʋ(��ZG�_q��i����(�NW��+-�k>Zi��]�ۇ�7�6���D�\�~�j}/�S�wc�@�/'9=lt��ѣh�j���ݜ��[��I���M5kg�L׳�Pn�j�T?-j�JUդ8(.���˟�Q�g[�������{�=e�2�S��>UZ��?�T&vI�7QnP�n's���3�����'S���K-H��tA��_�3{G�xѽ�t��{[�/�j�X��^��z��� �0�9��Jt־-nȍ(б���b�����jە���MG?���Bxʜך�
���.��V���ηuYx�c	N��P|#�j���8����9�ҭݽ��TW�z�ө��3�X ���V�8��� x�+��]ٯ��D���PQ�hcaf��T��ސV�Oow�{�^.Ƿs�C��P�����A��u�R�k:+�+�X�4���u�M-�u���k�����*Ó��g�.&4���*�Ҟ �v�u����~�X��]T��$25�_��n�y"�Ξn[o�&�+�w(������MJ��,�h� �3>i���E�s�gkr�+ԏܘc�/CB�,�����S�z���B3U�T>���4J������Ӽ>U��.;��RA�;�%���\�-�nۼ�Vf�8�Ք�XnϠ��'�;;jT�7褪Mc�X���F�}��#鰙�nc���tK�Tm5��b�mϝ2ʭ�;�$7�2��3G)ʜ�#gk+t��ԯg�*��-��og�Ҏ����{��ԅ��P������z�����T�)�߮R��= Z��Ǌ��K;*z�Ns����m��E����b���>ZR{ǽ��%Ӽ��jS��F�]�+��h8xl�li�]�ݛ�7f�ߗ��^&���ܕw�ش�8O�!$X�٣�y�ʍ2T�-�z�:����]��2SОR��~n6n�Ӳ����=���F_p];�\E��H)V�֢B��v-+oѹ�:SY���y~y[��]��e�H�g�ںe�ؘ �jڗ?����鷱�\�T��R�#�k�� J+�h9�^2��z���}��b cx�x�-���&��������kc��wP�r	���:z���>��+�p���z��L_��r�<2��F�"��*�񵽊���w��-������1����s���N���49��,7�i�ȯ�c�mn�rWޡ��fu�>f�9�[�wuF�z?�x�%�ܕ�r酁0�l���E�m ���P˞Q��\(e���v5�]}��7�Q��A;�%��[����?rg��'�)Hmt�>Kȴ���S�(���|�þc��w]��W�X�!@-�GK�-��=P,�h�T�/��֯�3�5' �c9��6%?����{�������ɌRɫ��M�;��C1ٟ���;�iݺ�!�^A5���x�0w���=�?;nѳ{�s�� �;�t,�˯+�]��f���'�䯩Q�J6��&m���t��,��Ǵ�9����]hh�\��I���<�C�����8���d��~c~���
��c�1p�n�i����W�E��m�U���TjD$I�Sѵ�j1�M��p9�����߬��9��S�	]���3z}[&ʎ�U�֒ɴ	6Y,)L���<��#,�m�`��&Cl��&&&�X	�L�,2�W�v�&�$��ԩ���E0��ﴽ��iU���ru�Q�?;4���~��4qB���<�K���v�v.uύ��Y�5A���DG�����Q}b-%#U(=u��L`����{��V���U�M�~��Vv������b.�3 �c\�q�`�)m��jB�PrL�N�5���YX��	K���TB'Nr�bS�󧓱:/�pQ�j���X����A���?��͢[j�|���1R������b�֙��b9o��&����X-*ժF~s�?�=�_���=ԭW�	��wC��ۿh
�R��p�W{&�
�&�������AT ���>��+����vb�����=������}7�~Uiب��HG�゛�ᛞ�V�Fcl����IiD����N5�J�lb�sw-����(�>�
Xv��`��2����ɓB����^��D�}��tM���wy���XU�+*�T~��/�1�|�hUw�lB����}^S������p,��xWq\؍���W�8��CV�\'��ݜ_�(e��Q���+��{\�����{��u�wPM���	5��!U���ͨ�����f)���M�;�����δ����WWby�"ѩX�vi3�kI��5(�t����:ѳ[�ՖB�k���ם-k�lpAQ]o[�j!��/��yw�~�}'O�,����j
?�&Ų�dѓ;pRj��V�S�cAN����x�@}��4��54�Tvg�7��>7ޓm:�U�	��f�VZ5P%f��u��3���;��MF'�� �J�k���c|Y�gXR��_��2��N�n)��8�w.��WW�9CKꔼ��y��$d@:�o��m�a�u��Ȗ�i��S�o�T��|��2p��J!K��W����;�j��R��{Ů	�)��b�Ϟ;�4F̡�q:�+W/e|]�#MQ4T�b�0t�f�
4�Ӵ���0<��̴�2K���g��Rέ�	��

Oi^[G,N�[�Q"�Y/�=�nִu��;�{��|���"�du���Un1�B������J]m��Y�	[@��;�V<9�RGo��A�����G434���b]�(���S��2��"�'Rs�K=9[z�O9��F�M��$UgGj��M�s�O�>wǠ���TD~y�y�i�Fb4bj��ɫ���j'��c��5�*�ރcs�ͩ8Ħ?[����H̶�[eH�E��+�4������X�ߜm��/ħR-n���Ks�
4�g�|t�<�Zo8��Dă}˖PR9�����_
f�jݦ�]���u��"��o��M���~�|N����I��9�W�1�
�z!�d�T~Ӿ�w���'7vk�]�s>2Fӕ��d���������e�i@E�SvZ��#?m��9��%�z�5�I����^.��v�D�nA��2��)�Z�4�2|��O�U��xl���==�������|�)K��s�wܷ\4N:}�݁�{˹�[�ں&�][�"P3a[T��+C�qK�8:Q_�Z�U��T%C�T�{>��܆������i���޷�����ԎT82S���ܤM�,�v�)�c}ʶ�J63�b����DA2� o��kw�{�Wi�W��;��Q_��.�����p��u���&��o:��$c�`˶�߅�:��H��R�_�g{M�P5�7X�WCy�h����++���������ڗ�B�>�Ԛҫ�9)Ճ4��
;)a�[K�9-�����s�X����X���P������y���>"�~J�b���Y�S����D�>c��?�'�cX��-�ڂ�k:��qP�J;�o����;�I�_ԩ���dMNMAYaꂣ����m�+�H&zNy�S)����,�#(l��g�w��Sׁ����jkj0�6N'-R^�8�ά���鵠Xn\f��X;t�kI��`�w�	�{�*�Z|���J��#��?��^���S�0P�UX�g8E�6�]�@W[��umݻh;��R�5��4w>e��*�LMS_Ljc"���$0����}�b��)��P�s����I�X�aZ���@U�L�g��A����9F=>H��''H�?qp�9��,]s�.�k��Ğ���cE�0��k 6�xu��4@�չeڇ��,5U��O[�V�,��S>��ɽ},MF�Q�a�o\�zO��~�g��AW�+�f������[����������7/[�c�ڞC�����eM�)6�b�b��k�N�µ��W��+1
P$�h*�^O��
tS��:V8�~�+9]�������x�>�2C�yÍժ�w�r��n�g�i
ݦ�caپ�^a���+Gpz�V���u�xw���P���j�z�ĸE,��Ȏ��gZ��VSd)Z[XWm�N�
�E'�c��?{o��ȍ,�U$���}�3������9�x���RK"Y����H�(���{��e�%q-�Dfdd�-YaK�.C����?Y	������7��A��=rG�ۭO���dgT�ٻ�]���>�6�ǂ�����^P��',�����"uX����"���mϿ��B>��n.����G���(o~F����G�w��Em���8m�q�A�'ݚ���'>��6��uD��(��.�ޣ�����Qny�Π6�D��x����v7B��Φ��3�o{��Wo6�N������nyݟy�0ѡWz�}7�U�筧(�ǧ{�mP���.���Q���������蟂�E����o�L��/z	~h �?�f�����8�4-��L��YC~�j̉�)�o���O��#��#������j"�{[4|��������'Nؽ�LSj�tYB�>k`�ˏj�WF�fV�{U.¸����p����Y��6cz�|���g�HޞҡF��_|�������O��۠�rf�o�HR�u�{zx�b�R����R�����|���ڧ��I���U�����xysC�|�aTrG��=��֤T�J_zz�{�)i��ԃ#8��;oN���ۼ�����3��&ͷ>��W�}����:/s�A�n1��X�RnY��w,�]�)���/º�x���nE6T����#��Sm!��g��cڛ����~�mP��7����l��+=�o���ɞ6��sn?���5�Վ8۟Z9xM����ݎ۽ѻC��n4��w<��mQS������E�����z/�b䛶#�>;d�F"�|m�_v��-��mJO�Y��C]�Ӽ�o���4����R�x��V0������������];�<�c�4�K;賨�������
;�?��,���7���<��-�A<-T'n=�ÓhI�|����]砋�?��9�4��fq�F�'�9i��*��d�tP�}X��E)�������O��V����v7lr�%��w��Z֣��zCؽ�T\�~�i��~�O��������j���y�X�z\�����irU��z������OA�ǳ�zj��V�u��u� ����{꼉�����}s�� �r��'���w���h��\.��uI�w=|zi�g>�*=�缜��al�����}����~_�V�{��:ͦs��q���uH��V<����⒩N><c�·��;�<榁!è������{aTm�����R�浪X�#/[��gr�/��C<G'���"ǿʤ�5S�ˡ��ǁA�+fM��E��vœz�GL�C|�nA跘2��6�+����XpO}�4Ǯ��n�b2���s�U5�X$0���Jj>6O;;�uN�O��-b�Ms�?EdlgJ�Jᾡ�9M��r���L��0�Y�ڗ�Н�ͽ&�&u��G7$>,IC�8���`b�ٳ\�ˆw���U�[*)���m�oit�fa」��C��Q�s �����F�a�|�<�uH�sf�� >>�����\��3I	�3��3�C�"��5�w�F��6ϧ�͵B'�<��A�F��NL'Σy��N����I�?">7�i�y[/T��1�ں�������d�y�����u��)\�������E;�>�z�Ooͼ��`�IZ�MS��Q\�z�գ�T�s�x?.�����vK���2���f���uZ���8?O���|ͦ�wtt��M,��5O�z��r��f7�����9�Z�@��^A��۝�_8���ɭ�{Sg%�|��%�t�f���cs5$|�����~�Y�P�}�Ӟc���Ҷ�vuw5b����������T�F�_�b�7�}S�{�����v۴��Y�+4sx�v[��n���j4��������5Q��㺬ߓ󯾆�uM���&����e�ut�(�O3�)��� 5cO,oΒ�����P�pF퐷>���zsaLo�b��^��M;��X��'3,�"�0��q�]_]�@�ie����>���������'O�e}��{������1C?�
?�3��jpͨ��2*��txΝq�Kݮ�����IN����VG[X�]�c���wzp��F�B=��̺��n�z�yF^;�6«:n��R���k������#n�8��\�QޯE 3_�������KIO�H����|8������~Z�\�e%8(�g�^��Z�k�ƣ�T��~ S�~��g�����L��Π��g�徻ͬ��=��,꭯�(�~��pi�0�{�-�{�&��F��u�8q���3�����e���]]^՟��ɬ�06GIڐ�'�����]ox�g�}��Q}������圦�jl��6GVx�a��/F,nX�k��/�Rx��*�:4w]��~�r׽����Ӝ�G�i�C��#:�M���S������Uz��E���7�u������_|�1���X7TFm��3}_��gϞ���/�#l�0��f����߻?=�����7�C��)��}S�g3p�g�������J��8�{�1��^�����"�����	���.�f�a�]^í�-�m����y��Y��m��c������=����lI�.�T8s^����^�{���c��)�%z�o�׼��?<o�����"�����NO����sA��Ϟv�ԓ�z��I�yT�o�������F�ޫwV���fޛ{��`[�#��Q�q��;�C���?�rS�}�us&�����?��ܢH�y��MNn�`�x�����@a�^�9���+/s���6u�=>>��uʿ9��|�ͰN�{�8��^�_0�!�4z2��W�?��G�=�h�����tT7�f\��q�w#�;��T��G�z���J��P�j��U��dR�h�k�bP07�����9U��rݮ�M���������;c�L�bW��7o�1'_P���g��A��87<�NLjS��FϡNp�3qк��߻O�X��ׯiD��.L�c���rr:�B�����>��C@Ux*�R��A�W?�{�7
��Lt��2��a	�~�Ds3n������rq��\���A͋��m�(c��^?a<Y�5<���_��������F�~dn������<¦Vmf��DC�yq}}E,u���ؼ�����3����3z���jd>|H��>�s	�.���yT�+�6!���z�!�%)
tp*�λ���9�&{���_8?p�_��r��,����G�}2)V�]W�t ��g	��!τ���.�e�L4��G�E�E��ull['=qRܷ��㘼��gi8�3ī��v5��-T<�W��O?������D-���I���<#,f�	���=�^�g��^���y�4�Qz�4�y���xc
�A��pl�E-nn� �B�����;��vުr�-@�-r��]�?a�h@�����3Du���%\c�Z=S��H�K��c�+cl��}��"��:'\�g0��Z9fH��)�����A���ߧ������J'5�'��hk6�}����AR���֡"^⻢y�|��y�B�{ϧg�,?��������F�,;��f0F�m0	��4����G��b�_M���)�oFf℆G�&���ʰV�� "���z���3z	�W|�{]�|z�Ր���ӳ��,� �1>cf���Гe�8{��!�zhH쯾�����[�=����k[������z���,w]��iH���7�pۤ{# x�KUY/�L}���[?8�ǵ�GDR��v��1Q/0b�G�\DfH\SA+�S�x-j�����)Dcs��|���å{�{�;�����0C�٣��� �U�΍b�(+�X�w��Kҕ�`���m�夛�x>��|��$����N,.�^W��}���ȋ�E�`A!r�&,i/[[D�=a���!6:�WQ��KOLM�W�����G�^�����s�=�~�����o���w�v�x�~~^1��k�f���X<x?f�����z�8_���a�Ӟ�(�J�ȡ�rn^[����k�m�܎��xSb�,���r�U�ł�)�ю�a����y�������7�\}���Wn��%n;�'k��Ɂ�V�;��*
�&����������`�T�@ct����~�HXT��'�I՛���#��?������~cb�˯�L�~�m���/ҪV�\���,M��G���Ѣ�C+yäf=�y#�Uk�
�zo,}��#0����ҟ�������n8��;zV�d�a��,97T�, ,�}5~�Q1���p��ta�P��Ͽ��~��Gz20d��'f��D��;�;=�z^����� qXsQcq�p���9ɘ� �W�S|_��z8���y���(���]�tc����c�7!E���nQ�����v�M��n~������igd|�,�����hQJX�&5�1����߽P�竗�hH��㦓��ZW��7ǆ�qE"���,����wڒ�jF��.0����>���������?�����_�[�MծA�e��[�sw�9_r��0I��df�&u�1�m@�L�����??>�z�����!����em����?�dx('��Ƈ�?d�O,��߸�\Px�+3���A��J�Sx�{�f_�|�dhT�� �蠞�8���P�{����(�İ�i;��\s����ǘ^o�ـH�IV�����L�KX�ϧ�"Gn�)�H\�m�V�I��nL4�u�ɤ�jɥ��
���Ƙ��zݼ~D8ú������F#؈�b��8�� ���#�DA��a��
��>>�n�?b���_���P�;�ϗA�< �����Ϟ���;]�X�s�u�Bp�|E:v�{JT�MXc(�Vf7}ds�0�B�R�H��t�>�oY70���'��B�����D��^7��Ճ'r=��y�Ϟ>K��?�K�4$$�)Żc�Ǫ�	�"�))�$&��D���&3&0eNiQ�-/��씆��?������ﰽ2s�'\�oa�e�`�������I<Ԟ�]I8�Y��cc`�ױ8�m�Cn�s�EU�;���X���-�Y>�G~bP����
�k��$z\#�[R	�玕j6�`h 6�79��\�{]ǙI�q��-�\�$�msDX���iئ�9���?��������Y�~���
�'Qx�����������` ��c�0��x�ѯƀ1�_��(�����1��h�E��&c�W܄4x�aϛ�gPs�ᔬauY��j��`��啛F���?��s୩�^:��`�v�eZm�L������l���~����eڑ��%=�� ] L��2}^w�髯�C�]Y�9[�!����O��'O�pa� V �'N��"S"��bc���jؚ��xOL~,��u�]�p��c�k?��sR���>xh�=[�/��@Ba���]6\�8�n�-���l��h	K�����NQǛ���_Rm���w���\��!�C#K��ե,\S�<C|O<����9��y�����=����#�{g��9ܸ��u�T<Gl�q;ZYi}J����|	$�K�� !`�U� ����	�5x��&�=ǀ{�� ���=�
����1����_չ��v�y���`�F��\"�!
95�Y�A�j�$�W���Cg+o���7mش`N����j�w��?K�[vN\����zɭ�/t���8����gj-i��L\����_XU�&�,&]��W"���_~�%���)(p+P�~���:i��=�yUB!<��A�I���9���X��0��������������T���q��4�;������=�0�eK����$^���yY"m���@�-��/>oz��O���_��P;"a}�6V�/���H�����5ƍ	 �О�?�����'�j%\z����_D 0�0XJ4a��q�0Ѩ����׫����� #���"��c���rS�c�q�\�y�&��>7YQ��]x�8��:��,�M�0����?�0�-9\�)I�׿��B)��VX�&Bd���v�Yo�^��B��;Z��ciB��c���Vӆ*/�e�A9��ӖIf�I3:�D�a��_������äC������8}��W���G\�=8��K|��9aKL5�Cu���X*k��X`�d���jᅧ*B8�Ғi0���0����\��J2R��u\V^'�c�R����|%���Y9��c���m��Řk����f�Ɓ�a�L_�2j=S�$�aԨ��d%��lcv~nb8�`<���S`��/�x�^j���0Ѹ�DUK�̼��3@(���%B�hK���x�	���0�L2�7�d��ܼs�����,����py���˚+�ȖPG)clJM����ךQ�o�mx7KO������[֜B�e���h���o87��O-��Z��T�bb)��+��!��&\u����p/�5'9I���+�׳i���p�y���^�BQ�>�±pyv�6[`􌧦���98�rx-�yM�j��aW#n&�|�ᳰ�.�W#t��L!��둊�k�[c �]���?{������1X��R��P�z��D$\"X������Բ�^�Q�4�0T�����\���@&���܀(θC*6ʕ-O3�9
+�n�(Xh?]
E�����s��0ϺF���s�3�TMᵛՆ��7�'<�z�(�������z�<|`	��c'�츪_��wk1��Y���W����w���� ��2h��>=�q�lj��[^�%S�Q�����0��a�WB�I|^�߱�T>��sz3�X�Gs�&LD�j;z>%���-ѫ�^�����2���L�4��-|�����{z���
�
��}	>�}~�%'y������C%�����y�ej�m����?<ߣ_�
Y3�=��v�؁������48V����I!�M��mYŰiK����5+�.�9�4V�_~���6�'����?���*A��oA�Qhs����"��9fJ,*�+&X�cl�*�&�*#�Ǽ� St��5o�@A����^��Zu��	,'�udF�폃����ti�?���y�o��E�!�;Sy`h�9��K0�L{�l��%�܏�h�<0 ���f�'��h�@��6*����Ù�Jj����]�+BÅ-����B�P5lQ��4�[�F�I�k�[K���`��.� -�^)����ҋ�=A�A=Y7�����c��K�����K�xg�u���,���LB��~���}P����k ����㹣I)��I�KVnz�ST�6��M#U���_�A&���f2/T���6H1�v���iqf�9_&���ʩ	��Gi�{�z_��;��-����X2�W��L�������uz�t�~"�GU��^2UX^�j��k�߻���M�I5�ww��?e��s�^��&�7=[F�m3�t��Bj���� �#��0{ݺ�sX0�h�u��sd=��g"��c�h���ł�|^*����:�8��h���YE��p/�Ax���
甇jB���)xh
/-��^49�9�-���QX��q[/]�XR����?5��!c!�/b�<��QL�1��qn1��+��1�l.'�d��
ùu�*�Hlʗ�v�`��Jx���+�&�6pN�:b
�ձp� �#��!��>�u��.J��e�=J��:y� ��|||7`�j�A�w`1C5�F��&T��jt�t��/Q�!0���N���滢VY��l���S�a�-�2B�[�Zۤ��GY����%�������ѯ�a��)Iٛ��<B��ָ��]�a���w��S\ST���c6O�;1c?��<��2�T��=l���F(�K���e���k�_>'���E��G(#��c�L�ƽ)W�@n2��`���rS��U��	�uy�+�׼�Ss����^�~�P�hL똁�ilې�u&���@X��a���c�q}G)�c��'w�B��uI�`B9]��m�X�ţ�7�+6E�cD�	��P����i��c|�k
�\s\1�8V{ƣ%��:���&C��?�`,<{���L����o�1����m˓��"w�w��X��/)u��S"�yv�@�r��ۭn{ngLU�4YF[}� �D}`QXL4X{˪��S�)G؂y�?��?���;&��e�7Gkð�xpt�"���e�3�0|,QD�~��k�jE4z���ᅡeߡ����������U�:�B֏UQ��'�/G����A�_���X��JzM�+�
�`��i�'���c�����aQn$m�o|?d��A�k�Z��<|h�5��q�HO��q\��3W/Y|�p�<~�.�5�ѹS��F1��z����QB��/�(~��VfjFW�_l�ڰ����+T���Z�`LqfH<�����ƽn���Fԅ��rl|'l�=~���G��\*�.�������<�"�Շ�'��pؼh�i���4���\�9�:�ՏH���'��!��*C|ϊ__^��9�e��b'���aF�J<��x�"���?��~��Ɨ\H�Q�w��p�2�L�L=qa^�5'�UI�+����)mcL�_PU��S�w��NW��ΐ6y�Y>�d���D̗A}�8��M�ӈ��!�]ֹ��������Gt1Kss�7m��H�2DrN������(���k�4��`5X��X����dq a�����ՠ^9���̘��8X�����%S�8�}O��Ә��������㨀y��@9`�2�>��fr$��F�.�#�Ӧ��'/!�#B�65l#���2����7m�ھ���{8>�Am!K�<��)����i��f��0��'�D� ���X0J�^� 4�����Q��']p+e�-;������뀙�=۩����3�w����B��D�hU�Sv��Z	�d*Si��hl��Mň�|�4/mZ�^Snp������+�W����01�r|<�pT�	!$� KL��T��־�/?nZԤ�6]j����.��b��~V�M���X�6�����)�y�J�`,������_T�z���Ye�G�p
Ci��a�,,������ɼ�✬�t�$�%�ګ)��K���=���wf�SQ]2COm��]^V�?��F��b������3$�6���R�@�.~/aX9M�n��>�� �_r�S[��=�8B�;h��cz�;]�K)3����n�/%Z�rB֝���=x�_~�=d2���?�^���u7R��D\��Q~h��S���5�Ƴ:юhx��r
�!&�y�V������k����j1S�=��Ő`���e�װa��l�6UW/#�����<��C�u[��)ϋ����dښ����	OL�:()-��H������qN����E�gu<���D|���?2�"ã�F��o�!�FU8�q2�����%��V��/��9 ���6O.�`Cx{xp�a��r���;��h� �O�<��o���@K,��"uo���xs䚺��v��:/�y�y��VJNf��^�Zb^j�)Yٕ��{�vB�������w�I��^lCU?�i�`-P�����|ݵ�)S���TR���u����V4���Kvޘ�x���~K?��_�i��������2�����/>�q=��L��&w�����e� �X%����)�d��}2Y�������;�b�b�q;v+,�s��z����i��8ۜ1�0���x��Yҳ�=޿G��<)|=�y}�BQ,�/���%}�h;X�����(W�jK�tl��x^2�ta}x��S�j�xt��s����؇�A8�ͩ3v��P���ā�M��Dc:�1=��0�;�W̚�p{y��U���'4����6��g���%ꀝ&��_���3�sK]܁�ð�Gׇ�ދ�]� �W�e_'��[z����i�O���[:Z�9��7�x�F�b�R�//������Xˊk����a�:v�PU�{T�4U���hY�L�,�~�P.�� &: ���}CmW����S	m��e ���>�ٷ�#�+�Ŭ�L�c!~�ヅ�����3�Y`t�u�^��F��mY~?���u�rI.�`��8��9@�◟~J��h�D���s���a<��	
%H�}��W�ޙMH|6 zx��d�N�i��|$���4�s�Y*̎J�j�k�aҟ�;cu����7�'O���T,��aXׯ��уtV���l cs�vOc�IM�`ax��_�����{>_Ђ`x��l�\�7x]�U�AA�F��_�W_~���z��at�VݸhLK����RY��J���//�Q�cl�,��b�hy��y5�?�s���Ͼ�A%��R0��_�����u���dҋ���/�-*�͛���`� ��ōцJH��iQҴ�`��"yz��G� �P0���*�j/�D��5��LD���1��q.1���=�ˋ�.u~-XW���cu..�����g��չ�)���K�"p�^��̩qg�(��U���_�ǳ���:�j�w��%XЎP�����dPs`Xm)��%���Nc���<��◹a�u��ӏ�_��?� ��l��% �d���&?G�S �S��5���=�k���w���),����1h2C���������Q��S���?t1����㓓��&ݘ���2N�N��B�//_Z�Mz\�u�d����/�\���zy�0ԒS�v�yy�ka�XH/��#�|�勨Ȳ�/6�YI�n��v@m�w��M��hwu���ю��M�ߝگ�(�Q��{S�S,��W�=gB���º,������������[���ٌ�YD3��;x�e�),T8�哒j�(��yV2Өw��F�{\=kT��`��8zV�[�#V�Q9*�(`�g�����'��c�q����`a��t�<ej`ۀ�����i�	%0��ުK����,��|`,�}���3���Tm��o��|�O��*��A]Ȩ��p墏?������aЩ	L
8W�XW�����=��{ϑx��C��k��;¸����b|�՗��;*M"I�/���l�WsN�d���z~� @H�٥��k�E�� ��e�[M�,�!y���v�R���V�C\gL{��w�x*ᘺ��`E�{�����Ԝ..�K=G��f������aCٹ�H�"�C��ί���:cU3(*���e�����e�2�ڄ�}T�L��V�J6x�S���X��a�T��/�;�k)g�|,R��N{��\��Kd���vk�mЙ"ƙ��vg�Ux���#�I{@��9�����; ������ow��1=����-������T%��(D�
2�����?�Vp_�u�Q�h8�)�crҳqI4k�'!��Vn1q��hR�ĔZEC��;0+@LF�J��FWܧ�p] W� y��)�mqRE�R֘p�, ��T䵾�r����H�q,d|΃0�܄dp�`��Hz0�W=ug�$)i��M�>2�=���Vtǁ��}�{�������j���:Y>K����5ϓA='��m���Ȏo�C*S�d�3l�����j�a��1e�owaр�kO�����/`�Әl��{�����5y�H&}��~�d�����Rl������l�V�[n�k(��1$7�[BлO�k�!yEW�VX�`��9W��b*XVܠ��{��YMɩU>�-���<T�o���n�v�bn6d;�JS�߻ʸ�U{��9��{n�pō�3ϒ���V'�v���IYn�{�΄�����ghl;�����ڗe�%��ٽj��Ym<x�x^�E�1:��"�#��U/0���x�ꝷ8�"&���Ȉ�]�$����◄�KT��j�HAO<�'������Zi�=1�G��W�Q��uS���!c�1����ppt�vV��=�z����lhC=wP�gV����˦ %���Қ��d�y��C(YὍ����cc��q=|� ���צ��T^����:X��0Γ'�'*�369`�,A�a\�\�f��m����Z\��1��^Ub��vHȋުs��&<M
U:M7���
树��!(%����f,f��"���!�bP�0�����û�-� U5��p��T/31Jv�א�����ֆ�������>�ۙ�@�	�B��pD5�S)�,%�WL>�����bY���D)�1�-N&�<y�p�4fR�����B�'/��:A	�]!�ra�$Ε��J`������o\��(~��\��{��coܧ*mZ}R��Z�=V����̠a�ej��+�� ���RGM�X+�Vj�,���&��bb�WM8ƥ��"�P��8JT�y�4�̬�ܛ��2�-�:��|l�.�훈6-$�pM�|	���^�6]��1�;:���@nr��Oη.n��^�a+��&��i?9�P���+�?⣞�_f�]?��5�C�@ʆI��{���ѦҊP$�n���hשKP��:ƻ�hcƷ�zO�M��},)Ռj
#I����]���ɝ�s��{�\��^b�|�����ce��:���b��6x�����KR���?l�Z�Jo�&��ݴ��������������*���p��$����C��P��n�Ņ0��Fa= ����y蝭�b�K�`PqQ;�Z�6��F�_����yBp��Ņ�Azfz�mq$[2J����G	������FBJl
�@9�v��4N!ai�k���no��1oe�o��rx�}_����J�I�J��Ӭݢ�5��"�`�ޣcoN��fm�WW��r���7�{5��v�q�ҍ䞺�%f��� �a�
�^����ƅyڪ��xN�.�K]mN�5q��}9��!|v���;W�o/-GLחo�d[��`\?lO�[���i2�&��f��\�[<�B��*��`]=5!N�g6�h$���fٱذ�c�-I%X���CcǷp����RO$�>Z]+�0»��:Kpx���ɒ���Ơ��=�R��+l �H�� %���Fѱ4|xhX�ye���if&�S�y�̕�q�9r�s&�����ٮ�P�Ia��bs��эtP94��	�K��
0��6�60I������L��<���<-��d�K(껪~�u:�6�<G�)�З�ð�<�n�[��KS�R��<���Tb������`�D�
�L �'Cʹ�rYB��Ґ�[F-�Kһ�ǘ�QXi*ڷZ���lv��ٶ'y��{ߴl��vڼ�y��E�:>l���94���;~W�p򄌅@%���idm+��]m6iK)hE�)EX�5��iL����N��-t��ӄ8����Ƞ��n���sṺ���^��^�)çE���3���$ķM���:� �i2���B�kq���UC���Sd��1uI/n��\��o�ss]Q��R���C�sygN�U�$y�K#�Pʌǿ�	�E�!�G�3u����߱�險��%q�+Fl��N�ӡ�GԠ�!B{ݜ
�0D҇U��0^8�>��+
�lCi�X�l���)Z���؛��ϭG��i�SҧpX�Ds`X7�0������o����E��ϛ=d�Xtє�t^7��5�ud`��,�SY��Vݿ��i�G9��9,�������fY���S�-�c�zC�:�։�u�!�����P�0�T�N������}I^jx*q����d6â�A=�JL�Ͱn�qk�^�ȫ�	?�!����@#��}��.�)ş��L-uK6��^Y�%��Z7VA��ܱW��؁����'�}, P���<A�����3X�:�L�77���Ux�0N
��Z��n4����dI�ŵ���{��(���>���M��Cv�z��w�� ��J��9�Z@�:Cg ���)7�:�j�>>>�e��x�~Y��!�i}�\35����Q�[�u/X�ڼSa��ԕ&Y��qhÏ�K���G�c�D�su�~���21�r�j�Z4�P�639vmZŚ��<(
(�m.ESn��$`'�ɓ�%���{|X�T>����P�[t
?f���)�xȼw����i`�#1����E�B����|++\y�悲��u�X5j!OT۷+v���g8�І��.@�6(a�wH�EIJN��ʍ)�db�O���wjj�/�ha�7kk&�w�D&m��������~��Q��o�}���oz��q:���cz�2��c��0hC���[�"?���'�E����ƴ̗�I�GۨI��O�׫���VF:��`bq�"�r�+�=P�(54�FI֌l����Ҁ�M��Fl�J5�R&����IW�hOf(�!\M������ުA[��0��h-�I}%����_��'{���ug0�.Z�� �E�'D���1썦]�NT��]Ģ0�=[ԏ��z�C��M㺸'���y�J�H�L���>ΚcbT�T/�xfJ�!헇�!E�;:�D���1���I5�Sݵ�J�I�{�Q{
�3G߽	��.��k�.EZ�j%�T�rd3��8��?3�!��o<!��H<w��P�b0,qE��x�XX����I5�/�����M������]o�DU��=����jY)t���_���a�}C@#_ޓ�؆a��|S��$���˵���1S"�3��H���ySfD�����6Pݯ�Bn͋�"�e	3ۨ%2�"����{	b�Q��N�	��"��Mn�S��`�f�LB�/��X�Se������פG!��g��"m���N��g�,[�4u֕8�����f��*�����e}�n0�8�x��i���( ����1Jȅجl������_핹x��EY	�H�ǐ�����Ƕ�������ݞ��tDx������	�%�O��μ�$�R^PK�9=��հ\��=���(2�Me�)ݺu������X��r/W�W>�e�������'���I��"s���7a��p���n��%�0�li�5��5��_}�T�
���5��]<��'~��ֱ?�Ɏ��{_wc2db��#�=�Z���j�i�."_P��l\[�0[�O�� ���~nZ�֒m�Q�sa/U�P�4zE��'e�@v�}T�)[/�-���Pr�Z���7Y5B���'2MVr����XR�I�V]�҈���ɳ>>��k��'�;�o���� L��lp������&�Y]��K�㫵]���u,��VR�(��]�㡍l����SDtL��(�t�RyO�{�m��mc׿���ν���B��z�~9�͕e�"?���-�KC55|����rpA���B�0 |���yzZB4�������$nUc�)$qx�E_��4-�1y 8�*S#1je�#	�Z��	��<��� f���`1C�P]\ס�9�����Rj1�EKj�/�c����d�ϯX�{���$�#���(�X�U��˙[�Q%���lf�s:��YĀm�H�x(�0���^��c�W�w]��2u�ۺ1ϱ!2$wc��17�c���3ePq��DQc����Ӕ�$��n,�g����j�������0�d�f�3`Z�u��^SLi�M"1?W�b��rOW���2h`pn�%`'��sN-��Rf�I5�!,VY-_��s3�	(�F�P%Z?'�i1a���#�e`��=���ƍ*���rɼT�%cQ��[C[Ϧ��*gz��g�Aw�q��<S$2Vο�N��y�1pF��?{�%<�����EV��M7v�9p^t)�ƨ��o�ؕ�o��o�ۦ�4N�lN�L�&,<kL�c����F,Ta`���V�L,{]�K���� ����� F�c�><"I������~�S
4���$�t��x��6o���6��I�J�G;V��~S=mz�G�������{��'0�8�GT�$;)Ck��M��sPsr\�L����1��i^'͓��o>��S2Jl16�gK JD:x Cm����	\I�a~��9��0��@a�qhדE^��j�,�<g+�\0K`��w��O��(*�7�Ӿ��At ti�4*/R3X�l���H*^f��:��\ Ye����0�ĉ��H|/���jMC���HCtv�����zv֊ow�����n�WfLGL*�l��IN#� ��@m�Ou#<M�?��P����$v�s�n��+��2� F�!-O�Ce-�`F�X�'�s?���Kb�P�BH�Ey��VgR��t��xˏ�>�Is�q-J��3՜�c�Y�Gc7�9�o�6M���K<q���*��F�����J��:����.�=7��a`vL92��宛�h|���I+*�*���!]��m��7���r��N2��Aul���T�JN�a>���0�E����q���(³2X�N�)`�G���ث�(���w�Ԏ�S*�-w=��޼�KtȰj��KqzL���/�/er�� �j��h��s��8�Q5k�L�䔡��jp~�����]X`�ɯZvz.N��1-�)2�2� ӹ�뇮S�\Z�ů����LA͒7��P�4�%F8���z�_�����D�cQ»���n��9igX`�!erK���+4$�k{�LC�sx�2�9�������^�������d�g���|H6nw���CiqZf��\ul��=��T��#`�kOD*4��^��m��H�*~O��c^�fLo���Z�R8?�|Wv�G�eH]?�6!�z�IH�H^�p]nHN%�1��U���׍��I����z|8����� T&ү��U�D/Nᏼ&*C������u�.�ɳ��ؐ�wĉ����b�j����C\,�(W��ʘ����Ư �Li)�1oKB��
�S��-�-^��� 5�_��6��S���#E2
	8��ٳzo��M�����Ɣ��� c
o�����i�徘��9�0�3��skF'�;�fKˁQ�qtx����h�%C�Ҷ�q�0
����7���X�&S3y=�U4��!�h�Z�&y�s�եl��Mx �x�Ba�[�j�l���� ͞aO%6�my��'D9+��jq��Ql���~�[���/�u
�x�nu�VY7�x�NY��%����9n$�8��X��)��$�o��ۨ48d`J�[7S�%�:qP�@8<?���]m-T��Y\~���b4�b�&������C��$�[2�l�*R����5t�I")^�\�\��{�����]�veZM���.±2�w�����K���y|􂯣�
��eM��3�������C�q�V��xn�k�)��s��ޙ����LP�]�!Ef�t����4��,� �1���Z�X��||a�J/!���"���e�Mg���������"�[��h�h��������0O��0{^ +3�r�J�a�J��������ئ�k-\l�E;��c�V��m�1����T1C��-!�>��:C{X���vDN���J���E }ܽ���JZI-��J9v�ɭ�-�dFŲ�r��z�quf		'�_�t�d��/��w}'��r@�k�g���&~���3��=%�Cx^�
0�y�P������F9u���"����<� L���	����[%%�3�����<QЦ����J܏�L �J*%ON�Gn�E�e���w�X��[R�,0�P]�j�k^vNf�����x_���������fu�l����}q��X��.����qC�����
S'�n����)��IA�'қ���1zYID%�0ඳ%k�-�bٵ�ν�����8SG/&�2Ĉp}���������y����Q�G���*�K�{w%��[Mwn�4EF89:�-��Di�c&`��#��g7dj1�����u��D�UYM@2V��k��i��I���M�2�ϲO�ʳ˿��R~�!�X1��S��z庬�������k~`�}�
x���c�=O!��:��o���/��~��jV0@�nL�,�/Kh��+zV�w�FQK�F�vU�<O]r�]ѩTZ
�r�j ���Y)(6
$����!�����`<��Jt<U��Ū�>%6;���R[�!�KP��&B>+��p[��]Ɔ�_�q����،/����
QFO�aSA��cks����vЍf�͆�כ�g��&�SW̑Գ5��Y�hB���6)�i�/B�r�[ݑ��}�1�����X�Ȃ��!Ns��i�A]���D%�gϢ.������Ⱥ}��^o]�ޒ[0����R�׀C���rHyV��	����y�����5,Q��ϳJ�*�/��m�.�Q_���M�{#qǢײ�w��5�}�s��a��ӧ̔��\r�oB���F�h�^A|+)�SU���~�)Q�M���м�(E���)�<q�Y��ݚ1���N�!�n�k�K�X؎q�������yB9V:�G*vH\��	r �f�!���9H�*�X�*��b��ۀ�w�f˦��>����q�1O���� ��0�l��<٦�����i*�L��o^ɖ��V�i��e�WYuaG��vҾkcќ�T�j���p٧�|uƘL�Ą���#<���.��%�T/�R��՘��su���d�*<����ExjJ��S�����	
��e����<C�J�Q�����k�*��:��D,Յ4`X=z�.��G���yV=�Ǐ3�3�&���mh�:ˁ���˶��+�������y�nLSK�L2���Kd� ���;�G���mF��_&zp��Q��9���2|.ǥ�g5�33V��9�*�@�nOt.� -�fΐ��������sn�}'i���G�3#(V���d� ?�d^�e�EA���W$&�<�C�׎�S�/�F��H��$�o)�7<G�7K�ۢ�eLEYi����2�����Yݦ9�x��l�d(�G����>��F\�䋃��j��%�ϋZӳU�>!�h9���짦u���)���F#���R��?ϙ�3��i��`�R��R�_!Lw��)S�BtM�@#ڬ�J
ڱ�� ����z��Y���M��u�"yny�m���?�΢{@Zn�s_�SJ�~���Q�+J���I��9��O��7�;�\���.�;�tc+���0�x�57m]��L�HZJ�������ͣW�Z2E)���*%
X�z���7��+G�v)C%$��O����ĺ]=+��Q�k�@s�=�;a�|���ߛ��H��*�S���ƹ|�ﲞ�H�݋��pW�ǘ�*" X��w���d!��Ah�"c����O��g�����w/�p�����}�b�����?#ކ�ޡ�0���Ķ*Û��A�}��:�6y��L�j�3X��2�k�dF��I�Q����	r ���YuCɻ��jH�alè�__�L/�� /C��jt��:�%��(Uw����;k��"O2�-'��e.*9ԤYF!Q�8䀏z6�
���d�G��J�E�bI���Ȼ�q���Hv�?+|�j ����N'~��摧�L����)r���F\]��D�ֽ�9~Y�9��W����I��!|�N�
%�!�V�f�yl ʁ�4��V��9�JDC���+���0?����ߡ�6$À��6���'��dǎђcy+`�7�K��@ļ`�\ph@�RY���A}sv.�°���Y ����c�6�W�L��R;�]�4w�i�1yPCN���{�����嵵%��2�$Lcҽ�d %��Yy�o=����O�s�"l���pȗ/���'O��\Hr��	�/�0�ae&}��S�w�~R��C(����)�7�(m���(��N�CbF"j�ih,d���6-HB��r�s�C)ј�N��Ӏ�ؒ��n�Fq8�-�6$C��1���%_�%y]m��n.�k�x����엋�>�ב��1�^8�����JTq�8��B�x}^_W�?i.&�S����k��>}�Į{5�(aUC�k���{�X�6iܮ��$v�ZEI�w�8�T��vrM�c�������z�����AQ�a���H#�8� ���z����������}@�zAg s�G����D<広�""Z�PM�֤Ri�J"sۅ��%����X��n�%�~������~!���X��*p���t����b�2+�a	�`��UA|�ѪX֙s,Rx/��8��\]-u�(!������>wa�_��XBcb��>]�X!�&�H�}����M�`Pa��8��h�;�G��
��8�{O�`a�mYj9�wl�c#z3��g
����&������~���r4�Sh���b���őc#5U���G��v޸�ղ�}j0�0F7^)7��`N�59�Ʋ+&��:�h{O�U�mo�7������N���zf��VԘfp.c�Ę {ǆ�β�R�8>�$^�i�nPw:+�q@�3	%�p G�u��Y	;�#��54�c���c�0�;���+��J����g�fw�0'��)��hD�=��f�Qda��|!��R��U<[Y���jod?���Ը�X��ü��e�8��
1"\�7�Z��� cLP���ϡ�����ie�!���o�R�S�x�ko��	zU��N}J<n�./7��J\CjF�[iL��:�$Et���ʵ7>[;E��<9��m����{���{xX�ۼ5�#[a�a�����#F����ae-S�'�L_�U�y� �0�1��u]x%�6�P�V����']ڷ��  u�IDAT�mY�o���K^�u��k��'kkJGLy���9gr�T��}�5T�i	���J�qt�p��6��D���9%�u��}���^�5�sk�b%E^�7��6P���6a�Ѫ�����n���%07¹�gƆ����R��M0�ޱ�[4�fN�W��S�"Ӆه�\���QM�/�uh����1���(K쇭�.1�%�]9��n���1z&IAi��j'�%m�5��Ϟ-�:��[O)�a�� �	'(�����K-!a��UEȞ����m�ZOsQ�����!��E}���}��
g��h��8��QQ[ �6.����,q�-�b��rN�e5.��fD7޽u���T�䏦�N���~/�E/�=�D�����Xvp�s���3�en�����#����$W��w��6�K�!�pɧ�s3<;��MT�tU�!�;�J�u��rcqX��3��K�=��0y�ɡ�����_|�%���dl��m�mj�|��.�E+�"�tq��W�q����b〱D�j��FwS����7�>L�]!�./0D$�X9���e����y����E�1�2���T�%.z�v�����.t[�T�#�N�3ǋ��UkEl�L&I��n`�V�'N&�D!3����7�K���l�c��?f���w}��M��=�[]�S�Ғ��|�����$/f�6g.Nqf�^转��U�LadI�)������זD����=�}��w\K#��"�L����xڡ�Kd |�/b��I�S�e��|Z����CR"�������[�:���evHu�1%�=E䂤���|�����?<���_,ǵVݫ�� r�ģn�Nɓ�1��m�Cr����,lH�B�s�>x�0�d���9��}��l]�1̓������g\^���ǕS�t����H�wڊRH!rsq�X��al%���U�R54=}��&��+�a���q|2�J�qc�ia�A-|T�Ju�b�S��@�:>9J�n"0������lB��3�k�aW%?^&4R
/�	/�Q�_����
��z�-�޻������(�')q
}G&�<,�R�����'��ʦ���DWTӼ�J0,6���]�NJQ�r���v2;]�a��y|p�X�6a_vu�R����.ø�Tm�}�ҿ���T3`��W��i�u��_*P�����v����g�>K���?�����E	.B���<NW+�L$��7l��a��=8�T�o�n�g�~y��^�y96;�����pup����ztie�`%T���ܒ�����;�x.�Ga��9����kKJa~�S�>SS�����A-���q�����bg�`ebnT�w=b�������1��n���-��m�C��� �E����;f^g��'����ⲳ�ȍ <N,H�Ѡ"�c��\�C�yժ�f�l1�SiF�j��J��6&h!����"�f�W�:,�|޹-�}��7�SRk ����%�L�`�.�a�,���7o��^
�F&xx�9X=��c�릑�����og׭M�sW�&�u�9ځ���[K	.r��c�x�:�m���!q�u�8�ǖV�A*���B�~IC�D����N����~���K����O��)�c��:�U17�a�)���M��YWn���1d���ȵY�񁎥�w(`S�V/�/��y�������ŭx4�s��;wa�t�u]��sD&pV(R��M\�a���?��$j�>C���dE���+�"�]"���a���_�_,B�n���qgJC�C��ݚT�:1O�����w��ێ��� �+T���P�uU��a��*NX?�
�|Z'�#�u��ȣ#�!^\Z���ΰ]d���pY���{�
��v�j�*F���?YV꺝;�lyRcsD�`�X�ֆ��1�w�wZx����x��zh<5�w������ߨ�[7�S�J�
��P�J0���R`-?ʐǱmt�O����1U
c���z/[Eqý3�ĩ�3���+7x����EQ��0B�����y��O�)�qP��)p,
��/.:���qx�J(i|a��Qn�0<�:>�i��*���O�䚒T��@Kc�-� ���"�C��R�2�����8�t�$W����5���IT\WZ~�,�n{�zWp�3�Ɇ�=�1}��j���o�!B�ao���3ǲ���/�=�1��Ļdz��!�{w�s$�����yP\Ҥ#Mil�E�ڣB($�e��?qF&1��e�,X�y��K��X0���#�V�]�~1"�b������e���v�3WAwṡ�^݉����?���{�A�E1}㝶k�F^3^�[ꆑ�0v�?G�jI��`��^�m���gw]7�����Y�Icؔ������Z��cC�a6H��3�Ք��I"��s������7��\���O��Yy1�nm�ܼvË��#���_1����c6�$4�a���a���*9Ĕoi",�ڢ���M����GMކ'�$s�)�PV���8�@IԹ�ǃ��b�D��^��]��#uc����_||2u�����; mhQ9���$���i=���CR	�ї�_��]-���J
��<s!��.Mm��	�X�]��H�",��93Ϯ:���4��U�X�j�Ke�P���?�Y��\�^��W���W�<��D���<~��]d�'d�'f���	s�5������{�m�Į��h9GG'4R(��u=C�Y=4.px����bj���7~�iP���h*�kh{*7�QEf�}�ZD،^"�Fc��q�26���]7���S�m�S_WJ��_Uo>��9�x[�^I�������ù��ECG-$��8Ys�~�����ϿDe柕���([�36�5Bq
Qb��Z����qQn��wx���Ob�x� �@~�^�d;���W^��]M��'/����S�v���a�)T
\z7��T�.ޫtF�/>>�Z��Het�e���-+�E�W^.&/k�!��6}���ߏ�2L�Y{+k[eS�G����d�V�V�-y=�	J�P�)�V=���5���M�ަ��j��ڽ�S{�ㆷ�P	�*��;��<cѱ�o&`U1�/y�Ź�������۪�ۺt�M�jvpr���x�ɹ1�OaD�-�3��(6�.�؏S?��[��.��c�cb��e(��8��sqW^�i����3��^["Ί1�C5�q��:~9���-���B���&�w�9�Wt�!0�]�&�/����WUn5�?��on�8o\���:�	�Q����pڋ��_u-
�Z��5��Ki�R/,񈹂s|V=d�?5>6�r�.�y���+W�W4]M�C�;k������Q��g�������Ŝ���c��P�Bo�=T���Eb?����M�����-���u�H�xHF@����ڥ�^�� �y;��T�]`_X Z����K921,�����S��b�n����;7FlO1x�� ���k�}�Z3�� ���f۠�`:m��ګ$�XK=��3�ȣ&L�P@T�̅a�zc��V�Wz�&�gL��8
|�U?+_X2��T;�,�U!��bF�ߟHj�b�LM�^X(z��ۃQC�¤�y�(�m:�X���۰h�ph�}���#�CF�T���D�+��6�j��񔉬�f��䑅�
�cEDc�U��Z1N����y����\��ʐa81�p��g����M�{==�e@A�/������r8����$ab�5,Ugޠ���Ko4ǺV�%��ֳ�TO�f�����������a��s(��t_s'��_�T�¤��d��>���A�����堓m<�b!���ρ�!��n��N2�~�H��
��*\�k�k�^J�u�]qIYai&0��عOOΌ�rte���{8)�R����>�yW|=8�_�5=x&�}�  �+��^F��	ҮD�8��$�ܳ�"���[�����,���`ԇ�<N���+�q� JB�n�F� �>*����d�uLe�六ʫ�<��n0H[t6>%z-��q�Q�9&n�+������*��&�2N���sv��Zv��k��>�o0��4h�^�R�+ֶ]��T�f����ai���)X�Gy�������ֹ���]p=f��c+�H�;xg�q�_�J�dW�\���'�ކ��k�X�c-6��D�Y��9���(Rɭ]��%��>rRKD)(Y����8a�o�c9������M��8�/j��p����a<����2��/2��&㫲%��B	'7��������JI/��;�0�\�$���\��t�x�� ��z��٦���ԛ�|��hܤ�
�g�O���ɓ �t\ptL�3��P�hԖW�!���+���k��o2`��0pX'#{dm�lT����`в�H��|�`S���V<� xM�LI�G���L���!x��Gy�1������b㾌�J@@:�k�r����8F�A\�������� ���K��BO�C�ժq0a�؛�n@8L��� �J���96m�de����E�Tr�s�(�M��S��8�|F�Q?���Gi��57���\ .
�U��$[Hml�.��Z���cl�>U�)���(�_�.F^�^ҒP�^'>��oʍm��SG���Go:��;}�(��1iX9��_�~Z*]�����,%�}�w�����0�R'<���fP�DC��2�Ԍw��W�3ݸ�=�o��B����\3����zut�Mҍ���㯣y <!�d����xu��`���Ħ�Cfć���f0�X�3���3k�I�r��ex�{6�9��8�Q��Bg�)3�G�[GM��K��j�lR�Jf,�KܴM!;2ÁaӼX`��!��o�	�@7vg���筪�*},1�s&�U��ݻ�a���~@*�ސ�8�+�A�<\�%먔򨤾�,���:Ȳ���FL��%��}���:���sS��7�^|�5�����&�C�ȫ���țd�2�{���Źy'ؕ�jWQ��c�)�5��!>/�1:�z�����A�!��7��v��_"�b�&���%u{zM�a5�6�Ff�>x=V��B�y�.l�'U�jx.�t-JH�=$9!*M�����S��sO��� Bhx��:#mI�C��^{��X�	7�����y�h �l��"��&��8����
#
���{m<�����l#�s�k�V��s�5���nY�Iy9�L���z�~8ۇ{����4��ԣG�.�C�`�#��U?o�-#'O1T�`��Mk�����we�<DT��b��1|Fd��*)<O&�<$gAȋ�$�kF/U^qc6=�GaC�;�����]D#�K�]��Lt�U'#����ykj�Rx|���b=��r��Xl@yr�T�Ul:� �xhc�G(I�fi����q ����q�d��A��y�0 �,N-|�y�^�.΋2�jTO/N�㶽���e�U���(�0A�+��*����J��O!t���}�p@�v��b���q�_1� �r��".4�����l���ɱ`,�k�;�J�cu/��τ�ޅD���ܠ5�3~�)3�N���*���W݂1��u5�D���	O6��6Zh@��]H�̱�#U�-�S`{^�̏������K�E_Z6;k��������++����Ɣ���V��񑉱�|�6��}"!Ai��2e��Fc��®���{E/�(����2���m�̴T��� �}�^�*?�Wɡ��
�^LcL�H;���� �r��U^m���(�@�`9^Q�z4��DT��L���A�I>�0ٔ���)<��u��/�e*��CB"�N�X��N��S��[MY�<A��F�����x�z��y(���IJQC}�-��O�~�K
ϋʙ��DL�_�/KI6L��c��fU�0f�l!����-�xΓ���"|��q�N�0��������z�=�FFD'���w�~=_z����\�[IO^bp�J���+���^�we?��ǒ{��>����).�\ޮp�P��X�)ެq�Cv�:\Su�=���x������w2¾���K��νX���|��"�禓�J�B�{�^�'����$$����.�ub���S�
=У������svͰۍb��n\�چ��j~Ҥ�֞�� �l�/�5���M��F�ע`�����4�e`?��0���k���9�Q[�Z�j��mt\�j��H¡^=+��`ܻ��o��J׾��]�iZ��<;�r���IZ�F%��`�G �!�U�}��}�͔/8�f'X���3Hz�\[����	����902Q��F}�����ƪ$v7YR��5	�a���6�{��?>�h�}��G�C�E��8�9��ql����ϝgS骃ɠ��re�6c���<Ӣ�sN��t���������v*x �2�l��Q��Ǽݰ��[2�*���[]�B?Bj\K�<N�����U��8�9�`<���~�š�ϢoOz�`n�]�#������s����l���!&R�� Pay`�*�EF�Ԫ%|��D$��sE��;/6ەws`����ӂ�C4w�~��'aPq(䋐Pi|-��@�g"�<5"�{������Z?��0�TD�]Kq�IS{�]�O����[���p�6T������ ����I��5�n������#�}�a	6�l�j���l��v��U4_������C"��.�kx�p�{���d�����Ttk�S������1�y4aDs7�%�t`$�p��l�;Mͅ��$�=Q��Y�<iP�u�m���g�Z%O����i|D��<k���GB6�NK��&��>~yl�=5y��D���(E��a�սO��к�bs]�ˢ��e˓k/��|�#!|�kcfI&���Z�x���6�Q�H�m9��7f�� ���M�����e��>|Տκ~2����L�})p�¹R��Y��r���ν&9��%v��(�&�s`�l�|�5�G��?��e=��62��Վ��K+Jǁ���θ��'���QCS�WKe�X�����-k��Bf����EDE*���ʓ'�1�x>a$=���t���j�B{�LJFD�C筈#�d\[	��wY�ҩҭ���QnbC��D_�'��-��ʆs��sV�g��s�;t.+�@�
?Gy�����;��l��u��GP����̔܊��j���T:�������߃A݅.���~g��4�{���{�I8086d|�w�hn�;'
Ĭ���ڄ�����#���;�#'�V��G}��C^l���5}�nj�#9>-�څ#]T�|�qݤ�D�Z'�~�oe�|��S�Z��%�Gi�rg��5����8��j*�ٽUw\yr4��l�.�0���zx�!5u���UՉ��/�G��C��p㸁�#�%*�
��Ӳ^#k�q�
�By���R�5��ıɃ�nH#�`x�B�l7��Gح��e'Y�ep~�X����V:��TAR�˞O�l$��O��}�ز�~.�AF)`zԍ��7�����6A�QT4O�'���=r�,�@ˉ%x�eA�|j����]�G�(��/�md<9�ʅSt�A��ì��R�Mt�i.qpE�/��t�Ԋ26\6_�	��p!��̍$¾�c�h�}%@D�Gj�K�܈.M@�}l�iJ�����;��	t5U�w�>�l�w���%��2���Ȓg!	���&x�&D�)4L��@��1���4f�ܚ�U��Ty�p�h1T��ٻ|Nֻ����w��hdj�,�T�:X.��á��6`���$šl6Z@�oI������/5Y6��K���K�}����Q���H*Kc�����G�N�6��rj�hc�����<<_ն��)��\��D^�B9��lz��5Γ��lFr�����MyW��\F��"���"����l��ޙ�cG{��rS���>P;�
��^� �D��
��׬m�ױ�F�B)��g�+ˣK��a�ᴷ��Ey�����0���ʟ�|my�ؚwjJT4���V�?4'�ϋܺ����OƠ.��rn��v�a��[���	2+�Q�H$)�w���IT�=�4E����
�j
G�kGAv� ������@�+#������%��H�P΍��!L��:u�<��tE�W�I�HpqH��=�g�~�2�6��y� �T�Q�N�xe{m,��=������駲X?}8�~L�"4��}�!���6!n5�Ҁ����Af����"�<� ��x��a�ƩnN`U��4qC/�Lb	8]M�=�s�1>�@o)�g�z��#&q�+/ع�8����� ��zU�~��}�.��ՐD�"�PLMl�mɩ%�J@5���9i>��EMs�K�U��Y�X����E��[���Z�0=�����k�jP������B
}������I��xo��`���m�=,��2�O(;�wQ��,��I���הI�� a_���{7y7H&�'|��Ԡ���SRK�������S��<<W��8s��B�٩\�<'*�Sk��Α���z��2�c�f/%�n){����6�ka��Qac��ƚ�U�dS��ug3��5!t��5{ge�,�{�~i 5�G�K�`�-�g����q���!6�w��;�4]�mn�P����y}i�
J"RHĄB8ր���݈ԥ٠��P�0���-d�M��R��F[n
�A���^���%�K�Y`�Yy��!b��W�]�&75�F���z�V��
(
�9�0xuĒb⬃m�6��[e?j1'%���U����"�0vo�8��F��G5%_8�j�d��DZŝ��Δ�[�Aj���7׿4�S���t8��Fև�Ss<����-1���KÉ]u7р�85x�G�|���j�cKT��Z�!�������4l�2QS5��I�R��

�d.�����ў�R�l)��񺐜��Ǝw�}rу�Ҧ%�ӖL�O�XD�\'�tou��W�bE}ކƖm�W��
�pEo�Ǎ�;Xe7�u4kk�\ťڼ�ja��M��Q��Ҧ��+�&ו�̠���3�������(È���1��o~��*�6G���Ş����m�[��y,A�v�{f�ٙ���og���׸ �d�NǱ�*�N%�u�x9<���\?<8H5����#u'����|M[����l5�����\��M���_���f��iΰ[��K%�*�����$����-Vh�R�[d5��b1>�E[D}���t�j `lQ��U��ށ�KNX����S�7A��$����	:nt�--2�ޫ<����!%0�O��s�ͺ����vj�=Y���m�"�KE�D�*�P�t��L����"�O�JO;l:�^�x�3���2Y���S�e�=��̰���3C�l5� �d������^�1O����04�8ozB�����_�	���4�
�	�)S��^�X�g��"��r	���.�������8��L�(E��&	��~���k�.� �t��i�i�#����Q��I�#��M_-�O���b�$�x���r��;����
��͐Fl3�1C�VL<�.��G��{�Su�u�^"�䟶ۉK��d.S�틿4�<m���[�a��c&��t>@���x� ��	7�*���}%��>�L������w���T$WPqmJ����A��N4q�W��B0��VkQ�s(���&4��uGl���zx��Y|�2�#<O�l� d�#�BgK,&�;�w���_�C,��q��'��$��5��Z�w�I��6$�z0�iF-8Z�:u�V�v����R�*�<�&��)$�W-�⢴����⟡/����6ʋ��wyW�f�Tc�b Ǜ3vU�hnn��1E\�,�	���60����Y���cf�`w�xpB�@���g@�,0����6���B�i$�9�9�F�X�����U��ŀX����0:ɯ%*�?�E�ڸ��Q�Vd���ǈǛ-)� '�'ASv{�`ߐ$a<6��RL���$V�$�?\~�� �n�0T����}��B_;$yB�f�2%����s�����G����Z���S�j�8P4Ip^f�si��E�Kq��PƩ	�d��I�tB�kA���uŲ4öՕ��^�+�.�lau��Z�WT�u?�b�e��4Y&e՘p��~�ѧ��dV
�Z)��f�_�06���\价(a�ű��(/ �w��w�|j�f$�ۙ�z>���O�`wz�m��{p�!�'��؟������ח��r꫐�4��5EU���($�N�m�ئ����xN�ĪVg�t��_�f�z�sp�j-v�M�4��m"*�9�'���*��D��I&�Qo����aoyd},�^�$�	�u��U(�[��ȁ^V���,r>17l'�탅<�)���dWg���!�lHWX��" ����z���+홹pNw�i�&� .k��.�Ƀ�D�710hX>�f��,�bA?]�lS ˏmS-&��r�,5Nx	Ls���X��E8��)�g�4mgLJ�eV^h5{��.0��>:$LU����Pw�1�����g��m����-v�HhF��f�O��ʂ�p[.g���qr��U_I����w����ձX� �(7�:���+��鴖-üh4b�,���(�^����V3J��dŗk��&b��!��kFYiuw:/���!�狏�k0H�ML�<(���<N�J�A}�����!.c�4��Q������Y�̖_q9*>�ePUr�f�A*����[x�x���G:�/����4`��<�%6��[�+�j�_�9��ߏ-���_��	 �-����~
0C�A���f�A�d���WSrϛ�K+���T1����)�H�{`�m�qCvn\��Vo�yŞp�D��y��b���I�=� � Y��]l��{a=�HH$���S�1��b k���mk)X9��E=���e�l�t�2���H��Tӿ2C��R�䯲 &bd�v�ߜ�U���`��dÃ�}#�;�*���2�������T͢�P�ֹ.ѕLx�Jn�|f���3C��j����P:��M֬�l�j%�ݎmEe��ƕKٷ=�ῩF�Ӽ�dos�[8����])�v;�����
������d���aAd��R�x���j�?Ҟc_����v�S��k�ò����Q�7�Ef��4|;�0��n{sW��_""��@L�ӛ����tp��f���n����B?\��k�.,�Am5�`!Z�h7�N� �M�cv�Ϝ�_N߳7\�t3Gxopq�j"���?���|J 
�9�da>1�݂�L����I�+�(�������e!�ǌu�u����},�N<A^44c+цYO���̓�wF�ب·�TG�o�����]SI=�uⓖ�2T�7�ek	r�i!O_hb>�� �N3P�}�O�V�ک��^���֎+� z��;X+��XgƁ�g��ǝ��2Ў{�f�zZ������bQWs}���<������<�����]ξm�ǘ"jLV���#Dz�F����#��:Yw�+�J�3�(��{
0�M�wh���[Ш��K%�)�FM���x`��	�k�d���|��1ѳ�f�yuc'/*��斂Q��ٓ� �*�Θ�ϛ:T"9zg�LB0'�c�`=�
0U/��X��S u�q�Ԩz0c������LY�T�~ɥ-梧��)���B�u1$K9������Yvp����c%�p���?k�\�@�^�=W0�4�a�uߛN;���q�F���*��` ���A���� � �b��P5`:��� u�8�<^�Ytu�wd��"�ۻ'6��[SQ`{�$m2�N������?����H�uc����3��Z�8?�^U��ș��Cz1��J�9Rq�Z��@�KE���OF���X�m&���F��&$�O�Ќ���I)��q��Y!#�4����?������Xʿ�X=F�e�ǰY�_/َ�7V�"�[��Tc��j��B��/O/� `˔\�N��'@��\�ĝ,,&Yp;����� �ܗ�!�dĢ:Sݧo�{M�.�%�Cd0��+�-���z�<f�>���s[�!��������v�E)��\�
d^��MR�2?v[$ql��9��-�U G>'Յ��8�H� ,�;�+�۽��ǀ��X`ޝ�4R]��Ì���Wb�U�W��ˍ�{D%�]�ٮ�^U�̀}#ޡ)	.d{3�E��ߕD\}��ʰ���XT��CC�� ��6$L>^Lwf'B�j;�f	/��Sr+�􀾡d�5�Y�}��o/ [r���b �Ҧ���٬��n�NY����� m��r���O���NxY>Gb1$�!&���֗:�l��>�YƇ�j'ڛx/?�d���Jemx� J��jL�8�U���SjRzU���qvk�` �'���\�)j0���}ɍ-�Gs&�C7Y�;�Q�jD��&3�pY�Z̚����z�Rk�};CĤAO̐7�@����\f�}y�]2/�1 ;dД���;E�*��!�o6�w^����[��ۙJ 9j0�Ơv0��U�AU�"3�y ؘAI����OLNҒ����r�� ��U6km�j#�d�8�p� n�д��gQ�GT��;��x�Ru	0�9��{���ns�]��[�� \5c��߹�~�O�((b�`�������[�f�m�yF��l���q��&Te 0�Pe���:�ج�{�7� �+�E�Ɖ�$�E�3>��O��-����E�2������W#�S���Źjz�7�$�A�<yP
�c���G�L�*M՚�f�����(��l��{G�"F4g�co���{���@դ�.��Yx��G��!�#".�ȑ�ESj!�U�5�9�-��{g��nj��`�$��?��z�0܏��֊�W**sb��|���at9X��(� ��4||1���'GE_�&��o�}�x
 |�����v�c/����]݉Z��n3V�0�	Y/
0�l\9�b�˗3O"���Y�������,��1���A�j����;��۱�\tʗK�LX
q�nfl,�Rku�kf���!�����,b��H�4E�K�Np�E6@���kr\��4.�՘�.ތE��"n5�����Q�P�JͣI�^X벘���b�u�`�����dg9�_^^�\�9��lC%O���A����r��l���� �(޶��$�C�Ӎ�a�>rY�o��n��b�������G���_�A����Y��,��6�������<}�I���/s���uz�W�[�C{�6G�u�(�ኄ�} u����}��X\�b۞�o��>�/�Z޻�U���!����֣�>3S�/H
��d��!UY�T��0 <e���\U1Jw:�b������1TŻ� ��F�s�U.n�!?U�d�)k�P@UPL��|{��n*��\%p�2�_� "�.rA����{����y���xX��E�X�-Vhe�oY'��� e����5?�!�������K��YE6kwnD�½�Ō����n9u�ɡm�30��0;��ڒA/����޴�8�G�-dU�]�|o&~.P�^H��96K� �c� �X\c�z���v	��׿|+��#�+2Q��D�W�Оm��m�����%��Aj��ҕKikqN�[\�]�P�خm`����Ь�{��%[������s��\$���"6��:!|��:��Ӏ�1u��S��-��S�D��~��T�ln1�?�͍ ��X��z�zU!�=�?�Y+�L�8�t��ۊ̮RpO��A�M��~�a@w��e��l��T�)�E����L�mh�W"�����E�c�ڤX;���,�����=�=
��L˶[Rk��G�j�A@`	�<�np@�d;Ih]���Z�%nnֱZꔬ_Ƴ��.b�]"rT#�oF�2~� �h9�+��{�?�3�ܠ��x�Hc�FB�ga����O�c����P-5��;�Fױ�������+����|eU�X�vB���uj)�E�r,f��I�8�\$LB�\�<�A�M19�Ų��)��O0L�HE�7�K�����%����p��dx������,��"�[n
�=X5Z���S����08�0��ѩ��y;z?��ҚwFk��Z�=L�]$�+cq����V�2��Mnu�ķT�=E�W�q�l���	����,d�ns�B:���,/�b�7K}x{q���&˶ ��ٸ�{t.YLw�ܰ��VS~����Le�����4�q)���c��j��'t�#�/�\�X��"��5D��WT|:a�$ˆI��,��M����H��u��xb1��*��ѦΡ�k��!�*���~���(�Z��s��RLu�wBJ	�1]��bC���ښ�0���������Y�;Á՚��iP�|���z�$m�c�{>R'��!��<{;��8]T�+������9�����{>�fXDE����u6�'��kI-���0(��i�S	�㩽�U}� �"\�bA_#��T%D����l�n6��  5�Ֆ\�?g)}X�u�Cm%D2���?�9"-5�=����
�����~���:Se� �)ta��x �gS���u�\�XFVæ���B<���{ ʒo4F�l���}D[��9����4�Ё�:�>`(:=jjk5�7E~>��a��^w?��n��Ȇ7��G�E��'�KIQ���b2�B��K���j��������E-�UE͂�(k5���	S���,�|C#���k�[y�(�i�L��]�$'������ܠ�~�$�������L����J��FU����Ã������5U��E,C>"u�i�%�SҠYJ�*0 S�u'2�֖N�Vl���(L4��Fjb�<N���Μ޹�}%r���Z���
FԠ]�1ս�0��,L�J⃤�������Y�>�n|H���U4����QWx��D��0P�� 2��?_�S���dY�K�%�g��-ʐ�MV�����5��`6� �s_���>@97 �~�h`�D���F���|*��]��' bZ�k�\�UR�o�����T�!:�y�6�AaclQ0�{O�oY��k6q�uFi��l��҉f���f��}�d�P[X��.X�eҁݒ���sd���х�K"Y0Q�g�]R�o�>m'���9ϓ3�QW�~�{ �s����Ѭ= �8��� �v|��%�1�<��aq�p����7�L�t�19��ۛ.��[���^;���h{��'l�Hf�Ѝ��:oU+G<ߒ���[���iM"�Xͬ�Z`�
i->bh���s����Jk u��nY�O�~1&I��K�@ߝkϷ)�_$�$t?%��'U�X��7�hFGܓ8�WK�+���j�"I������ox��v�z/-�d�V��H�̥~v�p[��+��,3�	:�������*��n��Mk	R�����O+���*K��F������A�Eފ�!h��'�T�ݴ�JL��.?�H��}T[�mR��OX��O�h ?�k��6
���H"g3v9�zZ�ɷ� � ��H�m�O0b׹NC�F���G:ïQ~m@-ɲ�_�{J1�Q���E�K��)Y(=���	T�[��DΨ�8Y�J�%�ݫ[;]'�wH	�����D��H;w �����jz-(1(X�MyVIe:�	ѩ ����ڔ�۹����X.��M����z<Y*�[�TO�Vr�_�����%��t��7H'�9Ö T����ƣuu�͢��	*��g	� AAn�&�P�v�K��q:��p�d�LAO�C��5?�7�,8|EїJ.�(Ā(]]���jv��v� L��J�n��J6���!�l��r�%��ݕ�H����'>����T�LJ�Cg,v�u�U]�jS].�������Ez臷����r��/*G{���R �!���A~��4NN�0��Jf��u��&��ug=��>u��;�j�=/������x��~T�Z�F��*˞ ˿nȡuQvUM��N� ���E����y]��z�͇g�g��9�Cc_���v��B���9WG�b�u�o���6���V��q�V��̫��3CGF�CG�Dׅɐ@�E#��
����6Ɏ��Mѿ�΂b���"a��D���F���S7z�`��}[<$�Tl�Q��ѿ����db��rdv�M]�{(�T����32#�7)0�$0�,��%��fJ�Ek��U%�N�ۦ�[s2�$!��#�����ܧ|m�V���ΟΏ��-�UUOhc08,�`��X(�C?� Ms�=�/���^��.��p%�	م,�;r��H�@0,��wb��t�C˗1�\e�J7��Y��̙���8x�]�m~Q6�� �ј؊VF'�NW�i��e:�8t�`S� �Ha�K��l���fu�h�'=�#g�(T�z�Ƒ`��Y(	�~,��Z��~\|G�X�l1ӻ����ġPo��s���p1�)��h�]J_�ģ�y[�wO�[�]��~�v���q����4//n�K�,�M��DxE�`�غ>���!	��J�w!ڣ�"������>�ʑ#*Y��S�q��BH�6�;��
0�\m�^�1x� GJ�3��T��;o��=t9���Y��0��~�gK���k��lT��w�铦�������x�Yc�$���sعC�l�z}{����QZ�L�r ���ە��|J������{tK(صAFn��h�'s���I(MVʉ�,��n>�tSn�>E�@ީ��|�q@������l�l����4@�j���*���uꟗc�V3r�͖׷���[�-�H�"��@GNb4�\0X u����nLxPk��ml).�����;�g1�bǔ/�:�d:غ���#�g"�RH��ޮDp��r��^�_�%IcA$J~����3�5��0mgNn�&b"�TF5@V::���Z���k��Klf���܀d" E�d�3ؔ0I�Z�@`wΏ�����,�� �(1��!���F�spI�:!J���<y�XOA�D��^��ܗ�oW\2�������_:���3�,�5����:T�'<�l�!@�h����DrV�D�?c��o��ژiX��u�b�����J���/���ڴ�#qp��K>to`q�y,z��ګ�J�F�T�
߁)��By��/.��)�`����Z��Y��E���F� )��[��|�&;3M�&��� 0�\��Vb���ٳ8-�gjq ]lv�>�,i f�@i�A��"��a?�`�8���Q-�vbsVzt �[�"b=yY-������2� ��1K�\��s��fR�&�[d���ϮtOxH���V����ڻ�X�~w�Q��Tk<Ìk�ހ��}k��x��
ʞ	�Tn�o���z�ӁiX�F+7��'���g��G]��d��Kr�
�h���6�eB@������( ��ʾ���In�;�j��,2[&�Llt\�T�2 I�b���τ������U���q]���q�$�T)�⦩~��ӶqS/�t����N-���.Õm=�&���c�J츗�Zԫk�[�=��U�U�J��L��P# \���v��w<6���wS��<Z�[���㯶ɯ���2��.x�y辫��0��&��`*]4���ZF�3��'w��X�ͥ�ں?Eq�?HE75X;Ia��r�]��RR��T��5?1I�fzp�S��?2ԩs֏@�.m���Ń���;��֝����7����K�2�p� .
tD���>�01�Z&��+a������y�,�ӧT�9M�l�ce��uP�C�:�1�-�M���x��C�O#�z���O/�/�X�'���
OR��!�{�n��dC������>�����͸7�e��D��^�t�c�D@�^X�C7�b���-��3t�C6�Mf�#�c 5�-���'�n��ɐl��v�*����; � ���!k`���?���*X��N���d@�	�@ߏC���').g�0�.��H�wU��W�m��i��0V�l��[p-[WF��z�G��;��'=h�������:�r_�2�/F?��z`��⭬��*>����6��^ :�� *V� �m��?���{��� ��~�V���r �N������f�j��֯�����T	Sq��i��ǧ�fF�Ty`h�;`�H�|'���=��l�f�+�$��I�ߚ�?�^*�`�@7����2<If����+k`���p/�,�ۼJ,m����,��B2$��0\������߸�>1��ET��x���u�Ym����>���||�~:Q`��SJ��:��*�f��8�Б�|7z8RH�S{&l`����ը��JA>-ub[��4�#�R����6W����e/�hX�F�3�ݱ�}�@3	4��ڦ����E�+�D!��IC���Ӝ-�Y�g(�+t���a(�n䆺3��y�I��n局�(�=mМ���Y��I`R2:2��qHqqn�t��p�U�^�k5_�Swi���8�����םc�c� ��B�p0�s���l�����������P&��`������}�ܪ���-@2�+KiQsv���}���"����liy�6��Ę�>.��~��<u��5s��T��*yE��н�������s<����(����>���Z�A*��`9u���LQ�wX8� ����8ܻ���6�su�χ�C;�/�y?���i���T7D��!���gl� �\/� ��%���'���ž�e���w
6Pm]}\�����R�P�V��ޙ���f�����big 57 V�j�w�W*��v\fVşG#q׭n�I,�`k��]���w��������>�n���K���OP���,�r,�w���$��:�)�'|Q}�6��kcx4(F%l�v���<&ƭ�x��E<�`ց�9P��t�o��,�1���5�؂�⧎]*�`q��45Dr�o)j�|�HO��±=��Ż�۬U�������/������� ���&Ȳ�@̆��$��^�dS�a������1�M��F���&���Ѓ�%�g����g��_�a$i�Yy[�Yw�����kiz��J��/��/����!�h[���P�~�n�4�ca]=���kT,��A����S�JS=i��^����a�6���y1<P��գk6�=�n嘾�O�c��Y��1mz*|vy��X�����S��w��q��s��hWg��}�&�N��I�l�b�,�m�`ѭ� ���kL�8�B�E5�83u@-q��R;�CWJj;`�Fl���F�e4ZI[�m�6|Q7�d�wݖ�+`e�l W�Z.1*cy`d~��35<�\]Xa�����t�t�W>*�H�W���
� ��嶌J�����S�<Գ���h�WH��Y}�yR��w��.(X?߻<����� b�Ev]R|<1�y6�TUI�W������:M#^-�GH������ٽ3�1��n��.���h��,�2����;�uɥl����R�>��v����X��+����ccP��eZc��F�����$3Fy���S�~���^�i ��A%N�Yi�lX�����/�J��LR�AI
��S�-�Q����y~ j�bBtr{G����f_)�����w'S>ֱL�����2�g��=6(�Y��t�+��E�Ygq[=�69�� ���<��Μ�=���q�r���xPտ�y��@�C����ѦVx�!�}��eKi��(A ���A�bT�4�q�U1��d�r���-�K����}d�\fz=�'�K��`F\"Q��Y�{��i<F�S���`0�x�� �V��\��	3�8�����G�_L�og��R�A��fU��/:��|C�X��;����+��g�|~����|D���ҩ���>�<�(uv� S\9p��Z��T�[q�Vx럄M[�m�� }�_���q�.e�䄣7�"��擘�:4cʬ�Ⱦ�=[M*��	��\��� <�[�8�d�+����yh��F�d�PԘv�=��]s~��@?�߹ �5�%z����ùd	 �믕�p������:�]l�.R�p}�(
�j��.Զ��W��鬻��K���j�0�8�eY<�3�!>�ﲲ�b�i��7 ��F�\;�/28�}�ى.�}8&�m8��C�����'V�]ǆ� ��[�+�����{܆���y������5 ���ݝ��z�.��w��R[�!�r�otc����p���@��:���J���S�_g�L@���=�?�/O��p0�e�"9r��Ψ�/�>B��8�%i��/_�@�ئ�Lq�Zҽ	��,�Jr�zO�� ��F�<�{��Lee��ރ�k�tӱ���O��>+�ɒP���6t�m�^6?�����A��ꁁ�����]rS�,7����$�,aD~�;�΃�M�Ck��Ű��k� ՘�h.'����VM�ʠ�zN	�V ��c(�QI�dK���I -Ѳ�� �ky���Do���^֟慨��v�&h~�yn|��� E�J�[z=h.k_��"?�c��kz�´�}M'W )�ں��U �����q��� cSto�_�]��� )������6����a2�(�{�\CF�e�Ӽ���GI��T��<Qf��[� �@e���G�D��o])�e�N�� &��8'7��[�3ܣ��Q��1�E'���n��&ؖ���o���ư��#���Р���6������8��n}����{���x&������V�W��P�������5�>=	ew%��9 3�9�X�O�8�-8p�(�T~3�	Z�v��wI�L� ���Ћz��=}�s�����休�n]��\c����]������Dt.*���(��yq?T_X�l�o���X{���	�s�P��ڒ���XVX�����;��r+��S�
�-��?�u���*�0n�qӎ�6�8���h͒7��`���W�6�}��X��N�6q�w�W��x~��իǎĤ��ş�Y'�@Po$�Tn�hT�\��e9�ֿ��Z9������W�=�T �ʺ`�7c��gV�:��ZW@q>����ά��ߙi�e���T��~�[%�m`|W+l�%��h�=o�t?��7 ��2��_���݁>�T�p7Β2�R�!^{�ۨ����^x �.��蛼Q��cq�����׃�{g�܍W=,��4d�����>�㻡_�����cp�yky��b�#N#
�nj:h4�3����"�ͬ�d���)}p1Z��?��4�����t���#D-߭E؄��1�Y'k��9�z��ze�x���Mn�w���΁�c`>c��e�,�˘�4�ߑ��2
�������n�\�%fhC�o\LK��96n��X��ne/\�YKW^��S�(�y���o����kW�I:6n���ȼ�4Ie�"B�i��o�ݯ�$[Pǘǣ���ÌR�)��Z�'����,±�[m�}�������Io��ߥ� ��*{���a ��Sߡ�[%�r�[�4(�5_;p�c�禜�G'6��K�Fπ�6���=r8@�3����z�ܧ������R(�p��o]o-YgO�d֧\�}��^�)v���X����2���Ѧ(�&��8Q������ƂC����~�d'���)��B_���Ѻ=�%T�J��;��]��_K_=�4З��Q��g�=�����e�!U]8w����.:$�1j�L5�#��ιN�V}g�`T� 5��`T���o�*ق�Z8?��2E�W�VcM6��PM<֋��i	l y�P�[�
�wN)�!�C�����|~q#!����!S��|��n��ǡ�����[��R�D�N'A�-�K�Y��t��M��%`-�ɟW�r�����'����j2�V����ʦ[~���rI\�����6��W���}p�2��}��/*6wZ�����%[�o��nZ\H���"���R��m*�p�l��ˍ�޺����,9��'�R�Dr�԰�g]�F����؁��5Fq�!i6���i`}�t,�z��ì�m��\�%��jL(��1�:�cI���z@}V]8�3L���#���هzܨ����
x,�B	����Qs�-,+���`e{�鿩K�%��[Oe>�$+�{���Jᜡ�Y�]G\����׈fƆ��- �u�lQJ�w�`*�.w(��r���n���D���l�����j8�'g�΂���v�*�2��~7r`d7&������h�o7��V�m���@'��X,���Z��mj[�k J%�9	X��D
w����ʕW&�y���o�";�gÚ����w��X/&�߻�
��º�@u��8-���ه�����p9�]n����	�vŷ�7z��Jo�7��a�(P$�RV�6~�}}�oIE0ia��Vb�������v9������c�ނ��(�̠�ߢhq�e�z��o��ZaL��o��9����<h��*0�r	��p?췣6�>_��T��|N��Ƨ�*�ߠ<,�~w�H(�t��Y]��
�ӿ���~���^�^U����,�3[�E��A�$�/' �x�o��(�����\�PS$O��@���鋅���^����^�<3�:�k�(B�ڱ�!
���������Q4�RZ3��������o��v�Ks�NZ%pB����z������7����@�9�+T��6/y3Z�Ae� UϺ8x��p�r?T ��{m�
@�
��=�Et%�%��u�s4�i�D��k��	dw������w[�ÿ�Fy�c�pG~#���H�^�A ���u��R�dw���m�DV��Ce�|}�!�ѩ�S�fP%	Cݑ7������F��̡�xf�6�3�R,�q��d��K�'����D�wQ�Bs��`����N~g��\����.F���~��f4dA��{f����d��b�U��8�����E�(
Ĝ����{��L���	�q}b�8�g� *�'fKS7@9d�g_����>�6'� xw����o��@�I0lX�-�'��=o���쩌g\8�%/�ݱK��k��:/�/u������s�7�,�v���1�_�"��z��#"{����M��t���H毚3�-�������)�D�<-}בE�Z�T�F@��<#�L>e��N��b>_Æ*>���rt�b ��P���jTc��վ%���: i�
�	���V���}�Oe`W�5�V���ڏl�:;�[���p�\�c�I��8�s��ˁ�ߨ�5�M/\h�O,�r��9���7�WY	>[��?�}o3���4�jn�t�;�)'DnQW���Q�s�5a�CF`|�z�$�"��~�z~&mS������c��������^@�J��΂j�|MxZb ,�&�oGө5^꬀�r<��~.�ӳ��z,-�M
o���6���>P�Ľ��D�^)4��{��X�Xg���c���{�N �m@(��b����/�ז� Բ���n
0�[sh\^I�'@=A���b�N!�$�����?55\1{=�O z��%��e�)��f�*"1����z���G�~�Y~LZ�<�ew�e���߬t	&I�:�=k+��h�����=WF�)�Qe��t��O/��so"p��j��6�L"�yw+�8Hh��߯pJݟX$��j���f	,~Ǆ���ܨ���Зφ���[%��14ꪁ�fe�ʀ�l�ŎMS�s�@5��F*)R�;:��I�l���j�U����l���ն�<Ի�Ȣ)V���-ِ�4�u�P�O)��tK��n�!m�S	*v�3����3���y���GJ)׿G-���2����P#ɇ��*�nN�آL	7,��R����Z'�ָ^=�Bqխ1 ��ԇj�SZ�?Y�16�IBL�@�&���lTU|ہ��N��CvR1��Ӈ�,z�{3������a/u�Ջy#��Ξ�L����{�
��ܕΩ��)اӵ�3uF�.���2�v�����������`*��ߨ�u��l��-��l �`;��o�l�绥���T��{��f�ԙ�BM4I��2��b��%66�����%Q�
Ñ+܋��׽�b@�/�lUe�G���{ey��^�C�A�/��yت���]_�x�+�[>�_�F���xf2�ϴ#�1�]�5eE��d�RJ�5�P��o�q�N}�	pW�$�B����L7���c�'��-�>�r��>�<��_�q����\!������t�ب�),�Gjn��tG[�5Q_q�*��F�~Q~^O��u< �+��֊����O�n���jj��U C�Ѐ�n8�-��Fq|@T�':F�������Qt��K��f��>7���%A`�n�=��<���:��x�Zj�����d	���{��˰�j]�<�R���<P��	F��}.ZW��Юu]01�eJt~�aճ]���Wv(�p.� TI}M�^/
p/�~���v�A���5�Y�u�W���u�)@9�Up��>d0e�U���X���/sC}��P��<���WZ5K^��s7�0O�r�XLL��x��Ub|^�+�?�����\u
&1��w�_%ӊ�//a�wW[�kUO�סH�����F�1a`����|�X4�=iAO�^�Q����Yr-�|Ր�fN��3בv`3�`�`}&�1��r<�9 ��P��[��m��g?�p|Б#J�|�:���N�Ux{Q(�(��u��u�ۋ�~͝Љ��=�&e�#�#��{PM�V�	�8�7��HTd`�4���sp�
�nl[��`������2t3;͏��:����8)�)Y7�Z��O��t��w���B}Dh�ߑ��u��ӕ��'/2��6��`��1��w���fO��;���������������L��:�ћ��V�5�ۃ����:t��$��(���H�Z���F����UEP"¿�j�m[�-�pϲM��X��X%�4hh�����v8��{pT�GO��\�`67����z��y�u7��C�̰�ϫ����9����ifxd�@~�?��G������g��h�s;�bn���W��	�`�<��9�z��
��i/�+�Ղ$$�Q'�q��V����
���`5���G��3��@��
^Z�f��b���N1�LS3T	��"J��-J��(�����qzf�7� ��ʹ��?����g��3��j�9٠
�ᚆ�/���U�X;aU�3��b��ts�|��g�>������V�%����ӂ�#��^ۭeu�y���j�qq*1���祡�.�N��W�b����v{fKs����z��P���o�>��|����"���s��~�Q�����h�f"ӱrǏ&�5"B�������ig��N��[���'џw���i�T쒢z�"��dw֣߳<c�t)E;����U, 5Kr��`�-^�[��?��i�
��_Ӥ��D�+[]��Ka6�i�=�wc���7�n�9���]%���=L{ ����Ҫ.�o���}q����
i@�e&��Fã��}��D�S��o����"����Ӣ�e<b�J�L=�����~~���r�N�16R���XT�Gb?�H����zx��m�났o%�;ϭ�*<���Y���c�S��3vц�A���n�� u����Yw�N"Z�sa{����P� �8�� ���6HKl��,��3�Q$����y�)������I� �MS �n�d��w[���*��Սt��u�0l����s�>���WL?�`Դ�ft9�|2�Z]d�d�ͻ��`�h��oZ�!h�JoÑ�]!JK�=�F�:��ꟾ�7��o3�
M��-å��{��2�4:�S��Uۋ|��@{x�]bI^/�W-KZp�@�؅��P�;��� m��|�-��#s@JF���L�dAW��w[����1ԁ_wl5��udB�K��B��C�v3٨��O��%L�(!��T�����m'���$+�B.��-�u*~]]��C�D�Xd˾� y=�F-�?����tC3*;��&Mx�dfg� ��pʳ��M�� v� �%��*�Jk]��u �f`ZOma���ӫ�K��ľ��kd��u��ޡ���0�u�.~ﮯ�z+�	�s�¤k�����3L��i��7�ˠ��&x/���q��l]���Ii���v��Kg���P{�=��!�]-���r�tC��h�5'j�j���7����K7Dd%&Ͷ���y��ƚ<����f/e�ǧ��<0����Id(���������t����Y�<j���_ ��<�PwU���n
U�U^Uז G�[�BΉ}1"t[�������QҔK���μY������ ���?Ix�x�=?��v�>���~m�_Q��*����Mn���%V��o��A���Od0����;���%ݥG�UkV;g3fD�ڡN�7�xZ��q�p,�)�����$)�s������J.3,O�1�څ��i�����o�\B��$��u��$ak�<��J��j'�`��� ���ȸ3"y��+��02��B��T׉�W�J�	L�!܎�2�@e�Y�ud��%=�I=Q[��75�Y�&؎�ǲ� ���K��2�b�� t�p��ʒ��j-� Ҥ�����^π�����|�+���*3{�1���m36��q�����P��������xX�~���*����gHo�z�m��B��	��G���D��6���C�������%�.۵��������x_�5�|���� ���9����*?GN5�vV!����Kj^t�g����D1I�z39<��'��/����v�ݣ������o��E�_L'J�Xl;*��Rf�^��/V��*�)n�c��	$1Q0i�>��'��cM���G�p��2���sh��:���Y�\�GK󎟹Xϝ�
�P;����Mq�� ���Ys\�ȯ#Oʈwsv�t��F&����"=Q�P����6j?QǴ�^ǭ�x��hA%���lil�z*֮��F�m�XZ��3���[��ז�2T��V�9�g�d/iF4�[�Tk[R��Y� 5?"���vA����ύ���Ϙp�� ��:Vt4f%�`Ө�� 6T�`N���.,A�՟3`�OSu0���	|m6� �Q���[\�R�:⃱�J��N,�E<k���j���q��
 ��O�U���`O�PѦl��������u�Y�k`�9b~|�$��G$����=�j�i߹n��^GT;�~,լ���3|�4���:,�Н۽O_�>������^X8���5�0ϱ)ht"УN��$0��<�<L��a�vG�<��i� �<i&��q���3��6�9�R�O.uZD��ϣ�H��]�HE5BKz��0�U���M�5�j@o������ju��^��d�����s�䅀lҵtj�̢7��$*�^k[p�Q�;	@�hZU�3�OF��Xg�O.ԏ��9~u��Sl��>�e�t�V�������.�b�������YP���w�j��� ܮ�m���4�p�
e�+���+[�Û��-���FW�<4k�X5�F���b�Xn)ПV?nج�a��{U��7�AHA����~�n��K_s0C�Dx,>OK:�(��a
J�Y �u�):������:J߲
���欄�y���a;��]��8��NV�U�g�^��bɦA\s"��}�b�Q����,-/C(��y!Ȋ?g��I5 ��O3�OE�n�BWȳ����@;Xb n�#���ق�rYR6�P��X����#;���n�
�p�H�uR_��1�6|�����ڕ�|�bl��K��K�3�>:�MR�v�@��`\ʙ��h�IZ��c~���X��&n�K��g,4���?vbTt�J�˽��3����x����hi�"��1����":�d�&�M
f�M���^q)�-�����^�<��F��:3!}���x=�30�,���B1���5��H����H��������*p ,E#Ȕ�S������(N�[�Θ[	�e>y��:Z�Y}l��S�`q��C�Y[,�k7�h%<���J*CR:;���6 �Jǚ�O�Xs_m�B���}���T[0�0LƝ�3}�E���]r�E�;��,�`�w)�Np���[�f���*f�j�;1���p$^��.�7�ҥ���~F����"�X�ॻYNPC�dlJ�B������-���߻�����]��ի�ATfs��u$����G&0�h�0�	���hI�j�v�������5h+������\���s�ݖP��kP���8��J�
z���T��f�K6\����}�1H8(o�K~�G��0t�����e,s]��w�[�k�̺��a��u���u��?M�]ө%�ȴ8�}���Oq�\���A��2F��1���K���c���>�N�>:�wX*�����_t84������¿D@��F�/N�F�4́���㖺�tQ��<�~7�Ȯ�`�HKJsbz(O]k��Ƅkq�d��J⽶T@����t:�B�5$@)�n5����[�sw�~�VH	�Ԏ{�Z��y¢�"���-�ܿ/0pŽԓC����Y�M|�S�����0i�7�#�}}�9���C�u�=e�bYdG�}��X��c�Z��c�fĚ��ñ�vY���}F�x���^�G��ӵ�9�-[\E-H ���J_�\�g�J,e�<#�;iC�Nfi�:�lR֭^�u��nr� "V/��T|�.�����:��Y��zݥc�W7���(�� �t~g�$,�}��z6Gμ��^i�wLɥ���I-�X�O�=M�=�� ��$Jͳը�nr�eۍ��6'�6���o�&��}�gW[%
V����A�����]~�U%7��q@�5��[��s?����1��u�n��|O��󌠊*�q&��B���==�Q��xoh�����㧗�]ESl��i�����kʕ���/�������R��o�n~� �����J�o�G�k�M���w�3p���U_�6匕BBe`*g��߿ ��g��"������tӧ�����(�"n����ޱ��$����������~����Ӊ|V2�:co��d��%��~��f߹���2TH��~���ݖ׳g�A�g�__�?��V�_��-�ώ���|�$�c�'��R�]'��������+������VuOK'���<��סn��.��޳!�*b�Ź���%�{�GI?�,_2��G��������{�v�^��%�2s�E�au��K/V>��K�񳗒���������xQ�	��O��9�}P{2�B�L{�b�.��><I�U��Sӹ����O\Z�X�|����Uz���| n��}M;���ձ\x����蟗Oԭ5�ry�|ß~��z�K�����Y��(�oy��L�-�w+����R~q+����. ��Ģ��qe?|�Y�������ӷ��|bmw}Ї�㱓��"������B�B��dں�+b���ָS�o����{t�<P�J��WO_�v�~�|���#�Vל�/�ț�+�%�'y�O��ϖ�ǅ�=I����+��}QG����K�'._��lbC��E9s��y�/3��,���~�|Y3}����+��V����?*���廜)�X��O���=߀�]��w�.�T���|���]>�|�w�.��|R����]��w����~�]�#Mi    IEND�B`�PK
     mdZ��S�  S�  /   images/e5551f5a-2fb7-4493-9527-57db21faeaae.png�PNG

   IHDR   d  �   ��'  0�iCCPICC Profile  x��||eE���Vx�*�g\�$�{�R�f�IvC�]�%�lv7��l��U����E�4��)"ME��   �4AiR��=sg��E?����d�y�3��)�s$���_�`Ψj�̝�h�{���{�U�J2:�T�͒/�,\���Ց�'�~��ǒz}���J��~֝1�p I�W,��K���- �~��g?G?K�0��g9z�J�'�7q<�ݭ�S�d`���>Iƭ�?�ha��������sA/=a`ͻ����;c�I�*$�̚�x��ch̹���A��$c�\�?<+I���g�\�FЭ�m�Ϥ�%�����2���L�Ve)cͩlf���:�����y��C�4MR2M��4�1�5�kʴ\����Ӕغxx�ඝ�{Y��"��t%,I��ݒ*��,iƫĿ,1h�HZ�Ix�:��&��;�%�6I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m[��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����,��qA��m�b��(I�x0I־<�m��d���䶶H<os
?>Y/�*����������\�\�ܖ<�<���|аJ���a׆}�5��pm�C��Z}T6jڨCF]6�ѕ�;���ţ�����1��yb�cg��b�?��qG�{`�F����J��x��V�b���X�UN���ʌU��j�w�ֲ�-��կZc�5�Zs�5���'k��k/[g�:����7�׽�+����p�m�y�6Zg��7�k�1�\���6���͏��~1��m��~�u�J~��[l��V�m}�6�}y�/���EM��w��W{�+I�ͮc����r��[O7]v�v]_����w�񀝎���-�M����I��y��[���>���w���η�n�պ���K{��6a��ݯ�c�^S�q�7���侳�~c��N���L6����۸�����l��O����[,9���.?x�e�|w�CN>l��O=r���>z�1W�k�=z�~'�;�SZO}��#N��ߞ5����\r^������{~��ŏ_z��G^���Z��p�'�=u�/n��/�~�˭�ܾ�����;���{ο��yp���,�����ɦ�����y~ʋ�_������ޘ��No�w�����?���-�D�X���3�0
�]�ɇ�׍�`�a��='���W�4n�q7���Ru��W��r�*Ǯz�j��~��׼`��׾}����z����kn��F;l��&�7=u��o~����K_�дE˖Ӷ����m����^�ts�ǿ�B�f�o+�5�zzc��m�n�f�o���;v����>���']�v�ΏM~i�w�>v�M:d�nS�N=������~�w�i[M�e��{�����7��+�Zѷ��[�o�ϔ��s�<`�wf3��}/���9��}h޳��\���*7^Դx�%��ׁCK�t��g,��;7}��C�=���W9�z�8j���8z�1��=��?8�ǟw��?���kO���מrթ�/������'��s�g�z�~t��G�sȹ�w�����'����-��܋g^���/���h��+߿꣟���r�:�nv�6��׷��q��7��r�慿Zv�Q��x�Y�_t�տ��o����w>����z��w���������?���{���{��?�������?v��?|��?��§�yzڟ۟��/��m�����?���^�����m�+����߫�h~m�ק�1��ҷN��eo���s�~���><��?��֏�[1Ɲ��ɿvo�a�&������/��5�ͱ���t�����J�\���%��������k���kݼ�=�<���������������	�]���'��֗�M�p��-w�j��{o��ˇn{rӏ�^��+���gϱW���ߪA�7��5�[���o��rǖ��|��-�'�z��]��o'?������Z��b�W��N]�u�n�u���Ҵ1ӷ�}�{�y�^˿q�7��?}�����o�O6�6c�`�̡Y�g9tھ�w����>5����ko��-j[����t�qK�9誃o[��w���|�f��#ڎ�����;�裎9��s��q��	w����>鹓�?�S_]��io�����=�3�?�}x��|p��}t��?^q�xQr�'?}��]�Ko����O���+�ꨟ��S�>����~q�����ȍO���/_���z��nk��r�:���7[�6�s�ߵ��{���u���ܿ�s~?�����8��=鏧>���S�8�O��?=����L�ˮ���\�����~a������}������m�^������.~��7.y󊷮���8�����{o�k�k}8���Ώg|BH�#�Q�Zä�s>����G�ї�i�_{Ӹ�ƽ=�ܕ����ʯV~�ʕ���ڙ�����k^�ֵk߶���>����_��FS6^���Mo����/nո˗fN8|�s��q���~y���]�i�扵ݿ�o�,;���/W�[�=�Q���v�n?f�uv�b'�������:鲶_����o����&����;�N���[���ݳE�iӏ���=~��s{����ߒߞ�7k�C�O�犁�g<8��̧g�0�͡O�[mΦs���8�kA����p����r������J^{ل���~���C�v��q������Ǭ{���Z��<a��8���'|ʲS����ӎ��Q�}�1gsֱ?:���9����;��������p���s�~�����K{��.?��<��~v�Ϗ���kN����~�ˮ����n����~y�����<s��r�w������ѿwW��U�Y��U�w������s����`����������cW?~�����'�}j������g��������=��#^�ދǿt������W��ο?������k���[;����}�9����]��߿�?~��_�譏��ɇ+���,/n�$����]�b�No'�Ӯ<��wW�x���a��R���k�L�R�H`�k��$[�̱j�Ks����#u�l�)y`��������%�Z�Љs���־w�N}'���ڤ��������8-I�w/3������u]�N�������x�ۿ?���x�̞l�����񊜡�!�*n�Ff�����+x�O@����D���W���������M��Fo�����/�����o��*_��'���c��㎡�m�W��#g �N��޷S��a�! �~ ���C�B��9x�-��|K�_��	�v7����x��k>�b�|�x٘.;�LaaB���}�A�U�����߭+Aֱ4�m�'�lP���T�jK�$�����o��ȍ�7"����T>ukjA>����AYƀ[ǀ�	��ݴ��P7�N7W/z� ���!�)U���a��&��u~����X�~��,w�����\Ɠ˰i�
�>w%Mu2hQ�IԞ�m2�N�Q���c���\��ȌdD��q���C�&���Az���>$d����fh�Z�'���t|
�RY�,��b��O�!�/��Mg�5��d�!e�l4�W�1���,��6n������>��m>�b��;��bNV䝽�Z�V*��zZ�ۻz�vW[�g-�3���?gh���EC��U{��g.���^T�7s������2��}r����]g-\0<�?��������6���ӿ��ٿ��L5��I��d�:Ј�������v���T'��tu���X�i�2���oR{g_Oo[�$1��ή���m{m�sZGo{c���jc��}�Í�ޖ��m�}�Szz��u�M�6���=�h�:�U'a�s��v�o��Ο3�s���B3V����wϮ6��sw[�.��)S?�-=m}��o�X����jk��n�ȻuL�Ԧ`�X\_�NVm����̘�jmMp�XZ�R[˔��4V�L��l�h߫mR_�Ծ=��4�6����X��>�mj_Ǵ޾V0L�n�m�:��kjOO�Ď6�T�؆�����胈����Lo{*�K���Ϯ6��T�[���ՁP��U[q��gTZ4;H�Ty��l�W��ͨ�'���Se����͝8�����6eR�ܕ�{ں��A2˳>�4HqbGK��B;�G��6����o����l��Z�X٥��7��x��}_�Wml���tN�ڻ������]�z�v�ֆc�6N��m�{_8a��5u
��}��V�L���݇�����1�����'�����L��[�i���pJA�������u5ɾ=ܿ{��rB�{�=m�=�L�sT2�v����Z&4�#�dk�Sa%�Z�״jT-���U5�Së�ո0�����|��OV���g�"X�E�1+MZQUvSߏՌPR`M5��Q�)SVWtU���/c5�,SUY��pK�	&S!*&J��%3�GGX8��S��ظ��~R�D&9��(-m�*��J��t,�,u�gBXj��GF+�⺒�И�?v4�yVe�k�a�c��d#T��Q�Qe5w��"�i�0��2��T^�b���Yn���2)-��M���(;��1���"���L1[5�$�}d��������יѴ���(Q�T�1�����*V(3E��A�d��8F�4V�Ɍ�c��:�d��wj܎>K@����u^� �h���F,˔��g	�	�&B2�II)�
���DZF����f������D�љ�)��ĖZwdҰ����X��L�-�z6)T�Å[�)�Q��pH���� �ɌT�&d��Y-���:S#�z��!�&�f��c��3���VO` �rͱZ�o�Z�yjmN!�0jR�z�՘4�\b��6�*�ak�����$U�,�*+p��aF�jR��	N��\#�q� �V*���he���5�2)�r#`��=PY����	I�]O��X�m	��b�ؗ�}a	Ο�贄PX2�P9U#�ġk�R�
[�X6�hN;�#�feʉ�ڹcq�O>�s��#��I����N>'��N*h��,�B=��$�!�Ԓ|)�Nji��n�c&ͬ'���(�p�b�Y��*�5o�uDF��Wd��֑��d4#����� mWp�ďȝ
Rc��0h������ؘ�QW3�0PZ���P�
���{������V0v�c���P�GW�4��)X6l�,��.�9X��
�!�
�9�[G����9~��;l�(HѺ�f�S-S�e�)!x p�
6.!j�T����(��?����g�(�����"��U���6U�TBR�
�#�g�k�C�GX�)q�>@9�(^{^G�PEi���p��A3�6��[=� �i�������a��hH��K"�:�+���疤
5�)Ed@%@�f�0�Ԃ��@�pĄ�2�+8#�j�FZF`|!Nj{���6�8Z���7VuA��BpO%N�W�)��J���F��* M(��JI��p\���mf��RZ�@�H�X�V+1�_G��Y/!��R2L�,ڈ
,E���u�$G��¬�z8;�pxX�2�����$M#,�(nY�$����q1����% �T��qdX���i�F(%�:��f@V
SK:@& {��ZJG�CiZB?&9��ٚD�68����#��B���Bt *��U-
K�YOh�m�f�U'U�ۑ�`�F�wrHaL�>��@dX*2-�aF
VO�&a���dH�Ҍt�֎��0Π��a�a�{p+`W�ϑX=��4�גpp��wX�EE���!&: u�"$\�%,��(]�5D�����ı S�c� ��)����W2�>��E$geK2��[��4�I��L�ɠD�ӒL��H~�4�L
���<p0L�_�+Dֈdڥ~��5���e{���*e����8t�đ�U4���u�b2M^�B9%��W-�=:��Q��:H�'���j*��b�����H�#+ ��'C2���U}GA����#�t�^
�uI���(B�(��(��g��z�-�'�X*2�|]8aC���
$\챾#�#<�Qsʩ0�Ó|3b��%eq UC�AHڎ�,EŔ�q�9��!�������{8VSVȉ'�����J���LX*/Q�(.8C�����<�BF�E�!GqQ���cF�f$�.Z芑%E��! ]�<���QM��|ᨒ�#� �t��
�����[�*d�xc=�g >H�E���H�tMZ,Ք�1�����Fy�&B�V1��Y��%�֨\J���nIu'�i=��u D�����Uj5:f%�@�`�P=red.��paι���� eU�:p���:��d��/�� `d��i�@x6+�XZA��?F$Y\80��2b��T���9e��UB�����P=^���c\*��8xPޒY!]� �V��Ǒ
��"�{��b��2:S��& �!�:�hH�(�� V�-q�EGAZ�H�sN
7I�V�Ҳ�S4��"'g�z
"�U�Ҭ�g\,"��J���L��|�
I�GV�Z?�MK�F�\�5�r���K|kT�T��|�����@��%�5�pF�.��\��\GU����\�l8;CU$��'\zH�=���EO���\Ru&���qFs�U���%�=����� ST=�j�EONY���*ydEU ��1Z�-�:~��6p�)%��r�YL�d���b��e������9a�Գ��{6v������M���'+�& 08���34�=y��D	Q��a�������K(=E��B\Flir���irƥ�lG֔�{"IǏ�'�Hwa��o�T%�&@oq��q��ʼ8_M��%3�ۃ�b��V�9��&S�l*+�AظO��lJ�3��L=��9mI��R�|"	@LU"CY)���be
0@CN�ƔH��
��²��b�p����"�p�1V�5�e*` -�s��6N�SF5錕=��� ߗRM2/��:`=\`��g$�p<B9-U�Ud�J��%^3�SQ��rߔjT��D�r�J�f�d�v-�Ne�ڒ1]�5�JPq�lؐl54����֔@ˢ'U2*i#OE?
��dX����k�U02.:OH�Q�N%�IoyiS�l��xIFu[x�n�>H\�����)*�k*�"�PO%��J�Iт�)�r5Fኍ�)�`ٜ�)z!*N�*�@aX)=yL鑘(�&QBS�Pw���fS������ğ��fya3��ss"��<y�����%'8Nk�uC@���� Jz�����?���\����l6��T�'�/����^II��i��lѓ�}�]	XC@N���e./����?9˔�G:Lm1���\A�	T>���y�U�'�,�����9HZB`,�r)I��5	5԰�
���5��ꎰ.W��*�ɍ��e)|�I��)0r I=%�������V�5�
�R9^I��=� uTCr��X0C���2Ms��}Cڢ��R�l�}�O�Ӕ���27�M����C��
[�oG����U�YQ�Ӑ��e�5�Q��<5ݏ �q�!���[f%�6��R�EO�$=p��D��IVҳ �
�vT� �ߑP)�[�K�m�	T�b�S�`gy����S�[��(�
hKF�`��=�Td��~����]ʧI����Jz��39��T_�G����2Y��>i�,/=��J�?�GOS�ocO*`[Jv32q����0�Q��I�  F�ψ9=n��JCB�4u,.Уz"C��j��V�a�L�F����B�\3�S�+�g�%��
�8��È��`�);��)^��O{��y�f��H�4^�%D�J;��pY��H�M�,�a ��E*3����jUYRU�kK�\:w��9���.U�����n``�0���m��}���7R 0x�D����C�C_�!e�BX�	˥{% R���(��2Oغ� �]�/��'�YHH�С��p?Tc��VL*���0����H?�!��j#�I�:�r?�8!������TN�tY�4ܕ�'�7-J�1�r{� �	��T==�AX��7�DQAf�f�,.�U�&��݁�4�dh`�SWa{�/�_����{����IlXn��ɪ��ϭ6/r�a��q{�6ς��6�̈��-��Y�y �K�U���dPt1D4�;`����DO�讑�HXmރ��5{�������?wh��>&��x|�������}F^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� WuQ���   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    T  �    p  ��    x       ASCII   Screenshot(/��  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>1392</exif:PixelYDimension>
         <exif:PixelXDimension>340</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
����  ǸIDATx���$Iv�<"2�ή���ٹvg�b��hF�J&��Lf�*�>���>���H`���ٝ{�ﮮ3��p��;�=�2��fz�SSY������{�7]�E���s4�O�7���A�h?8B�>^�HkY<
�w��G�_��}�� H8�:��ȓW�x�g8�9�>��ÓB��El҄ z��Y��;�[bϧ0gP�^A�hLQ�5Uv�\��nru�@_;����9��O~���]���w]O�ŜNNNh>�Q�u���3�Ni>�1��J�
B����x¿Gc��Q�?L��ф&���J��z�o0A����oi:;����� ��ތ'|Ѷ2����9::���}�p�&�ի�hē^U���d̄�CM�L���m��ݣ]�=ij��f�|#	�&Т[��Ǐ�	O��l΄��ʟ)!�u۵���*T�߅O�>�G�1�z�|�c�'�an��],��e�4��ss����6����b¼|����7M�,������ղ:`�xzx�Y�)s�t6e"t�!3!��/���%������d���q��mnn�(�Hk�3@|O��?�}ʢp��N�:{��{�0|(�E��F��bd����E��1����&ƂuH+Z��T��pV38�.�(�A?3~o�?��)_�����f�Ҍ��ڢ��ѽ���ÜRQ���oq
�Y�a�ȑꂕ���)�9�6v��1���ų�zs�0,��YO���	��n sY�u]	���P��������<T�ގ�p�Q�� +��9�<��?4V�)d�H��T|��mml��/��J�a��
��K�;;ۢ����D�=d�r��]�L\�6s����X_�|�����TP�u��o6A���Eʓ��+���=���+��W��KL������{�f<�@N8�By��'"�	rt|$bp�����Ç��`������}c�i�#�5�O5�*sk���+���.ݼz�a�X8F�ȩ��$�1yc2��fE}��u�tbӴ<�?�?��?�����;����p��o���GTc\Pӫ/�B/ݺM5�+v�����L�Rxܧ���!����A�<������(\���Zs`B��U��oP�E��P�v���VxN���9�_e΃�`� ��"�����7� �'*���Zt$�c1�g;9V���U�#���ǢpcB�|���l�l3��Q��~K���$�rU7`�*�1=!��`L�t�#�_�儰5���-r2;��!�z[����E�Jꩅ�� � ��*ӓ���X�#�m���>���d�t����9���3�y���ٔ-�y����.�>��	D����Gc�(�&����.�{�ŵH�1�<Χ�1}!���2q����	����>��cz�����^�I�s�y*�Ť�?FT_ܿG|��k�6K#�*7���A�G{e°��7�������?��7nJ�̑"�@��(�/�_����4���ǂP�P�q� U�������+$.�2.���M*c��K�m������������[w��?w�n��5�W.�X$E�;��&�q>_��ֶ�#�⏂���	�0�����0tq�ZM�X�O����
#>���|e�Ŷ}z�`�����L���v&����b��{ e�2aqs�ݽK���ّx��,6:�d||Mx�Ă����c���b�����,	PݼyK�w8gE�w��B�i��ϙ,&>�/�t~w\�f���x�3-d�Fu��K��N=�_��h�z/�(���#}~.l	(�$ܺ}����Т��9u<�LD q����G��FB�-$^a���FL�_~�^~�U68���rΌ��a_x�ga*�\9AVX�xO��U���e���?+	s|zBs�j�`һh��&�3:�XT�!�}��T���	��F���ߘ'n����Bxiu���l�!V�Xt�1(��R4O.�jT' 4cV�x�k/�4L����(�$ $4l�P��Q�͈.s�����tFǰV�9����R������Hl���3/:ԏd�I���I4&F����[k�	��>�>1k>JЩN\))��#N����ʘ(�<[�a�reHb�r��ǡ3`sd\j��"�ܢ����(u&����:% ¡��b٘ �r�-��Gq�yP)7�o�: ���KB��r���0
��Y�&bq-�K ��Sх�M�:��z�4����ct���ϫ��\	��U�y4sI[B�/K�ѐ��a�C�R W`�c%���5�AH#yv�9���f?������U2įdfm��wo"� �O��y��#-h{kK��V�DW��$^b�-���r[�9�7�}�'�)x�[x=
<��{t�c5AxP��N�Nh�ga�6xh�(P��d*C�Zro�� �lY�KsX%�T]��X��\���d�0e�������'�W�������M����K����������� �P&MƄ���𺣖&�?�;}q��N�@~��rP�жQ�%'�C�\�4:ɑ�� �d�yR�Lt�]b��-��bF"�@�d0�c�����|��xT�J����O�Ν�d�5��J<���)L����f�h�b�Kg�>�V�!z�����&B��#�:�	�_i�!XS�k��R+r�i���>��666��W_�����CU���H��JuKWB�>����$����H�Iq��-h�sg�
==xJ�!M�J���1_��	�D����E)p�尞HC𢩪�c�恣Ưf�x��ұ�Oy�AD\��K��4���.s?�%uE��J����9����"��{��	�Z��,u��R6 �cU�h���,�3�&�[�1�pQQ��Z����x7X�x���Ǵ����z ��8!��s��+Yf�x
��&�1`��HT�W*f]��nȗ)��"��.�F�WI�{n�b��I�n��٢s='�8Ӊ.�ϕ+WD�!J_�qCN��R�$O��C���1�nHDȋE�Y�p��,�7!2���I�'�2�7X41�r�*qA�p����.��p�FY醫	���zC8�$/��SLi >1���rY^`��ݢ'�.�h@M_'B2�B��@Q�Ϩ5�F�Vɹ�EsIYe�j�e8�9d���ɣ��@!����W�Ĳ�JX��U��r�ؗי*C8��A5 UAg�$nY��&MP2TWf�+�9�y%b��Գ\���,#�L5��	������Od��� �k��'(d�g]~�4y&��7 �{�zU�A}Sn����>m�h�ِ����>�������}��(���M���qO�&HWD�(�=>9�����ޡ�W�"�ϲr��֓1cr�����"��t����`+Ox������ӢKˉ�AFP�FIN���|�k�Q���C]�ɟ�JBE��P�3���B�]6<���}65� Āa��c[O�g�*9���*����pD^��y]%���j��?���|�,)�����4�����mߓ$��d7�5r���q��Q��8�)Q�'��ұV�Sz�J�y�����zkkC�+=L�ɜ-d��a�lln�R=|�T��Z�z}��� �����"������ə�B���������r6޵|.�#�m��+vʥ�9�q-�
��'cqa��y�"�F�M��G�.I�5�������+���(�&����܋�wC*��C��CD�1���Vc����> -���2�߰�aԁ����~��)��H��K=����� "������+1whq���l*��|�pz|D'����,��+爡.�b��\T��Y�2��0�uX-9�t�mmo)f��W &��p(������J0r ��&��X
�`ۻ;T�c�+�+�n"C[�][�#O�<���C���T~f(Cూ��PЃX�[��(��c|��U�.�[��ń1��
G�1��L����3�1y,���Z4��V;j-���ȃbՁ(X�""�Dd�9(9��ꫢ3�P(<�X�{{Wikg[&�\��K�0:;������}�tX�O��������c���`Ԟ0!��, |�T"f���ի���_�^ ;�7
M!�I��GV%�*�@�@{"�(s��s�ITȨַF�0yw���ϱ���#���Ipk.���)���xX�;L &f�t��^�f+�SWM�א���*���Z 5�����C���������O���;�����]��A��[	<b�=~�^�s�^z�e�q�,&����]�F�PW	��	|q1TƵ�(��~CƢn|�ɾpr�0��<��I��#�|�(���G̖;q��@<��۷�&?p�"��	�x���g���E�� �yҎ�<�O>��~�_�o~����L(���ߣ�B�)s;)p�����\��c;x��N��B����z����W�\a�>���+V��~�L���ļr������V7����7V6V#^?z��޽G�<���B��~�7�HP�E��M�����������d�H(����I��=�Zv�7p.������k��O����޽�Ro�_�����L�I<����t��=A�o�񦈹��{_��.���>f�vI?5�͢�⋲�J.'W'_ٹ�bʅ'���WT;&`@<����C���E<@q޸~�����M�{e��rU��i�_�<���ҟ|�1����-=dN��;�0���c����I'�B|E���8�U)	� "���O��#�޷^���wK��,��?~��P�h��Eses�~��~@?���D��g���'#)��ؘȂ����$���ʒ�s���	C�xˬH2���\��>sB���O>��>��S!��^�W^yE"f��)]i�D����ݱ8
�88B���@��/>O�Xo�����?U�2�OFX�%�&z@�/>����/���C	���#��1� �{�!f16��ڵkr= ���(O���/g�S0~\�	D��jĨ�},;V�X�����B��Պ�fu(A�	��?ؿ������w�cA�[:s��@.S�߃8�W`����ŗ^y���'�|"Hv�
��bbϘ����_����i~ʜ���=z��!�`p�A��b�����8���7�8�}�&^���p=��
��d��t��f�;��2o}ᠤ�C���:���ON�ʂ+0��ypX�x�	�	i{��6�`�#�T�� �b=p�u̽�w5w��	t�)O�w��]Y���|�+qc�ĸ�G[&���n)q~F�/�����E'�o\��vö��77oܐ �'�X����a���Ct!�;`���r���|��y,���( (������G].[�"Ab�� �@�۱�Yy�ޯ~ŨE{��^9a�|��_����tN��) Lu��WĜ�k(k������$�u�5z�����?W�΍k9o�_�<yN�t)���>��^�U�!+���pL����5o i��a^h�x��[�fx*��_bpp����<~��������S����x.�}׺���I]��Ѡ���H)�ho��!�0�;lW	F��z��u��}��Ǻ�q���Ao޾�,r�o���^~���������WR�4�x�2��\c������b,<�n����g,j`�� <@t����PY��}4���`��8�~[3�>�ЗDY��C�ʋ���≸��L�'���3�dU�uֹI�}E�>�:��� �e�z? +qƱ<Ɗ�����ؚl���҂Wrz�e.&J�l��W����X�w�z�-����N��Sq��L��(}A����Z&
���@�<�ڬF�8��a[l���LL�L4,} z�w�b�O����ͯ-�q�<~�evF����I���}�a�O�ܲ1l��BN�{�{��������"��_���y" �o3���/~�D��av������f)�P���S0Y�*T��f�,AC�Ufb�n�ꄛ���N��k4�Y��u��)�)ԗpjP�Po���,,x~A,ɨ��]���>#)�^��\n�/_�#a�L�j����y��'���'S�Lq[�`QN�a�hl�`؈�-�M��^���$�.&m�>��3�Bh�d��=�}�����l��9jS�:Ei�(�>16xR�����LI3j�P1U-4A��O����Zý@D�ۛB$)�K�g��DJ��ڌvKی�m���_���o�N��(�����ՊT��4�^���8fq�ڌ>g�E����ӎ��=�ʈ����x���s�5��X��3J����Tf�XYA��ύE��6��g��m�G�V0�+<�G@5��Ome�S��H�L�t�ސ��ٞA�*�ߖ8~-�>V�c����
�ؒSVr�jI4@��M6���;�)�'�����n ����ߡ�_�5Wz��n�}j��>��b����X��O\���hEac|��;2�O�}�Iu|n��r���}��GP?7�(��,� {�}�Tϋ +�t��Cf6&�eR�=`t� �F�t1�x�gG�(2Zy�7İ���g_�O��oX�?�*��}�{�j�� !<$�yf��oj����3|o���~�0􅱩1��x�5[?Z��T��D' �q��%\����N���m� �X�����[�!{.	��Cؒ�A��9�)"	��3���W� �
ԅoAΦP*?�_��>����k,.����w��TU���$MX��1�rT)n(a�^�1 ���8$9�n�G���[Ҟ�n��6x���K�Ӆ�23�?�VX�Y��b��J% �B��Zy�R�~%�~e�H�I�,�^B���$�X8"	��0UjG�D���T�&1�-���&O�|!py����{t��)�?�������o�K������Y+U8��خx@�H�e��'�`g����؎�h��7b����CD�0W`��|,�ƒ2���0�nr�b����M^`*b�a�ci�)��n4g@����#X��W6����LV��#�����M?��OduI�a�ڪ���G�lmo�_a�y^υpG��� 2����}[�_���d�a�v[Z]�&
q}�����q�!�^�c�'�g!� 7���<�c�� C�J̠���'J��⅀ژ���b=~�̮^��P��A�=gS�.s������?���`����������>�7�z[2Fn�D�5�����槴�l�@�A8:�;��?�w�N�X��MQ�����˯�B/0�x~V)	4� r�a���w��\�3::=��-�ܞm��_I�B�@�XD��7�^�-�p.$�B}�Y ����W_�#6��M���M������r�:�'`���K�gFW����J�ӄՄ��3���������o�@���>���[f<����D�Jp�[̅/����v8"յ�[��L[��]���/��~������?	A���񓁊��Ap�/#D�7��D���L�;����`|���bh���H��6���Ap��Q�� y�s����=�^KJJK@��m'�����}���������C&�(XV�s�X3�j�E X�+	���߫� ��KUB��I�������������D��i���P����ċ�˟�\�B?<��6��D�A�b!�$�ϻ6�)����G��;[t���P.�����LH�GN�[�[v�P��J��	?R-
~��?��M�����|��D������s`}��w���Ġ!�g����7^g#�����<���{�Ͼ��d  ^ʅ��v��֑�� 0�/�տ�{���1��m�#*��oݠ�c�C�}����5�� ���g���2�T����w��o���gn���-�RX�M�$A�
���u��{V0�&UC��H���^`�o�)+��u��WX>���_�k7��ہ'�֋��ã{��­�����/
Zdz�n�y<-)�"�*a��������/�����^�Qz`���7/<���0T�����>}��\{����?��pߋ��l%���\�9�����q.A��ue�	b�z�k����A��w��bE��?�Gz�_��@��@�7�}9�2nؒ�[��������$���������B�eL���[U^���`��hr���,2��B���G����O�#{̡���gn��(]�- �>�HԸ�G�o�F?��w�����/��:R{��$�TȨzE���%ɼ�J	�ߐG7��mO�>�������?f��%��?���� D�泩X��$ �N���N���������N�r��$e5#):��e6.��Z����ٍ۷��-��_��x����?�1Қj�-�? @$�!!��<���">�dD	��sb�H��R�x�/x$��.�F.�:�+_���͉��|T��Rƃ���?�_����|�Մ6����6�Q���.b��5��M���=ԞG/G��c�y_H��b�be��ٛo�E���=����JB��|�$��g�\�1|��7��̥�� g�+��E�r/Җ9Mʏ��~?�CB
�g��J'eY@Q�s�޽k���86�����*�����s��ce"!0�߾���&@T�7��k������[�Z��\w�މ8+���tX��~�;�o�����a����Aa��G^~�eI��v�m��M�؍&�F�}�(���P� � �~I�8����T8�r_W�����N��ѽ��Lv
�[o����@F�SP�#��������#$��w�O��-��Eٵǲ��Q����2��(�f1�}�;���;.��#+D�k�m��]��">�RW wU³a��<������������ڝ�paY�	0�6��H�6t˶�N#�5�D���:�4�
�Ţ��i%k�o��B鲇����ؼ��>� ��r_CH��\���:��^Wh� �$Ҳ����[8��e�ेT�n�+n�Y�.�U�  Ψ���e��k�D��A%�	+��ioew�F7�2��+ԥts��X��H,���[�)��Wg`oL�E��U�,�֬�����;֢,���D��v�o�X����U���e�2��[ۢ�և.d�L�Ք{�`V��Y��u��Q��c&�-�'�锽sV�eo���)������w���YC~�}������E(䖀_� �j�k~�>������U�<��D�^�T4t�+�w�&�+����r&y�t+2����uq����<�%)�A�1!���?T%HO�ABZ�Q[�4-��(��EN��$}ˋY�`�_� �(Q{��]�#��z+[B�Zc���#{������±��*:��6]GA��C�I-��e��t��ظ���H%��V�lib�SŔZ{�g�S�~'��_]d�{���C���)W�i�25��I����J�%��D���1�3ܓC�V]��r����=Nj�䟅�8!�X+����o�X���R�DU,����9��{>b�&RF�h��^����dj����+��	鰕M5�I�����yw��
�	������W6�uA��;��r\�mց4\��G�*I[jP��ˢi�y+�H%����`[ �<������
4��řn�����C�Mn�`};i,+��o^ޣ<�a��s�w^(��W�Q�(��=)��瘣���P:QS^=�*u2�i�S�t��:�~Mz#��??��ׄh�b8A��N��1�χ��6���j���/3	��!t`�ڊR�2�o��Yk��ET$嚑S*Qv��)����<��M��,�x�����>2��t�`��E��G���2��ϋ�K��^+~)���W	���Y���YUt���A�[Ɋ��1ĳ��pE'�ťP��%����#o��� �OZ}��� g��}���_#�[�DRR8e�$���v���t��Q��Z}�u���@�\����*�9(�_�l7!��-���t��!�M�IG������ϼ�2��h�|?駸�����j3���y���[��s����� ���a&�*d�ǹ�.�!�?s�$�}<���]b�=.2ₔ��ʥ|��t��gM�B_�{���7�xn�2�[�MT������eb+_ױ>�J��D���ɸHg��]ĥW�ԗ���и~�N�e��n�++wώ����c9�0J~v�!�^���%���x��n����#[X�AC��]5���p��]�W)�"p����YA�@�f��{H$�G����|f���g*�����:<���Y��o�B�������}�sˢ/�)#������]8gb�۫�SH Cq�x�e�9��a�������q�\�M:���%�?+
�V��|B��
�LI��Y������tDg���g����6ID��s�c}к.Ëg.�^�����7�lQ?�Y�y��.ow,����N������.s�{��岾ş'���E��aq@���8����9Xɫ�]���_u��i)��Ķ���znyK���9%m�OKڢ��C���Zo�0s�?�m�R����#b�/VF��]t�r��O����.��c���Y\�x��z�@۸|~��>5��Ĳ:��]'�BJ�;#V��9s#�o�8'�zh�����2�xdL&�}��AO����l�h�K�Ń��зH��������Iٚ�qY}��<c��0Px�2˯д�d����i<�C�O�il��_�������-�pF^Vq�!E
�Ͼ}I�<Cd�U�:߁�ş���ϲH;.!�pH�OHu�ϊI����r6ܸ�м�8tT.�,R(>S2��3[���Y�c&���I����yw,\$�~$$�k����-]9hh���J�%��@fյJ�}P ��]�r2\N��l�f�i1�"-W+�jh{�;�3Uw��V~���2i�>K!Lq�'��d/��6͉�-��Uֵ9�6��2x�ٽNV�y0��zXz�4_�����6��5��(<�̶Jƥ���O7J�i��K6��b��Q#��R-�ͭ���	��sj����{ai6��q�w�@�[EV	9:r��4{����r����䇳r��IRr��3b1!����r9[��9}f�<���w�v�B�/��S����I�&�A~g�b�s|�����+����$^���~��a��̔�Pv/+�s��dm�ѐ��I#8���B�9Y�t�Ϝ��}ͳ���&p��y�i���RiA�0��w9��vw-y�zo��OX�5�gՀ �:'�n�Թ�*�B���s��,7F��)WG	��l�T��UH;�{���i;��_�+D���	O/�ՋY�}�2�k�,�ӂnE+��]$<r��ד�{k�-z�����(�����{^�T�38��� ��.���0P��Q�_ł�tD-�������l�߾����[��ER�wu�D�uι_������m4��x�AdX��TPm�R3[�,Ψ�.)��[+։^�;L0F%�t0���pM��}K� b����ґ��W*����h�^��votc���UQ�鏎�ڪ����LD�g�����&�;q�n�޶��y����j���t��m�f�1��]���'�r?D�C~������E��w��mp�ŷ��M�����K�RJ�BK4��?P҅n�*"�vC�G�� �W碆���{��"ֹk�t����Si�!��G�%�t����(S�h��ߨ�G�H��*�jk��;��@����I��믿&פX	�5�Π����F���r��zJ���r�1�����1m^�J�3����dF���-OS;x�L՛�o��u?©m�����.�x�)�����^[P��ڡ=��/D�m�(wB�!��:��*�zhT�"�\?>y"��\�����JŽ�����Ûo�\I��q���wy]=��{�Ԋp�Ź��۷^���Ѥ��TfK�}#+���CQ�~��v��؞2q>��s���|��u��sE���A���}�x|@-+��1��������՛W�f��������������ͥR�6C����X�&Z��d���Fړߌ7ebd�;^/�������t��N,Pa��.��2+6����v�e��iׅ��ފ�BE8�1���������4���%��&�\&}ww�9q��=x�s�\TO}z��$�n�o�AT�v<�tr�m�H�-Ni�=�'��������H8�ڵ��V+�yU]��l�C���K/�@���ZQqh.;�$^:Cs�mG������>�������.�C��r�c�(1m|�V�A�tM��j�w4�������}Aw�=b�tf�/���]�3���k,�1�<�Fs��	�lT�-�t�s)�D6C���vI̝�+Bu�(���tK�H�GҎ�weo�&hj߷��Cad9!�U�*��^�"��K����H'��,��'{�O����G���B76�j���>��c�W���+���b*�. \�s�QE�vJ��Sِ�ʮ6���-_�X��ye��G'�窝3G��L�?x�7�,b4t���m�W�	�r�b���ū'��+ t��u�2nA�ob,��Ë�V{�o0����iGF�o�cL"��e���h�t�Џ�X<��O����H�.��[&�tz��
�nD���=�-�����]e����O�0r9��т��m�(A��cFs&��
�;�mn�HK��m���;�U33���e^�^DS���pG��r妉676d�����#�gW?Q(��N��\c������G�0�?��um ��4��\�/4
��-��C8Yy�!�g2���f�|�Mǰ�W�T�l��AQ(�@	5Ccl�-�sZ���O�y�u�X;�������AQ\�$�lpZ���ъqJ��J�-E����������r<�h <�v6����~���߻+���YFj7�#p?m�6����T�a�9�HB���\}�U����}�!�0vw��b������#�˖�dd#i�i�ؿ��{z���o�(_�ER�i�*�A)���H��ޖ*�Ѿ��Н�f�9�>l𷷞\U=O4�����W����
q�b��-;)��b�޽����]���x�m3&��l؈��bH{�/F��������EH�����)� ��uM�ܿ+��mb A�,Ʋ��DV�CA�6�]kH��DU�E��I�֖��c�=�;�|����G�����d�Ȉ�&�旓]������p}$wP��j�6�Ld%������j��ڶ��R���G��g���6���0�$�%��h�{����+$��P��F3�q:(7 ��|g2ސ��z�_(! E�.���o�9p���g:����x��dSǊ=�f�m�<�}��v�Z�
�k��V{s��H���Zl����!�H`g&�G���<����{���V=2�/m�:�B�Mnc5a�8����PWI�b"*k��M��j��%��@�e���d�����CF4/'U�c��6Y�C7���=*���K%������H_��;!o#6Gٍ�V$�[��6��*�˶N�/�)�����)���ĕ�m������d��Jj�4�v��d���,O�
�dW�Z�!�C��d8�����["u�>Pp��b�g`��Đ��W�ҫ�T�t�W
�^�p������Ψnd��@Owx�]�q�J�ʔ�"M�d��6�#O< ZQ�cSv�Q�)Ȁ�1 ���@p�p��eߘ�H��,Fl{���k%z� �>.��/���z�-le6��1��C;�IY0���T���8V:��5���a ������'�%�Om����-���5?����)b�U�X&i�WOu5�g�[�`��T�?�p8��L�@g%
�jl�:pވ�ȸ�N��Q�.E]�a���<�P\�T< .�����6�nc�'EF��3yyp����H	��0�vc��yb���U��9*�]���f[�J��^�L�m�����	��o�W��c{�Tf��uѫ��O��`a�o:��e ���mX?��K�V�P�>��	Z���̀y7O�Q�х,u5�h�8��?�˓�ӭ^=7��w�@_�c��7�m�v=::�A�t�5�5V#<��v�t)�"!��ģ�Z<�����8;��TBi����;����Qg�I�I���ݷQW��4���gp�x��y¥2��ql��L�y�܉�(˛�$���9���*�X�ط	�zg{��-�aU9�p�9�͍�1j�'GW�K�lK:�O�_�Ŧ#���2$�X3do5��b� �l.����o�����[�l��ZDܢ��c�U��֎n�Luwk��u�8�H��	b>��2��P�cV��҃�+���ϱlT�6o�`%��/�N��4���.V��3�011c햻ay	E�i�5ڇ�'2_��h��_��A'%����=�e�2<m�20)ň �X�Q��b���=b]�1駧3�y����������'],��.�C4�+�>7�Px��Q�¼��K�HvS���b�kyR�*�>�1-eEF���܃\%@p����R��;��͐w-P�Ge�C�:&��̐�;�W���-��!:������l�K�k���Z�ksc[�ۗ����GʢjT�b���E2;w�@G^��&�Y��ãC�zz�l-���>#jG���8��
x�����nI_��1�0�X��Q;�m�>�Ő�$�egJ߼�řl�'�F���]���wc�7u����ͮ�%���%._�LJ��e�!8�����A���:���vK��)��r�6Gb#rK�(63��bt�^Uw�d�l^;gzl���e�¥bPAenV��_f�hK�WKO�pg��ed�Y^0X��Ƃ�2��8n	�a*��AʀØpз��(�i���+�
��'#�7/�lt]٣��m�pVA�7����5PR=�+lG�d)[�5�J��5w�M�(��vz�������������DJv/��%�=7��ut%�m&����mf��3���ʍn��[��g$��GPt>e�*��Q������6$6��V��������U$; `��� .�m]7'OZSn���t�?�CI�59�M��f��G�7Ţrq�{B��G,�W��z�����(�m�1nl�h���I�%��y�ߛ[�	ek�Ⱥ�"�Cv+�]��沽����wY��H
��$1�?�r���U1	�d���w��l��gœ��0����!���R��H��7&�����EZ7f��h "UHa74aTV]k�!�C�g	��*)1�l�Ӳ��Ԇ˝ �ņ<�û<��ֽ���LYF��!�
�'^���?�`"�b_���?���h���,��H�()o��6�����P���S�b�g���{��+>�)�{	�e�*�mѠ��97`0dpW'\k�m��d�V��?i�� sҵ������
)C�?@�-L�~P�!#D.	���a�bro����`��7��i.{~�O㐑������]�8��y��5)�-|�H�q���½��鋭���˹�y���s�Z��y�Z�Fq�3�&�[E��^~��u��G@uZ0~�O�[������_�k@���:�8��Y��±�_��ڶM�����{��0��X�u�R��'l�^�h�;���х����ҵ�=�o���__����X�PY1o�g�E+��q���.�ʀ�3-B;֦�����S���9�==��|nѴ�"1�EN�7	���cik�|Aq�dQUܐ�@D���y�&å�S���=+#�Z��HQG�B$�#��u:Vf.�L�Kqu�+����,�RD�	.�z�J]�+��l@s�=�&�$fP����]�2ǭ$B�99���;[O.W�1��bR�]�C����S�X�)�Qz/���w0nA�p>_������m�Ήc��IVu}�0o}-�PO��٥�e}��e�L�x�l��ގ�#.����I���2�#Q�M����9K�\`�5vX+�o��(ɘ#�#�f�o��g��]�i;��q�\�(���^!}V�����4y�]$��*��s7+W���#f�!�!;2W�wu�NP��rJ�!�!���".��Qo��M���L��D�����
�V��tK�.�%BN�+z�%����� �W�]��f��ԙ����x��Zaz��:=@�Q�dx
N)����4��dD�pV&��Fhf��>��c�Eb��m/���y����2�H�*�g:xTM�̱s�'�ȍIu�6*�ڋ+	sֹh�v�*Z�MU)�b/���PCZ!]G9ju�JW�_�8��b���]��Pם�z��lW�m݀���Fѫ��#+�&.���9�����dz\�8@�N���%�G��"���e�EGT+�]��ι��`�8���p�u/w���XK�leD�� �C�-�lAH&�/�Ե�U�ΪnB	g���*̂�������=Y-{G�=31�� �-����`��9v؝D�E9K�Q�=@R�
8�h�m�%����)xY�x�������5��ؤA)�h�<X�l��\c�?=�&%)Y&�{���TI�L�9�+�Wk��r�ui�H��n|V�<�d2_8db��3��3�0aF�����
�+Q� ��H	���=��8=��b��G)���s������*|^Z����p@'3�3�NA��{-Y���L�/���9W�q8̴�ʘx&PFK�	�n{d����H�I?�9s�(�C��x��		�\Pda��c�w�\٤�{��4�(f���\�3S:}u��{���NTw������g_Թ�,]#v�Ɇ���=.O��
��K�P���m%Gy�Hyc�$R���!~nk��Z5�.n!���"�1��jP>�3g�au��&»7�ct#Y.qhݯZ]C�d�`3M�C�SU���V�]Ht��57����l��a�0�}"�K�^��g�Rﵴ �tA�Y���.)���!v�m�E�?`�/_K{ )%�Ī][��ZN���!A�7.�X��lp.�=�/Ti��}���6���k��آ�^a�_���m� ����jT�dH�|�D�W���}(�a�Bu
Q�����4��8����G�MV���>��=|���+�������Q*.x
�����]wf���c���EQ �K�՝MR���>HO]��I���c��Ƙ����nOQ���r#�5�[r���y��;�l2��m��=�4����
�S�A_Z�ꮷ&8��!Q��B@��I����\I^�Bj��8��J�AA��>Xs�HR��Q!��tf��F�C^�Z�Lw��IG9�By�h�Y̢���&���g��z	��1f'bL"�av����"7&�������ɹ̜U����
WAH~�!��[R��#���J�X5<S���|b�=F� Q�%��|�	qH+ñ�=_��eٖ)}Yrm�=O,�G��j>����|��R��N>�c+��Mr�d���ڹ>e��}����\����C삳�p���3�L��+O溭���ͥ�hϮ�<*�R�vȉ�n����Uf�{i��Y�.�{�J#P����.7�$��zI�S��a�+ev)��T �B߈�`��M�P	/
��2dNpc�Aa�����MϦ��aP�+Mg\_��:��U.�g�~.�BY8���'D[��(
.�ͺ5�JcyK��<]nq�b%���J��n��bN���@\��Rb]\��1'*�T�Ø��5�<�4���+4E!+�G���-��G�g�OxX������#�T�Z�țx��fa�z�����R�R"F)ˋ��Г�V�P��^&B��^�ԥ���jQ�����J���@��F�q����9O�K3^�H��>_�	㫎�M0M�yU*�����w6h��fS�*�$����%hw!eϋ6+DU�R�%���8�'e�t��	^���+{�H��K%w�˟!t���VL4��S�0x%���r7q�0�|��)?�"q�C��_� F
��XD��N����k>��fDG��$�2"b(� �N���6F3ea��fªc�_"L�g$C^�^�*{�]HVr40�(l,�TcS
�����9�C�~U!�x0:�U\�m�IHWkj6���oT��H�؍y��苲�]l?� Q�s�}h��A*�b1���#:A�%�Ç��=X)rm��9�g#�|HU��o%��^ߐ���SZ����s�e���mob�<�֍!�8Qʭ]/	1,s>XR��?W�����*h�F�$����?��৒��Tc����%V�.�.���K���0�^T�0q�Jk���c� "�6��'7�$�3Ag����'0����۬XAj�[��XJ(b4nk���l2�r���sO^P
8�X��]�R��X��[��l����0;�������"k�&�2��ʚ��OQ�L��:�ʩ�*<�������U\��8+w.�)I��>rC��gV�����	�I|iYC�DK�"B˂EY$T�q]�`�s$$����Nf��x�>�
(G��y#߱�(d����h��,��Y�Y�E� ��"B<D۵.���b?|��>8~BO�<�I�_WQ��G3�&c�Q��BJ���j����ȚsEY_�=O�sJ�ER��ԉ>!�����B�Q3�#���Ѧ0X �H�W#.n�,��״���J�U;�j��.z��m���3�b��1�&��Hx&ABFE�j5���%���'�bz�e]<0X�Pb����jP�+�(�g�͘����srY(::<aҥY�Babk�@&��F������I�s�ͨC9��;p����h���:�m��-JP���[(Q���r>�����"�ƩsD+�Dtr|��0�z�YdB��(�:�������\~B�X�>������&�vĞ��0=(<�I?9QH�"I�]kU����� 7�V�
��Co��xq��/�)��m /�Fa���V����h^Fa���{i���Z��8�L�gjm��R�kb
c��ٖ�׮]����'X*��_5nt1�ҵݭ��.{��T�_C1ml�⁏Y)�Є���J��E��^����}z��q�.�#��Q�;V�I��#+�� Z
wk;�ɱ���Q�A���WA{��E���7���/zs6�������Fe*�P��\LB<aqI#F�����p������^x�Ez��ԏW�Z�)�5���s��y�£��Q�,!�O�lR͊mc�M�͂��ڹ�r|�H���߿/r����&�&�9++��M�w�"9�أCQ�.]�V>͜1�TiU�o�Ҍ�_�$���f֛r���5��	�"D�d=���[��N�f\)�֜�xH���O���H�	�����9���xE�۝�e��v��넖�ѿ|҈B�^V�罗l��ׯ�8�I�����QZ����m6��-��Br���s�t�F�C�1�G�Dי�1�U(-��\3G7��ǜ��AK��7&��z,u���Z��S�Y��},�����v)�q�ĝu����hi�tڜ2Aަ�L�rj��Y�n��t$*�Ty���ϭ]��i�[��J��2[�^]dm�ð�R$/FJE�����
yÖ��v�b��=DQ���:qnH�D>�`��bw����5l�/dNz:=i}����m��ND�Zb	���<*�t��$K[�i5(��	�> |C���F��h��,~1�yee֪`�L�1���d��u*��F���M��27�+Q;��f�f�9E��I#��_oea�Zapt&㫄�iL�"�_�(|�X��%����J�R,�w�!T�6���*	�ɟL&)���{ ���}318:Q:)A�y2�6�Wr��l�w�:K��Zܷh�ZU�����Q��T�Vy'QY���X]1�p��si�R=�UR����_x_��C�8No4
ҚusuІp&M�\�P:W]
�[EK֔�ή����r4M�(%���t�ȈTq��r����;�m�ށԓ�jM`�Ȫ4+Z��mۑfI��6�ӊ����t:1����.��s�>�`Ī6�<Y�A��j_�(���h��$�n:F�ag(�u�:5����)Q�^%�A[[lm;���8t�mS$-��~��`jmm�܇�	ж�B�L�BЙY�
mq��t��Wf��Ĉ���|b\g�!���љ�q}��5H�W��?쳨�zؚ��'$8ed��ec��ڪ��_p��t�c��8Q�J�͍-U��ne> H��\�������D�ܼ~��<z��	��	oMay�,������i�TWS���-�Ҡ��@�?O �?�o���K��u��$�G�l�{`��A\A,�p��#�$J~2N�Ĺ	�[��"WI���!�/F�-��o�/�9�`�ш\�sg������0\�=|AY�Sy8�-��B�bÉ'�Lo�	8商�3��f'kB�V�v��qp���.�1��>�̀�	�U/�Ƀ�nr4�n���B��T���$F#����Wj�Q�ig i(]W�6S ��"�����mۻ;�c��9q1��Q�@Lm2����5���1=�*ry!����9�E���WKW!\C�8>��N� �7�&�:GN�:�\�2�d�"s6�<�m��o#F�����,�@EzC���X��
_Vj�	PQ7B$w\V�ֶ�u��Q�Md�bBQh0*Z�K����U�xYI3��o�;���U)� h����Jx�I��g§EA�� �ܕ��Au��h�j�ʜ�zN-m�tK�&���ģA���E�T��c9�&�2G*�L_����v��[p@?�X�����3�u��sm�$i�	��fn"B5)d}4d��.P����� �,=�G���Ї���T!��c��J��?I�fe����^3[̣$'��I}ukK+�Z�7_�kG������q-Ҏp��r��3,����i��lK�i��V���!D�`���܃9K��Ԭ�]��.bk��D�4���ͱ�teB ýc����������
v��t�&M�s��W�L�1�Gs�!�;Hdh���&��o^:MW�����j[=�� ��ʓŋ�1���)+�6�b��"Q1�}���d/�{$��!5�����������C��_�C��z��ڠ�޸C�?<�vvJ���%�<��	:1�Q�v�ӭ����"�AW�2b-3(���?�{�hT�I+XSh��=^Y��C�2yu��=f�"��!��I�	�[b2�F	���$���'E-���gm
k�%����J{�j��Kq�(M�ѓQE/^C{?�~%��%����^,j������(�[�)/�7�����5�#�ɤ�����+��	ʝ�r.���b�R�6	!�s������VV� �>��U�R6�ު^�d�'U���0�15g��������0��"��֜>��7���{4�b+�iL_�N�I��m�</V��b#�k��{OM�s�OU�dq�R/91�)f�q���b	
��Io���z��]T��"͛r?j˝�C򕩧Am��V>�8hJP-Vle�ϓ����v7�.�!��
-�$�?��_���ϦY1����݆�2�����O�N��e�e��N5!i]x�J�Kp��:z�ʝ�� ���N�b�Q�W��PLܵ��t������8Q'Nu.p$�yRO?iT�N�w���-��$���	1�M�%�գ�܈�v��n �d؀rN���}b�JY'2I��������5]d՞�c��o�B~�rR��bYt���^7�q��$�шW�S�坸]�( 0����Ur�{�LN�4ڳ�}u�Oͩ�8ް1/���MP<&���]�c(	�r���y�V|�Lɔ�O�'���ԣ.!�}.J�Ğs��E�F�)���fZ��1�"��-q'h���g4z�D
���͘�ؐq�jr�S�[���TD���Q�n"�L�Ę�(���&�+d�����7�\A}"`��|zh5x4^a.�d�Q����$�T̐�.@�B$�(e��ܴ-9M��}O��ő�mv�X�=�AM �ij2�z�p�Q*���>"�f�O {0y�']q12��_�)	A``�G(#*M@hs��K�sC_��uhr�תX��o��#M� S�9�N�;�r$�c�=h�ۆ�b��s�������y<3�ԕ"��p\M���WW�%���䩯���K����yVk^��&O��M�)s޼�-v�1�K&�5V�'�9�탑m@���vE,�1Uj�"��Q��_�h��mO���=l�o�,4Z҅D�n�'�5q�U#�?�f��� jz@WW�5�^%��CA/�\�Q噸1��!���iux1MJ�{*�F��������5�q谜���r�y�	� !��֊L3��m�][���zG[d�⸂"��3���AY�ت�L�޳����֐��9=ᠷ����/]�l��"UnMQY-�\��Ý��h�۶�@�x���ڜr*�є��#�0A��e�D)(m�Qiv<�5(�ܴ�����!��X��ܳı���l������ż�P.S�ԞNې&����#��e�#(���3'dE�r+zwSt�Fq���<�G����4�#e�Jƥ������1�l!�;dT�a�A�JPM+�֛~�E"@%�~51����4�s�,G�JNf��9%�2.�e"ߓ?s_{���eg�[���Z�q�諶���9!��^+h�;�s����܉ ��J�J6i�n�R���Ĵ��RC4J�(RW
&.)�Aco��[[\��Ot���R��Kq�F�&������.���RcO�7m���{|,�iMk�4�@��3;>�/>�BW���>$vWVG\�V��V{e�ݛ[%�����;�'���M,�z�)����,nߋ��蹲\ �1�-R�/&������A���>V9ggg���ZZė"�7]��|�j�е���ޞ�)t��]�T�t7]��J����{�z�?y"F�6��[����d-��&�|b\?$��s��6.Mʦ�6�uRV G�%�9
S�%-a�<}*�ԯ����V����?����x�]ǈY��m�\��G���1��H�"�/C�_��d�궗M�%9��V�f+���.BB]X�ya�(h����Oऴ�-�<�Ao��
{d��Pjk�&搉O�"��힔��C��"R��E$�z�	���P6���A��Ƙظ%ֺ�;j_�;��Q�õĽ�D)�dAĐ0+�4�G�A'�I& ���kS�����l�AF2WD	J{�PK��R�X�~���n$�5�H���ȶ
&P!��M��N�l �@&���.�@�c}J�KyQ�ve/���T��>oic���/�P[��ZZ'J$�*�n�d�����7�sE�>Fȴ�/�!m��S�Ѡ�6&nާd蔇eJ�t�y��`�n�����K�4���l����ȣ���P�
�Jt?�p�<!��+��f�;|N�/�n#���dz�-l�}WR��,�S+� cF�!癉�"J�A���i.�_<�;����yGd2r�~,�N?J�.����}R*�˸�ox�U�%��?�kf
�3d������ח����\��b��dY(�('�Q�h1y���b�`{�����H�_����qC[>����p:�LGx�Mko_� ��`�����0 Ro'�ۣ�W{��:K��IѸsm�{�mI9q��\�`+�7�D؅��N��8�c9W����X�jj:�'K�8��\�8ս��%������28���EJ!m/spD���N�]9�#�h��B �XR�B�6z ���Tө��]i/\� ���H���Ju�yKQ��Z�>[LU�z��ww��B����܍c���<p�]�~OY�PZ��t^%5դ>Awp����ھ��_#��DQ�(�*%�m���K�i0d��NR���:�6����E�޷=��A��5��$b�d�:�i���Qb�e»�a��Fck���v;���G�,�C���������ߍU��q(K^�zj��ݧlE�l��V�!�X��D���Ŕ�r�%�q��[�>���Aԁu��F���iL�:�J_Kϯ+��e��c�p��o�Y�&kVz~Xٔ~6�{b��9�e�*� ��$F�*��c�ɾL�B��j�Ud�B Mf�P��,�������T s^���gz�";�PW]��ݭF��:wa�&���L+��byz�:��-A�8��4�����fH�3���8E�.���Vּ���.���P���G�Z�-�T�UFun�&�)X��ib\Z����&M0��V��+Qc��zCS��^�Fix�vI���Z�����_� ��cR��p6s�պ�X&P��n;b 6&�0�j�`��ֽ����Y��4LŲuw��G诠���D}O�Y���3=P�<�>�D9�o=;���]�w
�Bɭ�g�a��Ů��|m�^ mT$���M��`���B+$�y�Z��N����8�Ӣ�D���
��+ە���ʲ�cZ-P�Bt�?!�c��~��_�Ri�g�x,C3;}x�|q�v1E4C�D�))]I��]m�w�龜���ճ9x�[r%Dj��+�<%�������g�Q�� �!�\EW bh�)���'�3�0���s�%5�&u��8�X$�3��&��a����ڹ�5B"���!��bL��n��JH��µI�UѼ�
:�@i���IkI�W�]���-�vۇ(/���̺EkT���7EH��E	"�kϭ�%�.�1ݩ&统�.�"��<w�6��dq�J�P�t0R���B��&G&]�PjE�i��uE�U�.q���Ȣ�-U���d�:i���"�)v��"�N���r��R�ۗP�u�~�B%��!^&J�m�D�kϑ*5��AHE4���EۢA+���壮rZS��;ӵ�6�!���X'"*zpY���N�Y]��E
�4RsNZ�@s�%/��V�e��D�금���2XDSa���V,K��4�F�:,�pb�*g�Q�:s�;�����)Rwq���A����hH���X�,�BH��sZ�!�9+͆��Y�:1��EY�#�IP.	f��|u�{��Y��sW�:�F0�h��\�D��"m�l�kkZ����޷���ˊ0�������o�E k+�h�<�o-�Ҥ%�Ɯ�J��DR՚TMEYE����	�r���%E	4����	V(j�F᦬�@)�CR�C�^j�~���r*ְo�͌�+�t��\'�;�V]Y���
 �o���e�?��u��u}��ƞC��SC�ucr�9G�^3�J]S��9ZB�hI�k���+Y��R����	)�b��&���8�*�{�6�)���Z�"�%�d/PZ�z/(UI����}Q�Y��F����%�Rnׄx��0���>�&F�%���#�Zعףxx�o�����4[�������b�k��˜ๅ�Ooݾ<At+�6�yK��Ѓ�ǒt�
£�pND!��pl���#�{�!e�ܒ\�75�c�o�,D�$	���	��	TF�#��T'n���ҾYA]�]�+�<��`�L,$�#�)�S�vXBGy/�d�TlL�̭�1���[�_� ��/��%�
A�*���a��9��SFC.�o� �fxT����)V����M1=�Q{<zR[�5qd"�]�{ac��	�ݶ)�$;�a�|`�fO)�Do���&z���+�E�H#��2��DG���4�3��{ޱ��1O���1��N�5
g�S)�|��Wu5Y/��t����"��Ӟu�aMU�#3�<����J�Y�Ŗ(�m���Z$�KX��u��� ⱞ/���dƩ{"����S-�46�l�����F�X������:K͊��?��Y<h���;;;҇�L�[���x{������L���S&���y��k�R�Z!��ʔ��T��V�'�sKtS����2���  \&3��pauċe����R�5R�<%	=V��a޻5�4���ab\!%�d�
/C,�o)���Y�&���{���tG�B�oy�/���iT���}
.9a��Nis{�|>���j ��ZY�S?�}^��hm[DRz��A;݉�B��iV�,�!�mq��Zx�2�M���
��)�*��M5�55�Wj���b=QE�&x��0������4�p>�f @lQ�Y]� `F�!����i�³:#d�{lܳn��h�$m+��b���˓�i���zKn��=�+ :�v��Xb�GD�"����ln,��(����~X�D�*
D<@%�	Ć���z̍JO�跘�"�V��-a��֬����97�wl����J���O�I�=�x֎ħ}/vs�td5(U�|T�:���7<�x�+Dɟm���#m����<!�C�50�Ѧ���c���\�9 I���r�f�;%q�i���md��p8G��O ($�{������Q{1�)3u�yy��+�Bj|��n*Vs� ��#%�{��8E�+�R��3Z�=�&UC�Q2b����XB�M��wE�2�����C���B�]V꒽���.��,r�ֹңt#U�p�횑%L�ַ�Rb��?g#R�tsW�.%IW��S� ٛ��U#N���ĸ�5�>V�z�,�����5S�¿�an�{=&Q��y�׀����L�E
�6f���0xl
P���IoK;8
B,��a�;�;��F�Κg:Ry�������Y0s���[X��Q��=5��$���Bx�nAY��h����6"������|�O�TS�R)g i�歕$�;���g�g��A�:	!�-RMz�-L�'k�d�P�;��n�[ y������eg��碞��a��(�#[��3���z�[���(�	����\�*�S�����M�[`V1�*����*X		 �G%)���ZiU�BV"j^�%3����� ���'dc~�+v��s*�1�PT��S�򹕻^z�%Y@ ,�ޕ+��q�[u�M���^����MiZ����Қ;d���5��7&I�/�~�9dSڧ�X�t��Y�hQ�իW����Ф��}$s��ڂKW��u�����MV0��4�	⎑|0�!E��Z8�a��w�ޕ4"��]�C���D�lܹsG~o1DwX_�ښ�\���W��&_#ZL��]�4 �9::1A	�(1ܓ����F�ͭmz�[w�.�{M-=M�=�ٱ4��saB��s��*�@~���aR��N#}⚩��8/{ݚ(�i+W��1 L�������roND׉e�Q���r@k�s[�@�i"b��6U&B]W?� @6]T�Y|Q "��WJʹ�XY报�K�*�^��>
����ll1A*1'��Ʒ� �Q�G�>�=��%�LФu,�����Q���fUkO�ʈ��81{E� L��T\�F,���F�>_��{c�j�U���I�j��i7��s-u�P#hJ��,�b��"ؒ�V!�䁻l�W�#,Y�!ؖ|��(]IZ��w/�5Opt��M�6��1s��:H��^R�
#�%�l���摹��X.�[TH*�\ �����1��R�s'nח9��Mqz��
�>c��fE��FY�<���p,.�i�X�"g�;�3�I�\���!'��1G&����V���/�W�V�x�NV����N���w��ڜl��==~�>�ͯy�3M��:F�K�O��t�S��(絖�����,x���ɜ���d��_�|X F��@����da�?k=Ax�hj���c:>�j|��ĸ�(ocD�-ɝګn�y�JTs�`%�8��j4������Л��Z��1�������1x��!ȍ[�Y�n�/~��4�oK62���]J��cB�nW]������{�����a��J�`����E'h�ՙ�C�Ûm�^��sV�s�� ~��[.̭lM]�~����gƧ@�L�rH+���R���2M�r�)s�w^�~�?��?�#^4=/�/ܠ�����+���GW@,Z+����M:9:�V��MD�>����;�ߝ���P[�6���ɢK����7����Dod�� Ip'�}II�v��v[���7o�O�f��{��ݞv˶lY�d�I��I�b%P��]""U@r���� ��2##���~Ϣ�h�9ي59��e�g�&��wb�u�Qh�� �Zq�J
xN+"� �1��8��*��H!�%�D��r�R���>z�d��NS/\8��|2�+���������hp�0��E���/ƹO>�r�z�(��������	���ŋ�����a�eL�*�r#��Y��hPٖaG��0�G��֓���~�7kqq�&L����y�]g��.-�M���{ڤ�rUY.�߯�����z��h�ĆjF�S�4?����0��!���>�jr�x�9��8Lw�_�^�PB /��������҆Ԭ�����s	WS(W  ���9Ym1���5,��~&��FP��C�XpJ"��nq�uZ��Y��i6��o��>��'���'z��NVi���L�|�p������&?qs�`N3�;���E�����γ��ѣI��=�	�s�h~i�f�<���E#� \`��B��OQ/��@��^�B��B���dA"��%���Erњ�},��)-�j�0Ƹ�����2�=CI�J��.�@���.��G�%X�R�2��3'���>+]��6�������瞣�c��ڻv�'�S^~\����g�j)k榘��x�Q�C��a�#884��93;�N��J,��%�xtW�F�4a4�Nk�����N�k#�V�i�Տ6뎚�+�5����O��?��{A�����4�x��d�����w��{��?��v��M=�=�e�ڵ����^�}Ė��{��1�Ŷ�*=�ߙ���܀i��C}�Ƨ�-f�d5�U�������N�+�����#_��e�a���(y�k��\yWD_�+�����-��cw���AÚ�f�"Z���������n�"%l�B3$Y����1{XR�#Ti�}�jt��Y�M����g��ChFj�� ��8��$���I�F����`�B������]|�dyd
��Œr�uf�o햆a��y���(�3̼�\������O?��'�rI�GDu������B85&V�U�/+�3�W�
U�5I��/i��( �T+�����] �\A��ikg���K�M.)�pD��˨���U��8�\=�q��K�B���Zʢ��*�t|��8!�n�S�ɐ�rj������5�G�����ac��څ���R�$�U�$ɫe�		S�).*P#�4��VT��KF��N�����-kM�eq�)����%ԡʑ�|�D9����QHM�A�€�2m�)�~���8��$<X<��U6��͝��9�F���z���Ӷa�i�'��45H,�|�i0��E-q=���D�D�"0���ՂOl�B�u(	l�|�8�@�
���nG��&�y��;_XwlԦ\��]X��9&�o`��7od��]V��^��'B�C�P�2R-�����Y�L��˚��q���B�j�[d!݈]9�KW�*,���Oa;`E�ޱ_L��
�^5>,�֞߀sp�H�g�=�,Jk�W��Р��D-�lzw��!E!WPB5�ؾ�*/��!\�5Y���w�?��U��������X;���&�ѡ�A
�gee�������]�d�X8]��֦�����9���6=-���,���B���ڂ�i:��2��u�1�Z^$�P�,V �"|���G��:�y"�Q�����������Ӭ�"��	nȗE]��خ3G�mt��q�	
#U[V���ұGkBj��vy��#�~�$N�x��q�����Yj���/��E%oW�!ֽ��H���H+�iLt�N̳h���
!����3�E��G6ӆ�P,���i�I�j9�8��~p|E&  m����]!CG��[���m���8�p�L�4�����Or� G�����Z�
i�j4�!�hx�Ɉ���$l]'��/���0�԰k�ڻ��j1�a4��`��|_P2���`Hh6&�9�ɒ���R�7�˒��A~�:ߞ+LW�t.���1s������� fI�c���YB1�_v��{���Ώn$9 �%Ӣ�ܮi� �i{ؽ핶��HY���
et�I��dD�N�q�A�qن��'-���@S�"�K�yM�͛EU��������0���+-N|/sI����53i]���]�"����j��b
��*�lLV~��2	�ARu%��b)�Ȭ�è���d�Zk�l���5/GB��!9d���� Qo��BhC:��}k���EӞ�P��EDa�A8=hQ�_��)g0f�� E=!�ܹ ��=C\A��<�N	��"]�+���T$%��(�`o������(����_�e��9m\Vj�5��z$N�,F|�>��<,�E�����6��K�,ءiY j/��ժ9���KJ��;uXgg����B`���ϑ����'&fH���3���փd��tw{��K/yN��]@۲$k>�R݊�"Cl���%����?�Y�q��.�#`Ω��+������!�w�f��Y�wU5�,�/qQ��������^��,���B��̕�/Š�=t@�3�n +���\5?�S�r+�^B.S��ly�ZU��D�U���D�
�v���$���p��k��$Ysj��SE��;:�������	���H���&
&����m�S?a.���$�W��}��zS��� ���c.��Z�ȝ�,���l�l��/�\7l��dA���)��#�����9�\���o��cϖn��])��:p��������(H�	:�e��?s���\K�k����Τdu������K1{Q_v�ݿ�rB�����*#�t��%:x� ����)�UKi~`�n2�|Q��{N�i���`�+yv���h�)ԙU�'�&���\��W�<?>������Ú�/_��cw����49��f��x�qP�Z�+�*���db��.]po3z���t��޸Q!a��C[u;�<���S�������JKʮl!�$��Ƭ,Z����wY�v�b̦����J5�in/Nu��տ�_H�ur��T;�%�h���XN�*4���dOE1`$k|����^zd��*�֘7�Ѹ��P��|��ͱ�n�ɯ�W���,g�QL9�4Ѣ����WWo7o�+�H�Ǭ�D'�p�`l4-���*�kK:h�G׆��]Ix6rǥ��f�ן\$�?�u~�x���]d�[t��(
=���J��	2d-j/1�X�����^�(?Xb�7:�+��j`�l`SaK'�ͺ<�QLY��v��+�OE�߅��z�����n2/hz���2������$ѕ�L�k�(q>�]�vK�%y�V.V�u���kl,��&W���PC�!*_W�Dj���LU���0�|4�1���>�)*	Ts��$Kp��1Y֜�H@�&+��� �W��9��06;�,��#��C��mvx�"�'��Uo)T5Δ��˘�r���H�ʣin�~�ˬmKKO��=t)�-���]��2���B��=iЬ�]�s�$8�R�^J��a�a�(k<�v��]o�.����-_ n.{&�Jz3 Y���A
�&�����6�mYS��꽆I���<�d1�E%�BR[4�I����j2�Obc�Ʈ��IJ�?���Ү]�X�=,��϶{�µw��c��u�6�;>�������lָ�#y��)��	�L?����6=�xě6�7�x�����Iڰq�3.a6`)v��M[�l!k8��X�eE2� &ߛ�%�#�q�u�Q[�	6� gϞ�������jt;#�>u���۷o��~�;��������� ձ����>�cǎѩӧ衷�~�o��_z�/�z���xG��/~Ovz���T �‒��>��#��p�GE���g����g��K/�Gę������'�ҙ^�-#[�f�<�M{P��Y]ج�z��V��+t��Y�=-hh�v���IZn�pj0��,Mqq�N348D?��9���͛��G�������#���i�t=�8額6Ѿ�=t��k��χ|@�=ݴo�(gȿ�⋌�s���i��Z���U�|��YY?�b�JI�P.6SEYs����֘��-�z����?�W_{�����wߥ����F6aFK ��Ѣ�g���@���ԃ�T������s��;H��G'���_
r�2��v����C~�o�E�ԁXv�����=t�0�4n{�u�[��w��o��QƟ���̿%��ѧ�|�.��J�ڱ�)Nm�f7gERUQJ�4��ϕv�b�az������5�I��/~֡!ř����/��N,�چ��t$�S����S�Am�����͡�Ǐ'=O�J�7o�}��ѹs�h˶m�9�
vp��	�_�����s���m��U"{���
2
�
�s��K7T�r�l�yA[�B���2e������C� �����v��S�"m����NP�8�ȭ����०UIEp�����)�}��y���L;��e~NOO���,uuwyj�OW�\�l'-h�z{�����H��z��,F.n0�j	m����{о�@짻��2x 6]w�TQU(�I�yA�Ø���^REU�I�sne��`���Oa�
U.Ɯ���m^{2�N$�=s�$���w���@� ��{���'�-��4�*P�����m.|E{=uإ� �E���K]��/�uw����ίpם�y�ꏟ7n�'O�<ݻ{�nݺɔ���ghӦ��y��1ݢd�$��cF�p�Y�E=G,8���� dǃ���K���{��q�}�՗4t�_�#/�!c�絓K�.z��)匌lf�ו��8��٪����6JFS3~_+�9�3�3�5���C۽B�8�Ů=�,KX�+�"yEa�<k�����_�~�~��_��A�bR������;hl�6k-7o����!���OyF���-����s��~̀16Iy�\-#]#�rQfE���Ā�)ܭ� M�5�s!>���A{��e�%�!��KS���q�T'Gs�,{4��Яi)�P�
!Z$����6od����:~��xj �m�Zǩӧ���mT���~ސ&_��?����S 	��OU]�8��!Y��w�f)�lĵS�"�q�JTE�D�V��e��e�P��j �%���H��\���0�km� 
}�����-QĬ�JS"(v�\k2�n��d�r�_�4���(B9uF7�ȃ��@�+�!|�"/����2�'�h�p/�2@#[T�ꈦ�;{�e4Z�~!.�S��Z-</�����O��;f���7m����f�lg�j5�6I�_|����C��� �d��h)�y�;yW�M�����s�L�ݝZ2�$'�&��@�����U�K�s��J��8�T/q�0�)ҋ*���Z�\�H䚈�~��>4ˆ!�h��x��}.\���7䰷��r��?��&;D&@�|9��T�&�!�>$�E�a]�+�����/�c��v��;�Ax�F����qn��jav������0���[YX�����*�nݾ}����;\o���G���c~��U�(r���o:e5���$
M!����C^N";���lsMM]c2�5�RƵX�XWGIVEEC�)bgψu�k����I����N����4���<ݹ3Fw����~@;�����"�7�o�|���Af;_�݆ɇ���E����	��_���ݹK;��.�/�{^u��^�4z̅b{�A,�t$�w�����F�O�*�qȽ.oc8x����7K�$o���H	/fњ���"kjŬ�,pӌ���P�E�������5�|���S";�ɠ��?�ȿ>d���>���:w��x����k^Ki�w��)������ϝ=�Nǟ��=���df�~��3o�@��<2���������`LQ��c�'�ې���͛7Fcr�c���u1�B���"���ƍ�&��V��@��BhW��qFY�[���gS�7~�3j����;���K��ֵt�����~��nڲ��4��s��z���)���7o��m������B�0��/�B7�^��[�r��4$g[��u_�n�$�М m�BH뾧�`�����h��^�L������7�]����Jp��I���)L�d2J�����%l��o���xgw=E��Ӧ��ğ9y���Qֆ]�k�N�qld\D˿��2����ǏӡÇ�>��~�6n���wn�	
|(/?Qd���QCq�DƂ�ͧ������6C;	�`���cw�!�X3O�9Wmd�f&2k�!�/[zMC��%��su�@8�u�W[^�.����e�\�]/�g�|8A���
�\Ԃ}`]�7o�Bol{C<�^�?��~H6�t����ܽ^�E���I6L��{8��i(�F�jO�ր�ooϨ>L�p��f�\��QTl�|���B���ڮ klJ�?a��4�~fz�o
`�U踷��n����[�Վ��IZ����z�5�9W+��/9v���&�"�&*��V�Lu��Zxc� �y5qK|嵭+^�9z��ܿwOZ�utg��"J��*$����>���P+�4k�k84�T�SX���}�)�.��X	���������m0��X�1WC65i�����'�����"�,MXH�<$YC���-�W_�~�h�6S�����T�nV�2T�{Z�X�o�x���2&*���2�g8=�?�\��������޽k��%M#�K&[9���0�̇��5��q@	�t>˂�[OK���v����o��4=�����o��6!�Vh�Z�l�k#4���~�nr"	���G�a��\c"��R�+�6��I/�^�Nz� ��#P���*�u����1�'tP˭Qvg��i�JA�<�%8q>p�Uo�/�F�&q�"q�5��������O~��Ң��z]}�&B�N� ��<<4��ŉ{B�?�e��W_sh�TjWݠ�%uG����ʵ���o�����O����],V�v�`�uh�mރ5-�.Dp��Q%G�/Ӥ����o�O
jA&�
8��ޞ��D�~���f��_�e�������}�����u��2�A|��ȞG�yr�̗vHi{�d��)��ڗ��:��4k`�C{Z!�ր����K��gg=�Eܦ��ݻK�w��_@�Z������Qa�[�N�Zq☳�q�� H��Y��+WYӲ�+�
�:�8ǎ����}v��������χ��*c�ט�&�[�eg_�ܢ�/0�D�zZM"����)΃%�����w�~1ޜ;��\�B05����;�,�1L�ƍ�L�'���M�݊��J�%�{�Ȥ�	����9�-�L���|_$��ݣ�鋳�Ӆ�.��M#t��!Am����[��{2�����=}��m���9�?:J�����D�B���	�Sݾ��裿|@����y��W5�����m�m^��0�3�\�����\�o�h���JR]D;{�m�@37�Г�'M��^e{�W>�}�$c@^�����NÛ�Y;4ӣ�rע,:���xt�Y|�K5u�J��!�g�}ڳ�?��O��u�[�p�M{=��o�a��^�}��1:��__�|�;)��?�OI!�|��/��2�9s��{���w�66>μ�it���%S���k���V�~C�O.��R�X�X��}�嗂ܱ�ܡA]���9��j�� �iO�&�ݪjoPI�Xi�q�ׂk��@����cGyr���8�Y��{{z����{�( �0�� 0�H�54���2�P�� ���2{C(��_�/�en�%����]l�Fc�QЗj�����a��Q)Q�ӊ���#_��gZY�Z߂��mᨸ�%-&�D����sž8��3�h���t��ֹ�9�%C�<o�ĚϲjC�>����Ň����O�c{yY���f� v�����kfZ(J�Q�dq���i�J� '�bea�fc�Z	�Z�Â$�kշ�����m�
��(A@G���B=�)�:Ǣ	@+N�y���� ��]�K������bæZ���7�J����!�;&vg!Ӿ���e�0���������D�,(XW΅g��=R�c��*�̓�N|V��~Nm���%Y�/��.�99ět�7\�32yw�k:�8����dJ�cc�MH��N
�@��P��g����T��Ɓ_i�[����jKag��J��H7��hra���3�k�>��m'Mb(/��,���^Z���eE�gŞ�U��G&�M7�J�X�K9W�Z,�-�ھT㴧9\lBw¢j�~Vxr]�|��J.)������);)��3��+ �K��)�8��'�^c����#���;c��M�D �ˎgAG�-}2-��Y'F�a��ԭ��֦��Ԗz�6&v������m�����HpU�A�,�u�����=^�d���y��"��=ӡ�}��@+M�Ak����H��a�p�>�%�Op ����[t���R棰�*�o��oi~n�)�c�s������eUAyxN�x�y�������Bej���.f]0�bᚻNTe���`����ʍVt��Q*�в����~�������B����^�j*$(C@~��g��1v/�cX�09r�8����|��e��Oz�	/��\�,���C����F:w�K?�3�Oڹ����u!s^@���Ů\��.�_�����ի��}���?�|9�ة'Sls�ٯ^��ss��-ڻ{/U�# ZЪ�b�8KkYgn�`���QXNo�l��e���jb�E:0�@��XE& ��������1��[�h�Ν422�I�G���v4���/x[����L�X���N1�!�*�%:XfU����\��E�hHSy��6��-[����,C^z�ea��`Ŀ��ijz���'G����dq��)Oy78�6�1@��%�'��5���jY�@QW6�IL>c��9��������l�tQEz��w����Z�|��n�'����E��.��o���2x�_ë��4�{��5Us]p���$�0��ǎq�-v�qOa����IW���#���~�o�����~���M����7������l�\�|��8@��s	�����~�c<e�L��"/+�F���'��`O�Zx��YKi���{Y�<�Z�~r�߱�qx��򀅸�')���&W0vɵ�$��W�6u=u�BA�H����Պ
�LUk��*�=�R^=��/�SX)�9r�nx*x����a�ݼy��ul4���:��i���rd]����P[��XU����,�J䩋ř�C�%�u2�P5.�����-[�2+飮B��EvgC�ƮDY\���[��١R		��{��7LMX��?��'�Y�XU���b[`,H��OP�YƑ_ⱌ���q�U�s!�po$�W�������\�%a�R��fk 3��j��� M sa���(��t�P��70�g�y��>�<����ܫ�+//�x���y�+��������� ��];w��/β|8v�hJN:�U�J�5�����Ԧ-Q���"3�Z/_���d����:�j������6m����g?�g�z��������,�0�S4����p��֭�ͫeB����K��u�Y1z�����Jc-����CL��<߇�?7;�ٍ��|oݶ5� "lZ�d�?�݌�2�;��< 7Ck��y<<.H��I��7�������_�С�L-X����Zӧ�}��xP2����� \�$��Rn�c{~�b�=£܃��SQT�� ��;����0?oV�.p+h#��u��	��燠 I���B-b��j�Z�+8%��\�f��VW%�\xhnu���g�xr&yd���߈���Ѕ+"+.Ĳ��H�~��Ƶ�t��>.��>w�4��w�`���=}��� �x3撤�wߨW��cd4K[�GGf#Bi�Jj6L@�A_Y v*�X�]r؋I�������3�p�pO�0q��?Y��Y�p���=qf���"����i��!���k�\j�Sɪ�?���e)��#[6o0���X�ͣ��&��G��"I�J���o� 	itV��T���X����Tė���֖kI���,[w�s��o���i.q���ơTP��-����iE'3h�cnS��?��U�}��^ظꇫ(�^OjOk
!s���W掗�@%K������.����!��#
�sp�(C5o���ũ)~��͒m#-ԅ�]iޗ!q�S3L~��#3x)����s��.��cv�4�������Vm%ѩi��5�u��G�]w�LY\0��-![R�q!�~Nn����hKH�a&;;��6xȐND��\��/=_2����`K-�Poi\���"�o�lJ��;�
�����!��T����6N�F~i�v�J��e^m�\o�]a�"�O���񺍎"쨕.}�'\�3D���ua��B[���7k��B~��R��^���n�V2����7X�
{a!>����ߥ�Ϟf�B�·��sg�l2�3$���[L�K-

���N7�����!�/��3�;C?�Ꮘ��d�MC&
V`ݢ49�V��4@`f7�b�_��hc��Sc����.�&¬��Os�|�����{���\QhEo���(���%�r�@�-�oE�m�Y.=zC�K'���s��L��8���\�;t�Bb{	`�Nٞ���T�$eR&K
��As�d�����cm���N˟��U�z�Cf<]~�5���%r�%Ub��5	�����������G�A����j�4�\Zf���pI�u���v��o�ݻ}�ݟ`�ڱ�S�����?�E�8::Jސ��W�3|�W3H�޼�a��uղ'&�֭[��I������1���t#��ꭄ92�fV�+�.\�C�}�;�BV.�:}R����X�Uo-�Z��[�S���
e*�#��JN~ږq�L?5=C~�O��5��d��f߁����&����nߺ�^���;|�#w�:�|�k�͚^���_~��=̮��µrg|�~����k�����PN�'��Dj*�Nׯ^����M��ũwZ0Id"�j�֩����q*<e;�Я!���xTR��B�.yæ���	����,HB)Ɵ�����@���i���/�,����}�u��r�gtI���Ob�!�g��B�A�5�駟���A
�"T@m��<�T4L|]m�v���Л}�Ν���|L���d��@�1j�&-Ɯ�����nݸI;�m�>��j�3�X&��g���'��S��_ˡg�$w#���A��~�,�*���V0��Wj�7m����B[�|o� R����h��[��՛�X������{@��>�A�L�T�o��o�;<̊e�uT�>$$���; ,]<XT�^�z�:���S���
=r���6蛒QO/|F?��/���ѿ��_���@L�
ˇB��/~�Kz���-}�c����B�(C���ߢ��^��S������t��U�$��i�s� �Ξ[�j�������*�r�S��3�Qg�j���zA̢�E��{xdM�W��PW'u��^�����U[�h�����EޑHzˊ"hQp�c��9�8�E�
o��`��.����&���K������H�<�<7�Tշ��p o�Hp�#�`�ܙ�w�ʹ\���&'����`�9UL����K���S�rÿ/��r��3�G�l��%JG�M����5-Q�`Y�=���v�8F�"=�°�����	7p4o/�␥�H�4�f߾��E}-����cw蓏?�O<{X
b��m�z�}�9)�l	^^8-9�N�kז�WS�1\�Y��I���6�,\��XOEdb�S�����*���Y��@gY�F����Y��2JJG��7r�w��Ӳk>�.#߰����/�ݝ���Ǟ�_�"~�
fP����?O��ߡU�������/=��^S��إ�g�(OҩS'�_�.,�sq��=p�*	��z�]�tQUu�c
@k�E���HN�g�7~�����G�ywpXMQ�%!3G��~����"�������H*�$�%�/�R�Iq^��� ��A��S}-3�
2g�q��	MH�������5U:zh��CԷuͣ�tq��<�k��%\���.�����z�嗘� U��4?���h����-���z������=���rΟ����2������6 ��ǎr��G���<(��S��� ?���Ƚʾ��~���� k������K��8%ɿ9���Ȗ��������]{uM�t��I�_QC4�׈�$.vB/�P.`vպ����4t��q����A}��	Id �������
=w�Y��<��~z��W��z��	pW�v` I�Ѽ�o�៨��L��Y��i�&����W���#�T\��;�C�G�'v�������=�M�F����RZl&��>*�7�6
j06ѕ���O��Sߙ�0��в��4�Ή1�7�PJ��P�R�r�7��4"~rQ�Ɯ���,���jh���~�#���Ѯ�հ�2�LLK�����fc��4l���$�B�J XK���F�"Sj��M���
rF��Y�xR׍�s�Aj���L�U�^�rx��Aj�d=(��8﷢����:5�k��X��U���J��x7IN��LPwc1kd��������,ߦEv�\�|p"����ŉIFB��	^i7C.E+��(��ؕ��m��}���Y�3ۊ�i�~��M�Fq%����C͚��S�IŸ�>����s�Ʉ��?��st�����vhoCk {&�1q��Z����LYD�P�g�Peն��av�
f/&~��Xk'Rg��ou��m,KW��d�\b�:x�T�H�*��/�%k-�Ү�B�I��hWJ�y͢�y؍�-/�UL	�nᕭ�T[\��$��J����J���������-�^�s���nb���p���)�-H�eDC�2~KJp
t�>fl�+Xۼp��mK��4�����$�w���d�b�\"K����8N�{6���|��K�����,�SG��d��t���"L���X��x��g0y���@:�� �d-
H�J���c\� �VFꊕ�ڬ��X��wJ��5��&�T��hbG� �L����vgdg����8Ν�\&)'jJ���!�y)m�?�n��
�ڜE[!��
�p�N]�1���~���K>c���T�N��K	k2�UT�-8�J��3�c�Cy"�&!}ؒ�6�B(��D0/n0�E��6�c����łv��.m<q���j� 4��i�X�9�R~/�U?��]��(��0D�-ZB�󳼀�S�8L��XM^�
��@[1�#��ΉI�J�(�"&�5�dQ"��S�UJs�Z���pD�V����N�<����T�&#�6�?�� U6v�j�͡5Hj��U=���_w��eq;��69��n�!Ι�!�9�/-d-/5:q�&b�����i	�ik$�f)߇i&����-���Q���4%�s�5^[;��n���p�G
G���f u�wv�S>��o���D�j"�]��
yHI�bE'4��&�M��6�AbM%,Q>����"�h`�i�Ѫ�P^B��e�Qɂ�A~~�JI��lٜب�xp��W9#�3���>���a��m���|�h���!��QC2�U�f�:Z�T:Q�#����N�+6Pr]�9
��c�\uf,'l�ɭZ�E'7��79�r�!�^*��"��Z�E�L�#e�_��s�]��i��u R�9-%g�\v�]�&��cEk�(��-K#+̹TV`�$N�5Y&6
:�ӝ�j��A�6^���Pm�B�,��,AR]��4[YJM+X�y(h�+�A�CN��(˛D/��I<�haSu����*�� ��N�1;�?�$����S:����?_��=Vequ?�r�-�������7s�u��49��z��u�s�V��b�����3늇���e�Y�:xJ�b�ֆX��Ɣ��!R}�X� �ǵr�B�f��ԛ�jz��9�V��|���Lf�f������i�j�ֶ �
ʋ�� B���n2��XŦ�ӭ`%��~�#RwQ�d���]����N�J���QH+m$0(U�[/ɷ�ڮI�i�vO�-�n�Q�N����N��o4�i�M�"��(�ޕ�����|�W!�u/Hr{�Iȴ̝�p���5R?��Q�JVA�%����&P���<��E8/�;�N.�k�!h�в΍�rsԭ8c� ����.R˛̈ҿ�m��Vy(�L�HR�0��N���Uۺ���Ӣ�3���m0L쯡`����.��U��Hɔgf�����gŘ�$L�_�h�cZ���)9���\�c�-�L���x�־�p��n�Őƕ��RP(iH��?Z��E�z"ף~��)	�u�S��E^�a(���ҪΝ�Q���SIv�Y���ť&�i4��5����}���b�4n�Fw*ݧɇk�A�j)�$!s.��E�����{�v΋b�S�����6��'�S�j|����
'l:q�( ّ��:������X��^Du��~�zv�ד#��G��[��RN*�wd��X�b�	�[� E�w\݂�m���G�R�JY��,K�	V��cmϾv�b:c �.Q&Δ���jr��-�-Fa;���,���6�����LTέ�06nC\�VC<2�<*7�΃�a����"� �$�[ӚG<��[4�5 [ˊ���3kç�W���a3k��*�̓<z�8��
��07{L��!�lĆE)�Ar;G!摖mފ)&�}'�"��&�Uȧ�;��o�om��k�Fa�?�R'���wc�D؊B=%I`��=3K@�$6���^��yHI��ՙ��@͵�tK���z�jV��b�N��m�ූ��a��zHD���ʣ�3Q������	��dP�yv�T�M?���%�G�0������6����QL�0�Z8��1�{���o�T?[�+w]��:��*�*\P]K*��WX�A���>#}HvZ����H�K�\�JklsI�Q��.�o]���k��x��,�~n�d���@:�M&��D	s��V�)8U�<PQ�e��Y�(�R�M�$jY���꾓F�5��ߦ�d���Z��R=Q��5�A�$��.\0�
�d��Z������eH²���Vy�i��X���u�0f+zMM�I�Ǻ����`�T��A�֔x��Y��(k��x�6��vG(���F�F-���E���:� ��Ag�0����uj
]��p����{�ɑ��ٙ!�S�2'�E0�jR��yh��'��P��� m>�oc�A���G�;�2��	�F���BYLN��B穠�T=8��{r�1ת�C�3v�6n`�ށ~�R�iWV~P�s��ȵ��ay�gp�����
����ѣ���������--,���0�!���{2��rZ!�%��Ѽ1�z;��cw��2���RP���;O�f�3'?Q�	ۇ�id�F���o��/�BP�=8����8F[�m\���@���%y�-8XQآ���T4q	3Iw`-�P��>� ,�L��g�qy6�pQ��c�.F#b6��Ď%�s.�se��y��ˊqf�E����ׅ�S�����皾��>?Fg�����Ο;��0�pP@��Lp
4�G�(�O���`��K\�qp0�oE��M<x�`�������8��8�h����wfj��͇7n�[�oч�ŏ�,�y����!GA!A%Z���ku�����B�e?���k�-�'O�`W@�h��^:u�U�n����4����`��]�˾�ט|��Y�>�?qo�F�졮�^���v(��%Y1~�7`�1 ՠ{��}t�������mz�]���E�փ*�ȿ�������
�����^y�Uz��3|���F1�z�"��)-����L�
�j��`�ܴ��+���;��Z����j�D��̝j��W����s����� 
��e��0�(������Dn��� @�uPpO Fp��%����Mbj�'�ט�l2`v�D{p�����������&���������0t�%F�
w�i�t�g�[Q���!��-J$��N�\�wa~���߸q��Z�q�� ]�t��:�u��Kw�*m![��S��%A�����ڕ��������366�]FF6�=���넙�.�ĵ�1�r
��_`�@":�Y�_�{������@�&�����vڳ/�z9��Ǟ������&@یL7X�&a���k]�NT��e^�)�.?=�`�߾9Ʋ%\�`��6�lt<,XX��rg|�*�H���橢�Q<���#�<Tp���G�R]o�׏<�I��勗����ڶbq�?{����w u���ԓiOM���+�(�Yi���VN�~y��<���G�n-�"��f��;�;.���р�azy���)@] Z����kO���b���w�.����l�����=����ԦM���_�����^}�5������k��n���&�˵"ԁ�R7�r�f�ܼz�j5�������t��uuv0�D�l��NVB�3�aPo�U).���5�-�4��H;���E����M~A:�����3?�w��aO��X����Ȓ�L��e����釬�c��
���]�L{FGQ�����y��b�H�z�c���k���o�}M>~�؈��?�b����Nf3����?��^=�����P�^D�1k�~" "P��M[���$w��|��l���v���Dz�t��]��1^��J��G,����_P��L0����q��Ӕ�O�0��m����1��&�6��c�:���7 =5�� 	(�%O���'H�	��	#��4<<����~�@��[��-?�c��0�	�Z''����]��;ζ�*{�rS�f�8��PVg�Mi��<P&�T�]�
H��6(��@�h��T[��kv�W�o���|�kzݬ���@ol<�Yjж����\�ԹjUe�kV{)a|d�Z�7��A�zp�>?Z=<��3�|��6"��a�`��?:F	�����pL����
|�-g(�^x�;�|��Ǭ	�����]%�s��d7�W�=�A��=�F)�+T�./�&�-Pk�@�X�-R��@-�� π�����=sP-�aSU�sA+쁁K�s�S$y��4��"�Ф8u����@q'�e����	�=L��ݧ��ׇ|�Ͳ�ْ��Y�2�;v f�8h�h�=�Gِ<r���h�� m�8���M������~����;6�Xo5}�f�P(Paq&���DP�{=�V4:<(�{ Rl
 ��.��+X����lP�q>�V�A]��|zb"�U�d�xYE���ĝ6���C>�V���\h3
����؁`Uv-C VD�c��Y��O�����v@���2�d��I1������"yM��c�>�S�������A����^�*i���r��>4f1D����î�:���񋰸$(v�G�~���:�Y�t彁��Ѝn%_�T���(��Tݵ��"��XV��;���� ����>�1�r`M�(( �����۹Q�]�K�^!�x�O�4�ۿ�SI?��_��R5���P|�]�3�D�e�P!���V�O_��Nx�㚗a�<�lP�����gՊ`+�5==���]��ĳ�<�I7Ri��EhNi=Z�ֺ fQ��a��7���� ����nO�PC��i«���Җ��x�w{{j��~.�$	�� ��N�����'���7fh��m��~��_ѠW�a|�c��-5��Z����\����-���<��Ը��S�T`�� ���Xx�:�?�����<c���,�7&�]� �Y�.��'����yԒXV�*[&��YGN��9 �xk�r�˒[^f ��ĉ��fp���2U�6q���|+~������2o�^,��̔�����=��۳a�qv%^��߽O�K;��|�G[��G�i�N�n��d�	���`M�~�OO1�&y��~U]=]�-����C�5�� c�A	/pM�pekW�_���]���Y���-8���,��G6Ӹ��!@/_�L�~��ݿ�w6�U�mصೋ�{��	���E�����gOpU<Y���c�,,+���$��ħ�4�
8�v�
�5y�������mݶ��}�9��[o�W���$��q���`
�Z� �w���=˪7Tn�%�>/�7P<(���;�Y�	\��4��/Hr�Y��]'�c��]�ʞ�s���o���;�-����������� Gh�[��<���I�Ȃu`��)pG�nc �$��\@W!�ѣ���]N��׹G=���W����^mF����?p�
��/��u�=���_ee�7F!�aM��A)��J:�`�q/��*#I�k.EMjY5�+Q�"�P4�Kj��L�����t��s~'-x���wӹϿ�ݽ}��t���bڳ`��z!��'�p?C�1�l���l������.ܺc'��K^մM�Ij�
�
Kl��_�p�S�j��]��9ׯ]g,�-ޮ������}�?4�<��M0�	o'!�������HP,Ӫp���������o­��x��:����s���{dh�0�>��)|Z���:��Y�?F�lea���N��72����(��a)wV=O�Aj��-�p��Q�4��:=B�\7�<dA�&YfHW
�y~��ȃ\:x�}��gt���^��o�ځ��T]�,���K�8/�����l�"�^˗��~Q�zJC_Gg;�[�����
n�6�(N��Q��W-����=���P&�i�8�'r`�l����vE��y�0_~�p�#�_e�����$�g�-�*�8�����7� �{�b�l��w쐟�N/s��\�c�!R�l\�vY���1A����%/&i�ˈ{���}=������t�S�j����s�<���	�q���E_���h ��!��c��%A|w;$9bh���;�n���$��^/KF��g �ە6�� mdiq�n>��w��# �؞�<xP��A������mF�_�C?�w��t�b�
0�XVX'�p)��0I�5`�m�~����r�+p������/�8�x�G��ܾq�Qc�ܴ����m���]@�|8,w����]A5䚸�\��,��Jg7�T���ϣ��=48LK;���=4�_����lᇎ'A?��^�#�)^V�^?q���EU����lgW~V���FX��q���2�������wqם� ��Q�M]Q�k�S^�aQ�a���J��{������D�������v��v��F�����(�)@b����F�	i:U�mY�/���'���1;	��@לo�!e�=v��GxbA5�=<9�Q!ɡTj��莃�����������Dlĸ8"C:x�繟�<���f�,в��sO�3lz*,�G�Zˢ�� ��]��Ӂb���U^���9x��u�W
��ɚ
vRV��Ѕ�n�̶$UfI])Y�,
"s�^G���v��_��2n���5������O�"��� b�Da\6V�h���eԓ�*,-��"򤽍툁���� `Q����q����lȘV� ���n��<ec�శ�a�J�[�XP�&u��hL�36p|���<,���p,DGO�'�o�O�"�5�z�����|��-SW�6��YE՞�p������~��� Vѝ��װ��ׁ��
kX^`s#��Bv`*P�=�m���H$��pl�ވ�rd8�K��2l
�)lBll�Я�iQ�J~��,˚��*�H�I�CfY|���#�U��݈��8ǲd�YV�^P�1���B�eg��?Ь��< ۰���O���=b�Mh`pC��������kI����d>�����,\����͔֡��l��e�мi�~�XR��dʚ.N�����0œ5�_E�z�/k-��������݊ICpd��Y�v5������q�*ٔ�9I�����nP���|�-�� o83��Axs�OP&��-/זⰡ��	P���PSbzy�:�K���뚼�c]��M��i}q��� �=l\���~��rA��q��Y����Ⱡ�P�Q���D����2�1���&+�L�
c�DP��m{L8�rq��j�!��(�+����v9/ת+Z�̨?V�:!�ׅp�m�"�]�Z�f��m�vpÀ~�L)�5M279_5�J�[	!����������#Ƌm�-W>��%k�W�,�Q��0b=��Dw��0LA�KXJ��ĸ�����7W��W��2mՑi�bE�^�T��-��Z�|\
�N7h.��p�O.:>'2kƣ��%d��������E�C�j��/T���̩��T(���1�X�Κf�;�<��ܢ�U����ֺ�mw��$)�+�����$'*0n�&@ƕ�_^R| �j�j*E���\�����x��4�F/�-'�&I�9�Xw��O��)�.�
QQ�_&�/�����5���Թ�Lz�c�a�&k�\�+�[Q� |ε�E}�:*ժm<!	��4}�T6��F)u������&�����ygU���b��z����� oI�]��۠�O���X�B��.nv�h_�]��8�����}:OZ��le#b����Ws_�''k�b��8~p���LvgK˜��b�`���$m-����NŅ�pB'9ˬ�(����9DVp(�@�I�m��k_}x��P�$�\S���E0�¨��Bh1�]�U�����QќZI-J������h���L6�ǯ㢁��E�Mg��f(,���r-%K7�z�<S^G'���ː�e]��%g�"<�xeY��b��]m��f��.t����Ƈ�Q.G���(�^��Rt+nDE!��48cG������!έ�i�u\s�h��nWp�xM�EP�;'��$�=��'$$���g��.hN�y��E�4�"�4�����J�i`�� &F@iva��+��b�3����u�����#�2X�jG�3�Tcrs�Hh/�0t�UQ����H�Zc�\�QG=��Aǜz}��$J��	�t|�2i�lx��H5Q�4m���Wctk���`�|U._�
���l��YW���(\�w�Q��;�(o�X�hlL������A�(y0xX�߫o���X��5ːT�;�/g�{v�d7���6�0�n
�奧�y[Qe����$�i�P���O>x|cJ�-J�Qk��cu;D5���-���m��\,�@��|e�Ч�,��G����0j�V�\I>[�����6�� �˵ؙ�H�3�g6f�<�R�Q�/KǓ�A���b��μ,�Er��)�5��T��֠jy�̡�r�� �N+i-��< 6��l�D#K�Z�%���9+�W�J%K�S�bzݕ*oLf�y�R_]V�.��WP��2>�^�,��xHq;Pj&�y����`Y%:��+4/�+NH�����2�D�����'m瞋~*#-+3��e�6�E��RO�:$��x���Z����Cxk��I�vv��B[g[nm^�zU�֬�R��"�� q��:K�4-R���$&��r��%-��2/~�����$��^���J�BNo�C���fN��v�	����8y�����kxR: #|+����@�'AN�VT�K*����a�;Q�MvvQ��@����a�R&系FUl���K�k��P�0tQ�P���.HGG�D�_Qг�E�v�s�@���i�i�uƘY-�]h�]H������~�-�jg��&���,����0.S͸�{�\2���3��Bn���p�M/.�Ȍ[�����5a��6�y�tf+�8C-9����-*`O�����Q��\�L��"���^[��[]!���W�O���-$��Oh����M2�@�"h]�L�.����V�2d�[)y�X�c��m���Y`�\�)�e���K2�/�Eܻ0���ιv�4څ��?�_Yc/Y�œ�K(�YR0�
˒���	N�U-D�qc��b��Xb��md�V�KfoFh�л0����-L�W���)� �Pkaj�3���������g{�w$�@Sv*t3�yY)��Ei<Īz�-�i�pQP(V4-���p����K�FZ�U���k�	�IpM�(��ge����FG��
����m>���l%�[}w������s�8�"r8�n�B�4S���&�7G��[�e���6�����p��he��0FMWYE�k\Ҷ�t�|�%��Q|�����*crk�4+/,��r�Dҫ~�ʻ����q�N�7��l�G�Q�.np��t_���K��vvI�6��wF�����Z��v�5���1�^��2    IEND�B`�PK
     mdZ���I �I /   images/ae036c7f-e258-4627-a75d-99715ec815e7.png�PNG

   IHDR  �      MI�  0�iCCPICC Profile  x��||eE���6�G��y�]�$�{�R�f�IvC�]�%�l�l#[`�H�"Mw�J�"�T�"H�&E@`��3w�N�]������@��79�Μ�=��{I���挪&��y����L��ǞՕ^IF�u����X�����#�Ox���{�%��H3������;sp�@�4,¯X0��Q����- �~��{?G?K�0��g9z�xǓӛ8���V�)�V]20}�n�$���^�0IV�O���Ṡ=a`ͻʅ��;s�̙I�*$�̚�x��ci̹���A��$c�Z�?<+I����{�\�FЭ�m����%�����<���L�Ze)cͩlf���:��լ�y��C[7MV2M��4�9�5�kʴ\����Ӕغxx��6���Y��"��t%,I��]�*��,iƫĿ,1h�HZ��x�*��&��;�%��I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����{Hl;�$i����6�Q�\�`��}yl���d���䶶H<os
�R�^�e���vLrjr^�<�6�-y y2y5��a���D�.{7�pfõ5�6j�Q٨�u٨'FWF�0z���F?3f�1�c����M��{�������J�4o�ߎ�x����<q���X�UN�����U��j�w�ֲ�-��կZc�5�Ys�5���'k��k�θu�Xw�uo^�{�W�?�~��6��l��F�o��&c6�vә�m�ك�[m�b����R��~?�-��f�׶�f����ŗ_�撦��;�֫������fױ���`9G�g�.;mۮ�������p���|�̖�&������4~�;��~��]�w���ִ�Zw]�}i���'̘��5���s�7.��ߞ�w�^o����3�ۇ�:b���6�7<�w�6�Ȃ��wZx��K�?p�����!�~w�CO9|�#N;j���=f±W�k�?z�~'�;��S[O{��#Ϝx�o���ܕ�[~A������{~���/�����g-WO��랺�7���C���֭o_�w~���w�u�=�w��>���G����d��G<��s�<?��/��ʌ�����oLzkǷŻ_������p�G>�+V�~����>��kWrQ�aCo�u�6u��7F����5敱�[w܍+�3�:��o����q�������k^���k߾΃��y����x�57�������MO����_}�1��&4Ml�b����Z��q_>{�˚nn����W^H��>�b�\S��76���m��j�ݶ��C��{}mA��Nk�x�umw��ؔ�v~��cw٤Cv�:u��.����Wz�O�r�λ����=~��/���7_�֊�u�ڪ����͜3�p�f}g��C?������s�܇�=;�����p�EM��[��{8�t�A�|�!˿s�w�;����;b�#�G���|o�cf���#����x�'.��U']{�/N��ԫN���K���r�yg�u�i���Gǝ{�y���\���2|���ɂ��]����.�t�V��uE�\��U�|�Օkֹv������冎w����C7/��!�}�I��s�%w\��_���>|�ӿ{��7�~�����}����O���~辇��í�\��������'���'>����������n���]��U_���F�<�o+��ګ������׶}�o.}�^����<��'����m?��Ã����n���c��_���a��Fm2��Q���Yc�{ĸM�ݱ҂�ی���wU��rƪ'�v�ꧭq��W�u�������/���Fo�ކ[m��ƻm���'n�|�;�O~�/����Ħ-v�r�V{m��ˇmsJӏ�^��+���gϱW���ߪA�dV�kl��W7�n���-;N�ڷ[�O:����?n�f��Nyt����٥���ίN흶���]/뾻��cfL�m��{�q���o��[��{���x�l�m���}�f-�}���^���s��Լ�$��1��B��m�nKfpЁ�/=�퐇���w�=l��7;��v�nG����}�ǝ��K����[N�������ϝ���/���鯟���>�ݳ�;��s>�ч�~p��x�G~��A��$�|�����m�.���/?񊣮<���v��O���k.����n����w�#7>yӳ�|�����[>�������z��l������~W��߾gֽs�s�������>t��G��GN|��?���鏟�������>���9�f�_vyv�粿6>��c_x�����ˏ���Wn{����������eo,󊷮���8�����{o�k�k}8���Ώg~BH�#�Q�Z���>�ר�G�ї�i�_{Ӹ]ǽ����g���ʯV~�ʕ�^��٫��ƅk^�ֵk߶���>����_��FS7^���޴�3��_ܲq�/�3ሉ�mq�m���o�n�6͓j�}e����v6�D\-oU��G�3�o۾�ݘ���a��k-3'�z����~�ӟ���>���b:v�\:�G�n�z�{t�����f��Ż�f���\�͍�%�=�o�^�������|p��}�����7�>�o�9��m��������?|���-[��%���_?(9x�C&|G������X~��G=~�k�4��q�/�o9����0p�ܓ�r𩇜���;��}�1g{�������=�S�?��.�鏯���~�=���O,���G.��e?���+N��ȫ��Q??���9��s���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\����<��ӟ>���<s�_�x���������^<�3^��o��r��w������X��-�����o���a��޲���]���g���Go}��O>\�p�����$��W�x�+v|;i��v�A���b��$+���O��ϕM�i_J	{�?�d�3�9V�qi��=8�?b��}oJ�2<88�?pm�|�A+6i����4�����c߲$�UW����Q��5���3�%����e��@����o����	���u}��_�{������ہٓ��z�7^�34<�W��M��(��y�Q4~���	�Q�x��׳�
�Q�uo�w4�)_������������=�� ����3�	���1��ch[��������1�����;%}�y��H{)��P�8|�/G�C�9����c~B*���~-~9������8�$^6f��(SX���t�{opPk=�#?�w�J�u,M[��I2�,�;�ڒ�I;�lż��[�{.r#���F�m0!�OݚZ�O��c!zP�1��1�g�i`7m��A����Ջ3��įyJ-#w��	�x���a�i1ֱ�>˝8�A �!���2l�¦�]IS���Gq��k��m�')ᘉ144�d�2#ѹj�g\������I�$�d������I�3�)������V��Io18�ªF�.����S}H�K�y��o�9 �fH�#���a�_�-=z���;u�e��O?f��>��/�����ygo;�V���䶞�����i��Ɩ�YK�̩����{����y����Y������U���3xn��X���>�}j�Ȯ3�.��Xi�nk�m�\m��_T��_Ze���m��V2Wh��3�[��Z;Zzz����{�:Z�h���O����7��������nZgWߔ�=�6�9������cZw_w[W��{ʤ>���JoK���޾��=���;ۦ�Vwo�Z4Xʪ���9�K���7U[�ϙ?ܹx�~C�����׻GW�ݩ��g�j��i��ˤ����v�7k�ĉ��t���v�t��:�wBjS�s,��ur'�6ZQSYfLZ��&�f,�f��eJYf+S�uw�t���6��wZ�}Y�V�h�i��h��6��czo_+&u���O���5���}RG�g�Lj�I�A{tt�AD]��v��=��%���gW��{�ͭX���@(IԪ�8�E�3�-�$�i��fj�ƫ��fV�o�쩲ZVc���N���Xi�:�t�ʴI=m�3ڠ?��Y�t:�8���ul��so���v�7��?wwC��i-m��܎���Z<s�ҫ66�xz:�M��ySWKo��}=m�NoñT�u��w��/�0��6KþHE+S�wNj���Fvjo��S�^ē[z[�v�����tvu8� M�v�Nq���d����=ܿ{:!��=b���ޞj��9*�;�O	ae-�ˑ�5m���v-�kZ5��A�xժ���U�j\�TU��p>�?�'�y�ʈ�3�,�"���&��*����jF()����(�?�)�+�*��헱�`����if������Wߏ��폣#,R���Tl�s}?�j"���^���6j�BK%KK:[���3!,�X�#��Tq]�FhL�;t�<�2ص�0�B�1�T�*SȨ訲��;�U��4g�E� WX*/Q��Q�,�R�V���W�&��Q��]���L���t�����Q��>2Yr�E�@ڌ����h�N�c��d����SS�IH+��"}͠yZU2]r#w��dF�1C�R�V2�C�;5nG�%��P��:�D�l4��b#�e���؄�n!ӌ����Y��~�a"-#���N��L��RCH���L��t�	bK�;2iXfhaIYa�jk&�L�� �*s���-Պ˨�e8$zTPB��dF�\2Nrˬ��W�p��=Q�ϐ\a3Hڱ�
Ù�֌c�'0�`��X-�7X-�<����i5�S=�jLm.�GB	�rH˰5�u��J�*\�N�8b�0�e5�H��'OE���8t�tC+�b�P`�2�_G�@��K��h�(��@�Lׄ��'�a,ܶ��H�Y�K����O|tZB(,�Y����Y��5t)K��p,�|4��`�2�DX�ܱ�����9����`�$�J��s'��fp'4rYc�l��@P����AjI�X'��TX��1�f�`Ka�i�q�Daͬ�U�ۚ��:"#���+2xr���`2�G���VO��+�|�G�N���q�
�Bp�N��zlL���R(-�Xr�U����=Z��z�R+;��C��x(�+lj��� 6KDHN���RؐU�����#�o��?B\�� 6��`�h]i	3ѩ��ㇲ< 8T��p*]G�L��
����3tU�FZY	A��*�����*@*!)����3�5�!�#�8y���P���#���4��G�Q��a��m���@��4�O�b�Va��La4�j	�%�����sKR��"2���I3�	�	djA@a�z8bBZ����R5l#-#0��� ��=[M�� �O�������:� �}!��'U����H��	�K#SY��&AJ��BG8.V�r�����3@�)�E��n�H�g���#H������r)&N
mD��M��:B�#f�VaVP=�� 8�
,� X��zB���S�,I�Le�uոF�u��E�J�82,Ug�Ȋ4U#�~c3 +��%� ���R-�#С4-!�aN��W��lM"��w�u�~�	!g	�}!: ؊ʪ	�%ͬ'4�6|��3򪁓����΁�HR�z#�;9�0&D�j 2,��0#�'��0n�V
@2�ei�:
Gk�_Gg�wZ�0�0�=��
�����H����`�kI88x�;����TI��:x_B.�����U�.�"T^Aza�X�)�1r��ʔdqFV�+Ek袁����%�Ṋ`�@��$�P��dP"�iI�St$?�p�Q��a��`�8���"kD2��?	���SV���=�w�_��Ffjd:d���*�����:B1�&�H��]«�E�ˎ�H��ړ�E�p5h~1Q}G�S$q������!���ܪ�����B�p
���	/	к$�ǁ@	��q@�̳Ba���e,�qF>�.��!�Np.�X����9�T���I��������8���!� $mG@��b��8���j`�@�
pP�=��)+�ē��QPG%a	J@&,��(L��F�C`^[�R!#Ќ��Đ����`�1��3��-t�Ȓ�����.P��I��&CA>�pTI�u `:Npy���RE�-f�n����3$��"��rW$A�&-�jJ�gGNF��� P�N!Q�[�b�{kT.%E�y�������|�: "r�EsJua�*�����\�h�C��22Eq���\|E�d��*r8GFi�zd�by����T 02��4P <��a,� {՟?#�,.��Ud1CE*XŎМ���*!j�����LUt��XU�1.��~� �
(oɬ��K ]�K��H�R��=�T1J�B�)q�Q �F�{4�k�Qj +ǖ�Ǣ� -l��9������diY�)�F���3�`=�*ziV�3.�TQ%OQ~&U^�L���#+q��ڦ%o�H.�z�H��%�5*\*rzF�Ukx�	 �z��U8�`�Zr�H�r[���^ZVE.V6�����P�.=$���eu�'BO@.�:�		]GO�8�9�*�q犒?�����r�)*��e��'��APM�<��*|���֖G�ZJ8d���K9׬	�W��rr�
�X��^�x
NZ✰s�YVO�=	;�dp�]�ӦH_ѓ��B c
�M���x����D����ʰ��PM�Rg�%���Lu
	!.#�4��l�49�R@�#k��=���Gғk���G�7z��Q��8O�8eje^����}������i1�xA+�Pe�)X6��� lܧ�Q6�ٙBl��Cќ��g�L)U>� �*���@���2	�!�ecJ$YZ���SaY�T1B�
�rA��Q�R�F��+�Ѳ0���9�L��)��t�ʞJ�U��K�&���\�0�.0Q�3T����*~�*2T�}�����zO�oJ5*�P�`9�T%^3j2K	�T�2N�mI��.�Q%�8H6lH��@v�D�dkJ�eѓ������Ch��AO[�5�*�'$�(y�礷�4�)�6�Y�$��-�	E7h$�?Nn����5�|W�'���d%ޤhAb��@��p�F���	�l���'M�w�0����<��HL�x�(!���t(��t
cq	���SD��s�OHN������9hp��FGM�T����ܺ!�AHka %=�j���z�Y.[�|�{6�~f��ڗj�
�H/a̤�$\��en��IپѮ�! ��
As�2�OX�QퟜeJ�#���Sde���*����<�*דe��dd{�$-!0|�����ؚ�j�Y��d��WKuGX��tr���F�y��>��EX�9���K�U�r�h+d�q�j������x��e�:�!�zF\,���V�P��9u	֌��!mQAO)X6�>�'�iJz�}R�����@�	���@o�-�#�	�j�m��(�i���2㊚��@J���G �8�Jz�-�Ee)��'U�8�s"�K�$+�Y�jP;�R���H����%�6�*l���)k��<|YA�)E��-zRI�%�B0Տ�t*�S�X?bvʌ{�.�ӤU�C�T%=��a`��ӣ�|NI��,�Cq�4g���m������)�'�-%������yM�Z����$W ��gĜ�QO�!!U�:�	��=��s�|�XV��0uT&U��_R\�G���)�г�F�	�A���aD�L0唝C�/�秽	��<x��E$���D����j�� PL�,�E$�&J�D��0 My֌�"��E�h��,�*d����X.�;Iݜ��J��k�i�a70��\�T�6��>MY��	 <�D���!�/���e!�Є����=���{f�t���'l�c�.
��I��,$�G�P}O���hr+&�~Nn��n`����i��פP�f�b����jt}O*	�L�,^���ԓЛ%��I�� N ��P������ ����e�� �p�L�*t�����N\240����=�����z�����^�$6,7\�d����V���0�{�=V�g�YW��Ɉ��-���Y�y �K�U���dPt1D4�;`����DO�讑�HXmޝ��5{�������?wh��>&��x|��������G^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� V�Q(&�[   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �       ��    x       ASCII   Screenshot�M_  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>512</exif:PixelYDimension>
         <exif:PixelXDimension>960</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
ǃۥ  ��IDATx���#�q����]n`�(�K��%�
�,9��c����؟���e�z,[�
�dٖ�s�|"0o�����'l�������\wUu�d6��P��'��⻊����Z�ON���1�R���8T�Q�s�(���ͥ:_8��U���b���~HgC�<��L�^�0z�N��?+��������m1�N�6��|f��ǧO{6�鏢�Yʷ�|��W��{������Yw��W��[ǥ��8��-N2��>�#�ļE���h4Jф|�<x��� ~��,"�<�d��a3��#���*4]N���ĵP���$�H�˗,>�N'���W�U��p�>3Z�<=hmQ��흠��>1=���g�Zz�\? �_U�~kݭ�"�
�
:n��-A���D?T�z�
�րc�U�]���6]����U�e�.Ҙ�?0��~�f�����s���VX[[K�Js�������[�ӫ�F�_�$\��8�L��c�TNt0�VOv�a���|�b[�����|������/�ЅwٽӠ��|��>:Ҧ�\�1T�~P�bY9.'���ӡ%U������Z�����;�y�pKZ���\���<�w��;5�;/���+_/�.�g�_+�W���<Fu?�`k�N�x:�+A~W!�1T.X`���=\�2݉�_�X:�q�`L�c���r}�1u*yz,���i�f�gss3<��c�ܹs�Y�-M�g/\�z5��λ����p�捰��_�t|��4�P�� Հ�N2���Su��G1��c����Z�frK��EU@��=�)N�����3��νC^��F��$t7�! >;*M���iUO�������30�V����I�[��� /�ʻ��)/�Uˇܰ��ד0;�LZ�$��w��ቡ���h���1z�����>ht��e�[�=�9?�7a��݃_� 0�
l�o��b^��q��X2����˗�K/��~��p���4gx�P�۷wo�~��_���_����67Z |��	.���i�nai�@s3 N5'��8�)-���'+�h4N�߃}*����֝i�Y	�	���5qu�f��_�zH��L�&x�L���x�� )N�����A�� ��ڟV�>�<�P_[�����K��-�����oЋ5��_�>��  |�v�r������YQ�]��{H�[� ;�<�� ޽���駟�7�|3I�ڶz�|��m=B��a3�r���g�Mװ�766��1!߃Fq}~뭷��~����[oD ����f�a-���ͭ�1YK�Qc�;o9>g-�nܞC��d� ��v}x�5���{�����5��VR�ș��/���S����YY�:���e���4����>��о�������D�)��=��]��t=.˯��׍�]}��]��A �����Z{��g�ƍ� ���,�C��>����x7���KН��#u�Xwem���b�ʿx/,�s��q��G�w�}7���;��;E}�����Hrun~�wvv��ޝ�����ك�o��W?�$�5�P�s[�a{}3L���H���:
0���w�m��z�d2�@�`�wn�����"|� q�\��6�Q���yb����_fNi��$&�t%�5泚�\��W��JJ̓c-��{�t����?���%�>���ԧ��,��!.^���Oj�+	7�t�F]v�6�΂�R����Eui����	j��<�Hx���+����[�� ^u�q��s[�GN$�UZ������A���>�����M�x`X��ӤU�>���R�a�%��_!y�<o� #���{'� l�Uam�����h���!ovo� x��#�򗎀������724����������X����3J���Z�[h"���g�Y'� X���_j�U6��{G�s ���q�P	�� ��T��U4Q���åHvՁ{h�ܥ!��vq*�w���{�V�W䯣|]��޻�ƙ^;���4^J֓R}��Y��g�B�4�zh'�K<X�~������4tO�}~��q�i_?誳��]u��(���^z��
�,����R9�gi������gK y�K��{�Yg"wg�����d.�E����D	�U]��;��r����9��q�=+Vb���`�&���+���d�.g&�T_���g����I|)���De����d���\�_	��j����d�Ű {��Zl� ��m~	���l�F`;��*�O΅͍I�6捛a��t��ٔ=ވ��~��<������L��k����;��@����!��P��?z�F;�ׇt���u�~P�8��Kx��Pu��c�	���V�w��!
������R?�y�&P��_F^3k��#�>Z�Q�"�׎v���K�Ք�n�c%_�r#B�˽e.�~�����f~�A�8-)�ğ�������eTj���rH{��McW��K��$�x=(��]�t��a�{������x-�?�}�/��<�?���JϞ%�r�燮!6P����K���R:�n��������������m�X�U?}k�W�u=o��`ݻ~�zq߯�Vk糖��A��E]�� ���W�l�ݫ��Y��*�ҵH�� �!J���)�:"H��Gv~S�+;���5T6Z�,>ݮ<;��rC��|�f�� 'Gc&�����L���@�L�ur_�Ų7�VXh?��N&<�o}��g'Mo�O2�l����n�[��aZ�c�'	E���a��Ԝ��X�����=s��z�Ĵ� �Ӗz�����:	��XvѴ�>C���Zb,J`�-��ɧ�*8\�|���C%��KNX/�siL�	�}�]�-�> �E����կ�e�٧���Ծ������2��oɼ�
 ��ǧ�2�Z ����_]�Q}<�{��>����'�qi���6]�<�w���y~l�����N�|l:�����궾�*&|�]��T'�G�Nu��ǰ�4[�,��n�J롵�x��y)�Y��w��E�_�[���=�*�Y ��7!,�dJ��X}�g����J|�B��m[~�J�����K��h�vm>�@#�6���ߺ��и��0��`v���V�Y�Z����0�J��o�[7s@�Q�����)�*<hћK�m���B��ζl1;��t�А�ى�.�C�9�2b��>��:
�Z.�{�I�p��Z�&���a��8{�-/	A� �;Q���l_�g�X���*?J� `�;Cv~����U��*p)�H9�v()X�,����<���UL���-����u�T�[շ�&�mo�Yo_gMj�E� &�+�z��d�g��.�-��Q߸��i��B�Zy�ȅ]����??|�_��O�����=�u�(��} ~UZ�E�3�A���|�i�~�N�-�%re�M ����
��Vm���u�$ =��x����$�'0�lT����,��a�Ϊ<7\�bk1�r�-�V�_FVkۥ��sǥe���,�g�ZWa��U*�ݒޝ�U�7}�:q�4�$�'�>p=Ԕ��C$���<>��!��V�� ����oJ�Ew���|o�'^�0��þ��,��K�(uKn��t��}�:�?����s?��oyź-�O�N�=_��U�;R�.�W�W�U�|�Ix���������$��F�b/�+ ^E	����RV/�t�U�c�c^ã�}����2���|���c}�ħ}�?3��.Z����\6'=�'��&Ϻ�M��}�c ���t&���ws=E�^�����D����N8����x��zV���	n�| �^8����_H��:����&�}�i���kq몯�Z��
�ǥ�L<}4DYR�= R_V�U_���4�����G!�!=��P_��C��%Z�>Y0_�C�[P}p��E��,�\K�^�K�����Uz���t��=G�oY��_���O�q'�! �ӽZ֕��ܒy\E�C�
"�3wr�6ߌ-��3gm\J}<X�1���u�« 7v�m\��u[���	�\-<Q�V�6<�c��z�kas�N�dU�Aճp�p7��������:L�JD��[v�=��P�m�u�Hi���U�N&|�|Zց$2�wi����q�i�]���t��� d�9m���˙�j!��d��	��G��T� L�R�,��<�Œy~U���IP�E�� �:M��U��l@��'��9Z�����2��q4���]��p�׹�|<�Q�xj��.����z�*�<����g�C}����U��s%�/�����!��~�z�U�U�Q�#�(r��ݸq#\�z5��
��u�����~�����gM��w��Dw��IF��c��͛i��>א+e)��0,���?_.��$r��y����GR-�Mb-�ۃ�cU��fweY�g�g�d�iM"��Xas����gaRM㇀[!�>�,=����<�r$��Fs���`~��RZ$�4�&s&o�3|pU�_HZ}�>+��� �O(,�q�ɲ6YF��k,�R����k׮�� Ki���[�#[��X �Wά�" ^�@�k	6���_����W��zDp�ڊ{y��-��N�o�{uQ��rde^�mK�WRT˒�jh�kW��"[6��R��<��.���w�eW~��t_m�Ǐ�5;����"��`N�d�tEж��Wd就| ��J<Z>}~�~d�~�+YF���Z���+V���æ�<���i)�JT���EB?��C+[.��%ߏN�\��4D���ѽT��r���q����U�:�|d`a�9a(/%9� x��u�O�8
���O�$6k
>��Io2�� �l�1'sR�	GIV���NA��>ߪ�uh��Vurw^_��q�܈1����z�X��'!E������F؏�wo/�iS�e>k�6���</��=C��w�z�tL� ��_z���3�$w��k���w�x�ôJ�9��ㅩ.A����=�G���n���2�o_�k�Y�Ӡ�]UZR*ض�ڰһ}��
_6��˗�ŋ�{�^��t_��U5p[����F�5�&D!cgg��T}�Z��y��CY��k�-�I\�H��I�7eT�}�
���'���X���� O��-'��t�R�����^��ޑ�FW���B�4�했Rp �_�;]|�OzޤQ�S��tIA���C@�T��>�S�=s!�O{�zRTX}�G?��:JL��Wikڎ��oܧ��|y��^�O,x����r��D��c�q��4�~^
NRk�A��W����y��D�3%����)O�i�,c��M[�c�22ƴ�L<��:���HSc����=�7��.IG�6�g���q�]��n���ն�S7v	jC�-���7VK����م������?�0��4/���D:��?G�,���h�]ȧ k�6=�G�N�y��dh�ɿ��Ɏ��ր��1$�e�Uc�O^�>�:�$O�� ��i�������m�i:)?�N�YA��m��E͞\�=���s*�$$��9 �k}�ތ���$.\qT��(oEP��HX���(�~r�f8��:�1�a8�� k�g�2ε��1�=�s�q��H�G�c��������7�x#|��	Pud	ڥ�$����t�m�E�@{g2o�?m*�!����Ĭ��!T;y���u�/H�:��6Z�j���],=(�˶�/_��|B{�t�հ[�Ke�%��G���|�+_I�@���)ݣ @p5�������>^|��������GM}�=X���������I�F�ꩧ����/~��ʕ+��'�̀׶(�"�~����^���o�@�U�|_�P��������I4�x<*�Iڀ"���׿N�HR9h�r���_Nc�믾�j��������.	�Hٳ�,H� Ud�َ3����'m�����S�׭`j<͡\��I�����sK��f����]�T��_�� Z���^��ַR{��'������-i7���ٟ�Yz^G��'m���v��6�m	x꾵<��ݶ������,�'���/$ ?�s��/�}X������{m�⃾�H����}�k��7���L�����J X��6Wi� ��d�S&�Q�����i���K��8|!��/������������CyH[i���?o��vۏ��:w�:.��[�ft�>�Я}�4'VV8����>�Uʺ�����X��+RV![&� �N���(|���_��ϒ��� p	,�|m}��G�cUZ��~A��,�^JsY>�i���ݯ��#�
4D�-��%����t�C��5�-|�;�Pr��q����~�^��E$
��J6��ֹЙ����#p�{�����|��z=Y'���w}��a
~�QH�sD���F��&�\E �7�4>7ۍ	OHo��%ñ/��҄o�*��[�Y��o�[d; �o� ��\쁅��I*	�>Z��:���Y!.y�G=��z��[�TF�]W��o���W&,ȵy�c�ҡ�R@�Hp��oq�����λ4w��G�?ib�� ��+�\�B��
�r/o@���_~�s�KB�����3�{&�x |(w+���F�Q�з_y���o~3}�.���K9b(@�,^ +]�I�A^ƌ����I�V�� E�f��x�	 &? 
B7�l�e(E�PQ�e�O��U�L�]�PB:�J��������n�qiN�}����������T�3['uZk��Mwk��²���!'�'���vPtX���+WR?��� r�ԧ����5�+���`���m�)[V	��\�?�H��7���|3����)�,X}��m �W`�y�&}�5`i]�UVՓ���,��t�Cx�1 �WD�%Ɨ�[z���yW<X��˪L���dƯP���E�ط���Y�*t߳�u����3���X�����~�Xx�'�������S��4.���P^��+/�߲���K)�Ө�ߟ5�S �_��c��%?� X��P�6$�㌇���Y��J)/�j�o�����A�k�<gd2���L��(����O���wTf!�����
�.����q����r���n�O��d-��( ��F��m��au5T�3��]�!�I;�gLp�+rV���j���oΉ
ᨦ�n�]Xd~����?��!>����� �RK��|'�{� ���@�q�%�z�o���x�tX�´��u!$|��?%��R&ͦ/K��`�}���Z@d��5�zhy*��ǥ���>
��!aW���E�DX���O�#���� �L.]�Jl�& k*��"�x&扒��<X�l��
� �����HV9,�X�x ���pN^�����SN��0�w���/@C�k҆�w�}7\�v=$����9����$�"|�ՇPB�k����T�C}U��;����q�Hm�t ~�_�>(�� ����T� `x��4kW?��S{�tOʉ`�c+��j�Ro��SYJvQ}��P��>V�3�}������c�O>�n��8�/�<,��#EƄ�W�x��J+x�?ұs�z�M��C�P� ͭ�O�ؼ=pU?�s'颸�?��{A�Q��ۄ>��	H���'�=ڍ��7�"|Ka�~C�<o�w�L�q�/��^��S�ȸ�l�޽[���q�y�@���%��2/��������-�iX>�<b� oɒo��R
��B��[}yڶ�s�_�|�C���Qw�W�!K}�t��j��i��k�;ݖ'x�\�l|w��7�j���v�=rR�T�{�Y�^o, ��c�0
��aInv0�� ���m,���8Q��zC�Ո���X�pn{��r�U�J>��m�T	z5Y�X��G�����ݙF!��nޞ��}
�s�&C4���]�6 ��oYr%�'��E�sj�%��Dأ��@�� Wľ�f� 4��g�=�>=-($`x�tq��i�U��L[&+T���Ez9 !�7���,| |r]�>0��V��;`H��P�`J=S�0�ǖ�
Q�u[iv	%˯� ���xF��h/�-e�9@��R�����(�uM�|��kڟv~����:>��t�>����*+��#��E>��r�������^K.���� ��m�5�4 �ԉ�zEM��r���~���P ��C]� ���E���/�DVC���/^­���3n�t�~c��o9��.���C�~�L��\�̌�J�G��{!=�#}��G���l�[��v��<�4��+Bc�׍���e����ӆv/��7�����æ��}���M��◲����|����e=����n��>m6j�@��Ϩ���ui>�B�ʱ��պV{e��ԯ����r�*�ER4���"omm�J˻��T/�3x�:!A��Oj�,�������K�ui~� vxmY,0�T���w�Ǧc�W�'��B|�ս~{O�*���M=�[�Cv��Z�����C���j��mz�V�sd>�-w�F;���;KF��5Q���ſ�yPPg&�[aa(򹹎!.� �:�N�� mr��A�I4��f���1�D}f����i�=� "90V���m4�#,Nq����Fu\|#8�~x3�eO����U
2�+�I�|V��Rm]���G��W��KUڝ&M��[��x��p_��W��p�p Ṵ�N�'��G?�Q�?�ߤg]����u�I��_��_�� PN�X�x^�5�
�"+���� ����/�2�;lJ����W�j�	�UP�KV�8/��=|����r�g?�Yڏ�}kV�n'���r�F��+շB!��n�K�}����G��
��ީ��~k��q��F Ex}��˩�P@�7�Pq�%[�<�#��' ��E����k꟔�2#��mK�Ҟ Tܘ�䵸O��=T PA^{���O��O��ڀ:��Z>��bY�e~ȏ�Rn�%`�	�]J&��\Ե7W��� P 1��@"]��8��S�♼Hߎk~ÿ�+�(�
c�|H����ɇ��7��G T�RQUIW�H��〴�G�ȩ��󋢳�*��/+��SҁOx�G��y!-rq!ݹ�>����]�}�w �|ķ��\����Ǆ 3��
�Fy�[|�5��@@N{��ԝڃ{�'ρ�|nn��{~��UX�+��������ǁ�7�)c��	���W�_ xU��$3�,)����Z@����vYյG>�)���[�B�+�炽fA�W�����j��ѯ%�i�R?��v�k���ȳ.��{�!_��Lp�<K������]1IF�Qg��P�C�|]ƃ.*)TV-�C�7��0�����jK�oi����x�c��~�o�8�b=u,~�S � ���QFə9.R�D�wx�V�ɫ9.���<�<^&��	'�	;p�=�����{��Z�{��n��Řg��f L���&k�I�<_��>����%
��8i=�=�3,Ur�fo�F�g����],����5yOhf�⎀���#� <� �V'�1Yb%d�R� �~+	�,ܗ@�V-�vA���ٗ�0�� �*�k߲]lĿ�R:�X�VP�B��A$� ¾S\fD@�.�yR6��> 	� ̳n�ǩ�� zꇿ)��o�Ic%B��IT��3y��F����f+�h Z���gd!�A�dŤ]I_��ߺ+z����(;�\�z8x���[>�!�|�~�e�����C:vo;��(2~��~J{Q��� ��X>ڗ:���On]��XՖ׮_K=�?mtc���/����������ܗ�ʺ�Rf�Y`�� ^I�G  җ5[��e�:m��Cc�2�?�×x���'�e�����C[��RvZ��
�iJA#�t�@s�~@�GI� hv�?Pn��j�>C9)���
�[�� �KI�D��]����@�x�7��=����~<�B�#��xOn�(c(#m�A]�kD��m��i3WP_|�k��%ڣiwʯ(�/o��أ�IO�C9��_<C?�2�&���C��[�8���\�r%�	������}R�0��@��hI��Z�EA � �o���||
�O�x�y���0+h��]�`�J��y.'�ȟ/)?��Y�=�)�A���,�ڿM�%�%�{%}I����c:�C��ҽI^!��V}��2i0�E��e4�k�o�� �-��J���$/�E��a��������6���&.L$+�8f�w��c�`���g�n�B6
��q��r1K����қ�Gr::�V�,��ɕz��ѭ��K�"?��ۺ���J�8L���y��2I�kq���s;��}{'-�|�م4	Y����Z �j1�����B�Q ���I(ױ�~�{�kݕ�l�䶊 ����M�ɥ��� `!��A����H!�K_�R��P�4������ UG�(_	�r	��^GdHx��B�=�\`~�<��T>� ����IhU�,��zN�Ԩ#�<���}X)�7 �K���O�@�/��5FV:�&��,��+.�\iK~�?yX����([V4�ٛm-�^�P�:?�;�8�� �� �
�����B�O���3ԝ���}�w�?>�a�O�,��3~˲I��]��?�I�N?��_��n���έ�hEXx�� ��ژ��7����7�=� �I��|蓌1�Dܣ�H�q@�xO�G��EٹGic[�n��-���?���/�՚�i���M�YVTꞺ����{�A�@?�]ȇ1%�_�?����$~�O[ǤIy�4���h¼'w}�Ń����\����칂b�rqO�ҧ��1J|�������'̐� e;h�t��^�e��d,2��Q[��}�S�-�[�Q���pT 6EZ�̴�r�k�KeMd�hS��L�ﭦ�(y��'쪙��\ؕ[7��|�� ��P�'<�����<�-���𨠯���f�%�A۠8�_<M������+�nXg�'��qڏ�~�v�Yk��gN)h����<��@S�KQ��	m���<<(W�~-n�E#P�9D�i������A%@o����n�i��6.��Q��!`�	���[��Q��ݥ���e�����UE�C�?ȷ�2�H�hq���\���m��ǥ���������=����D{��Oi��z� ���q6�$&��a���0�x-��ǻ*���d��4�Zܥ9Y)�y�.#��oHu�)�ܵ�/�&z~=<z����b:��YU8�@8T�q�Bc|���sa/�*�>���}�:OTnb��FC�i�p|���'z-�c4�y�s����YUR�<e��6] e� B�,B���%�ĸn!T �q���kr����\YI|��Ւ�*��m�����Q.z��l!��>n\������7'wR{��.K3�#44x���q ֥Ng�R��|#@�)@^n�r�%}�"]}�� ��y�)/d9&?�B�DP�_"�+������#�PG ��Zˊ�d�y�Rw�Ӱ_t環)��Gm��O���hb�O?�tx�qod�J���a��~S~���J�պ9R~��Q�\�x�b@
�.�~+����i#rMg¢�tR^�D��_�{�2�����v�b�h��y��	mŻ�-�0���Љ:��:^�H�@��'�I���Yꐱ
�L����]�%_�5uy�=ל��=Yw/_���2��l�d�>㖣� �
�F��/�W�4vc=P�:�6)o67R� XQ/�%7g�#�VSnU"��M���\�A>�cY�C`�y�jS���8Iq��z�Soʏg�h;)�&���(u�|@�Q��q��{�1�B���XTv);�+�C[RǤ������R�6 ]�&���Ns�u��V?{���bP��\�9����苾}�M4<����~k.�{8��/(
��V^}��`cԡ��l���@c��a�tZE�*­�=V�CxZƇ���5�*c��
�d)k�-GU�gv^�Z8��ӻ������C������ՃD+��]��J]�.CH㮝Sΰ_��v g��b�������F�r3����6��f\�'X������z�:�H����~���݃ð��u���dE��(��@4!~����"v��A:p)Ez��wF"Qo��n^�� _o��q��*@6�oD~�b�>�������DJ���,�T|�mV�.�����E�Te�M�y���_W�Ka��i� ��do�N�rSF��M�#e`�;� tL�pRL�X:p�xaPV(�f���<K�S�� � b����'_��r)��uҥ^�� XBy O�}�5V�C�X�x�g�o���;��A�x��)�%�G퇳�~��a�"_�2�K	)u�@L?�9:�^��|��z��%�p-e�����?j��,��|�.�?��j�^B�����3�K=V(����C��}Yۨ�#�WxF�ʨ ��g���!e��ְn�C��Uaq���rѷ��is�.e�ǂFIؖ����4�#훎e�Nȋt &���/S���+���_�������w��_�{�0ɇ4�O��G+�W���Us�N����@��Z�s���w�����_x���y;���w _� c�6�����S��g����c�~����FP�:�/бE�D�R����*.,��՞�L��@X�֒'�cȃ��M��|H�v�������3ڄ~M^̳� ZgM�>�ɋ^��K���2�S���w y�ԛ"?{0%eϨ�(�=ZJ*m��y)�J Qml=�P�_��|�]�����i��P는���)����F����u�B�4ֵ�"��?r���qO������S���g��@l���T�}�xϟWy����u��Je�Ͽ_z�$$��)��Gt�RlZ��>���Z~�<�ķ���Rz^	�W�C���`(�餖�������Y�Ϛ��WR�u)�:����j��̇�PoheQ7<��R �:~�@{H$惰��b����in����;����a��]�;�+�r����ڎ��$R�BFAq}�7���9_� �8s�oU�h����x���k O���i�qa�u�F��c�Cs��Z�����Go�H�I���J�K���9 ����j��-_�b��8��ל���ͻ\"`�]x6?FD�U�N�&�*V��~<�������}&R T��
��󼋰�`� ��G�<��<��ԅ�7��V`�K�΁�W�
��&��d_��LٴwӞ#�TW��ZVC(�m���ٴ��z^o,��!�C�H��{q�G*C�N�Q�����J���(8_Ku�UP�_I�2�>�#�y�=���HC���e}��;�J�����������6�D=�O�
 �U��T���3i��׵A�,IIa���G;F��-A�zuX `�Ժ�+-�`Y9�e����r�
h��d$�-.��� 0�>r�^}�2�(�H8 H��z�y�����JHZ
�E> ���9���#�2P�����qO�ѯ�3�^J����B��0#}���c��9 "�F�bJ�x�y�b�i��@A�l�y���� 5է<]�/+"|iϮ�xQ��?ˏ{; ���0P�P?�)�р`ޅw�˅_x�9�m@r���������@��
���E����<��e%k���8�M�Ѷ��'�	�EY��N ��-�=�H�S�8y�g�ğUjɻ���G^s��֒�N[�- ������J�D�E�4u]�pI��GmZF����׷q����q�ϣ/=�;�\"5wM�vjo�G��kB U��	ZOK�47�5��-�i�`��P�%�@�n��,�$����|�5Ov��R�)g�g����߫�� \5��pV!���X�p�N�M�� Ճ�q����#�8��Vr�$R�x2�GY��,8���Wk�5��%λ}*|��Ǣp})�?�~�}�f�WW�(t��W'��$��q��e4��6{�nD�歃d%��
�zr{��y;	߸�r��IpA�D�A C�І�d�3'�w���}M�}\ų�3���Ӑ�������"L �a�@`�� `</ (�� �\/���B>r��7麗����Ә��Q8���g?���*Kl-�7�VY�a��?�q�aa�!��k߶�a���-i><ϻ�b<*/��侀�y�.Fh
ͤ�����7u�3Tu^��,�/�qM.�Xv$�!���
�����>�/���p���R�k��(�o+<[+Q���C������G�
|F�����+����(�\��u;�|
�£���{�e��ZA�*3����G|ـ;}{$m]Z�"�Z��Ϳq�g|����{�c����J>��_���s %YN�(]_[o]�e�J��S��v�����4���k.��3���o����2��mF��f5�����j��3�eŤ���
L��y��h�><���	B(���gP)ڹ��X�t�~/ԩ�����8��^���z:���W��R���R"R�K�m��w�C��+�=妎���?�'<ۇyU�)�Jԟ�zS^Ə�Ǔ�׾��4gG�{ޟ�>{6�=ݎ��������b�OT>)EQ,P�ӥK���۳w)�R^YZ� ��ߒ�fO�p �A��l����W��w���m^��=����]�xO�%k�}f�u���ur!���{�N�On��z~�����@PW��_��'����+��uX�XyHw������Ί�r�t����O}���8�,�#�)��}|����u{=�U-\M?�g;� gov�����^�͞޴�wD��:�m����8�Momm���kam�R�<����������Q���"Cc!��5lmgK0^b��߃)֘�p��p��4|z-
P�82�f�ً@��"W	�mmr��d�˂R��ǒ�'�
 ��䳥��+i#L���6j�UU�����^�$u������$wO�Y�~,�s�<"���ŉSGs�D[7���5�V�-~,X�Ĥq3���w�FP��6�BE�C���<T�^r�~t��CJ(� z����Y��N�.r�J�Rm�U�>�	����6-S�^�[�oK� SWRL(xuhR0!��=	��O��6�ՖRX��
���[�Ɛ,����Ҥ�b�����v���0���r�]TdEI��B���u�ߍ�C
@&yP�<��Rf����G⣉@����V⾬t�X���ó���c� �Pc����s�zAy�u�	����<�j������<���(��Þ�l�E��>�ɥ��(8K������	^��}|Y[�u�;r�W�2� �����u#K1i�eYQ�i��>���oVB%����l����������y�:���'�LGL�e�m4�� ��W@�R��# ��S��������-0�i����O���O]e�A��k��]s4�k����lU���W+t-��:[�3J\���0,���I�iGx`���t�_�^R�x�n�]�f�՚Qʫ���:sZ����w�S_۟Y�/�������_�o?v���9����q��R��{��@��5�9�6VK`D�q��	��NXq���,�xo}#<u����O>�R�M«���}���λ����Z�w}}-�?�Ν�lą!k'���xk�RO��S�<ӻ����>�z#L�G�q�0�Ӑ4뀰����tD�N@�>��#d>��g��F3���A>�㝢��wܸOn6�m��u:���O>��������G�V�J����X�pa����u\���|�f���#y�!�b��o;	���?n*�L����>�!l��NH�| 6ʧ4��$6i+��)7A����l�W�ldʢg�u͂b��~5�l,K��_�]�*J9 ��s��Ӷ�}.��8����Qʥ}�JW��I}Z NmA�*Ye�Yp��#��ݣg�>@4�xQ@/> =�\��^A�#.��ĸ ����d�~�#���QO=�T��Z�)eA+hcA��Z��o6lD[���r<�g�\�=���)���o�����|Ξ],���̑���O�]B9m�����}�z%$/����a������?�Wc@��(жnlY��T&��C���u������@�:�1��� }RnI� ��g��5�xcQUtn;�ԓG���S;؈�60`�����s���k���.^���f=��������Z�=Ƭ�:nJ��4g��j�쓟���6���(~��$���l�y�̹�z�\^)e�I}���Y�6�{��/%0f�;���O�i�+]��oǴ��*���b�������n�w����e㼯����4���,�?D�q���PIizDq����S(��V������BY��c��?� �b���:z�v�KS5�D���%#=������O�g>w%\��D�qk�}�jx����{�A�Gao�z��q����v��}n3��n�ߏ<�A�#Q�:vvq}�`+
X��:.��A�A�8��
i����pc:��.��ᒵ}n�=�Bh�e����O�k7&�h�z� %׾ �f:[a�}j1 J����+�#��壣 tP�G��t�g{�j��@��L ��I�{%�'m�������F^x>GXŪ��#�R���CG��Q	UJ -	۪#x�Y�lQ>�'�Y)�\�K�X���Y��"ܒ�1e�0i�F���)����(*>�(�������B@� /�7��q�
R2О���-����F��Կ�ᴷ>�h�b#=������dy��I���^ڋ�{)�0����*>t���|ُ��Ϊ&}��z���Ƌ� ܾuۜ!�)M���~�����Ⱥn][���6Z�w'׻zަ+@./=kӰ�*��>���r3$]�s��R𮭤�r�~�5�jǀƳ��Y�M��U�����a�+�� ��\�8?r��d���mZz�ǥL x�n:h�.S����z��̕�2y�����@�X`�VyFiN�{���k�C0���Y�|�EױU��ҋ�D��3��ev,���m	*��?�btYw;�wU��>2�+ɹRk�JK}ƻb/�W�x�Iïa]�ܕ�2��x�J��gK�K���ٿu��7��=��>��zXs�����0�z�Ҫ�׮�'�cd�Q�z��xu[��P���<�R��jaڬ�^�i`�DH�`�_
�>�B�/��_�ֻ�����7�
�n^���`�v�Q �Ջ��f\�o'`;�[���5�
g�;JG3͒��(s���,�N����'��׮�{�E����Ih'
&�IxC��֙S�k�]�8�A��W_K&���w�}'	���0X &��P�b��0P�N�cVd�@�EC���P�ˢ�!�(% ۂ��н�h�?�y(�3ϓ&� &eH���f������,��*O�V���`��B:�W�L�J�Q!�׹��%�T�������R .qґrK�e����H��H��ԇ��_E����] 6rS�����v��BT��-�T$�4)�-u L�� u��*���~c��>^@2��R_�GM]S^�Β>ߊ�HQ�ʲ��k#�r��q$��W�Z�a �ʥ��Y�L#;qN���,���ZսuU?�]5��n��qמok����~�ׁ�JغXЄ�E@۾�����Z~ӟ_����/i���"��L����������*4�|��ߊ���k��W�Q��r�] ��o�x��	�u>�G��NR���r�KѸm�{t��7Tf�����c����\XT����%z/kȺ����MRF�c�wt6�������Қm��� Vv~󊝒h����6�x�.PJIbݾ����G�׎Y+����+fJB]�P����$T�}�iI ]<��C�)�Q��i �������P��}���Z�J�� w�[�%:~�D�=�����Y��P ��J���3C��zsT���9o�<�LA՗F�?T��z҂�#�.���ڵ�ŐL�u��fn8�詧�	/|���d�������W_+��Ȏ��X�QX�f@}X����:h�q�kq�g�s���Dp]�����4]� yՖ�+�t �\�`��R���TdU��e5�|��d_���݀��ͬ��� ����۩$�����O�&aS���0k�G��&p&WT���+�Lʹ���X�� ��"�Ճ�yJ(��<�<'K+?+�(_���"��o�#�B�Й��!��:�o�r���k����<V���X�Y>_Wm.wQ)H�G>��oC�f�tIK�R	�C{)��n��n��uiL]��Z+� �����I߂3�Oڈq  �S�:>L��|�*��r�J����\@��Ѧ�������+���C����:��|�u%��Z+XwYt�����c��u>/
��#�\�Y�ڿ������g�]�m�*���i].N���a׻�˭8��3��dS`7��Z'��<7lh��B��aqQ�e�J�4�Y�uF���9�:�(��Iˎޥ���qE@g-`]�1j(@tl})��n��S~>��b�PP,�HgA�--��`]�H����S#��{���j?�JAu�Y/���F�c�|t|��Y�qWV>6
����ٲqd���T'rL�@�/��v���[��)�<8^I����ީ
s��r�S?�-[�	���և��*�\�^W-]���*�/���<���P{�����:)�-���o�صt��Dg�>+�z�B���ԟ�&������������Z��P���R�B=�ىΞmV)A��.��Lu[ѣ[�Y�#�[������ҋ_{q���_�"��O" ���V�I�I�)�0}��Sk���\\�g����D<�U����qߪ�K�I��P�#��#���'?In��s�:�}xeᇬP9*re%��1�z��\���2Y�q�P�!��R�!�ɽ��b^�B����@��G�ڙ�;*l�UO.��C= �e��̓`zp�>�>V��zW�"l#�B�p��:�|$pC<C�Vk-������coHa^�]�L�ؙ��5���3�q��BN���&m�{R8��ԓ?��։���%ɂ�Ћ��o�/1�QY�s) ������ �|����.u��z�R|��'�� ��V��T�9�R,�8g�~l�ض��R��X�)���20��z�/������~3�m[!۶��Զ<5iYk�u������1�s[�kvA�.Җ7�7c����9Z��Ӿ���+��)7�R����^Q�ħz�
�& #E����ƍ�gun�<T����v3�`e�q���П�B��N9��5���γ�׹���D�-(���ˌ�0�"m���ҥ�)@�\�����t|P����&uOz��5���i����9��%c@��p�o(���<L�������R����G��@#	�FicǓMxD���/.�{�{@շt����Ӻ��%��Pa��u\*)���v{�ѣ�"p�|%����Wx^���8v�!�[\����SI�f�WH�j/Ջ��d=v����Kr�B}��д��$v��{����ï��]5����E���M�q��#Z6�{}J���QU廋&R6��Ѳh��_�6�/�_�E���.�d�^z����>��4Y/_{����믦��5�ㅹ)���z{fm��c�eR��3�}���c�8r����dɜqm�Y�@�rۆ��otX�;,�,��;��,�Ǉ���I���ÅIxkk;}䞬�S��!��
 a�<h��@�"M	��3���6��HǠH�Up	8�#�l���<���
a�^�ܥٗ�Ż|j�)�τ���y���:�D{���!�k��:G�P�������_��I?�Eוּ�jG���>Ҿnw�����f���
@� ʻX�li��6 㗿�Ujܤ	6E>(�LI3���i p���12'Ck[Bi�S]� G��%��x�>fޣ_f�G���bO��k�¦�K��kg�E����L�xk���ϭ˨U����|i\�g��(-h#�Y��h�G� ���q(�j��Rޖ�Ң�]5�5.U&��>&e��'e���g�e�y�*�le��1(�7���4?0�$�3�~ļ���藊p~�9��`O�,�ʗ�����NO�c��Gjӑ����Cs�Z1o�cO<yP�(luV���>�<����^(3�x��M���~��_�?�\�	�xi��
�W��{%˰����ߎm�g�y��ԅ�(�������
 {���sK��uO]e�@��sa����Y̧+�%Y���ɻ>�-Gvl��]`���5?Z����-��E��.pZzήh��|��J ��ﲶ�{�D}k��<Ϛ��l��pϔ�V��ۯ�v���ǽF���g����@������Q�6��*����=Q�Aŀ�a�c�@���-uQ����~.�_P��/~����(,|�ɧ�p�TXU7�Y�L`�8[G����(x=z��$��c�&U�^�o��'y��⽽��ٹ;��&�$ni��@��]�ٝ�wђ%��?�i�r�J�YT���0,�+�F�+�B�V���½����V:�xcs#��f�$��9��f��  ����c����dj��!�gy���0��/})	�X¨'�G8��c��ז�ԕ��j�'@�@:�!x*0��T�jʷ,_�O9$h�7�K��@�вi�Cҥ��Y�A�~�+�Q'�+��Zܷ�b�	Sw�,�оG�tH.�H���T7��O��j�N�eTQ�� �<G]�������8ξ��o'�y(�'u����i����[�:{������PY)X�������|�U�@�,���� !�G?�Q*;�,��{:ig�����&TI�� =g�&�k�����/Ph�K�_���+ �ⁿe��3��XǱ~6H+���q��cQVX 
i�����2/#ێ�c�
�k�1Y��N_U@=Ƶu�Թ��yc�
����W�W	�������JY~�ȯ�bH��z@a��qBߎ}�ʋWR_�ٹ;����F駹���2�/�@��@��[y�صI�r{/���/��+Q�����g���xDP.�:�A�:�H}�*E,��/�vN�����,���o}+)'�x�����i됏-�,|�h��J������.�t\*�v�Q�^^0.;�Un���N����kI��)�+~��j]�R����}�G�|ڭRv}R��\ik�d(�-a�Է�?]m�L!S�}�Ļ-��˔Q�.��v�<~4��I~Ϳ�d��zYRJ�ER
[��i�=C����� d X	�M4˅K�O'�oS)�B�;3B���=�@0�X��^{=��ƛagw/.����6߷�'�Ix��#m�#cΟ爆�IH`�k�k,�yO�9_6ʈr��A����3"�� �ܾ��X�_��[�IR�(do�}����3@@�dr�-6J��SwTZ�<p.�;�����SO��8nʵ�M���ZM8����.|�aLn��	 3�
�0�y�=#����h���C�IZ{�d�H��������J�?5y�7���G}k���R �𫽴rIV4g�xu�WC��H���ڹm|,�PDS��]�0����i�0�ߴ��g�y ���J��)�����c*փ�*�P/eG>��	WS����.�����,Y!�f*7rD�HB���h:�� �Oڒ<q��[�$��}�� 
 Z���"O~k��Lx�7��u�>M~���w���8e�����3�xO�?�����Ku/�q�.��&�S.k%�&@@���Q=M����;��s�gM�+ҐeM�@�)�(��M-sEcݞ�L�]T��^��;��B�o�e��<#�����붎W|j/;e���o��e�T?b�4|�@d^P%����K��<"��b��ʥH�RʳB�\�����:���.��Cj�x/��8�9��/~1�CY���׮k����<�	�.�Q��WJE�"O�]�߭0�s��v�����F���N0Pz%����\�8N�y�KiY��K ���%-���[��ci��Ζ߻�z*�U+d��Si]���|l>���_X٢o��i�բ���a��X��C �k������2@Y��n�7]
	�L�yD2��V�`�'���D�ښt����=�>[-�!:�U:'����d�u�a�0������D������阡�^���~��ߦ����~�q�V���*�<�8c��أ�������sX7աy����>�0�Y�����t��N-�����#?
��~�l
�K�4YYp��G��'a�g?�i��6��\��dU����i����uja0m�������/s���Lc�F�@�<�5 �ʢ.�"#�3�
��Ҋ�,!�o	�Xd�7�e3)��#E����rP��T�h��"\�X =Ey�b�=���e���$�Œ�ɗ�B8��3t��(��-�Lj[�a�Ad�R��_��������H�$@D�TP�����Xkń�9��<#WP�hb-o�y�ł����CZ�HY�}Y�W �<e������4�ƾ�*q&v���y/�/E�T�,��������GxF�Wg���ϴ'�9��]�@��.u�=@���� �����	dQ�<O;I�3�m	�� |�,i��?�C�U�@��Q����H��0��# 5���Hq�����4Q>@�jO��H��	ս�"�2�e�M�og7Yn)��((�ܟ�LU^�ZǤ���2g1?��<(+iI�!e_�{�oXΥPa.�x��K9�M��3_'��A�������=�e��N��M��XǸ����?ܮ��_�5��;o��}?܎kJ(�x��x������/��f��,ڿ������n�r�����A��Xk��f}Q=��D��_�UN���?H!�~d=��:�5�����D����;C�̕k����+ӽ�������n�a^�
��0�p2�4
W��б��o��%k�0٥ظ[���!��+PJ X'0?��:FU�C��=�;G�pC=�#Ϥ�?��͍laLB��GҢ�֛o��_{=\�v#��'��{w3t���~ Xr��C�'ι=<84�7�a�]�����4�#-�,��8�"R��rs#l^��������:9���f�#  �&7h��v��S��W���	�
$-�΋8��f@�E}�����W�'m=���Oe�E�HG�D���oYO���o�]�[{���i#��]Y�$TK��p��:#VQK����Ϛ�|�畯u��Ed�G2�Z���	��bB���ӥԄ*�z���s����FN�z4Ey��UϺ څ��Կ��R �׺��,�!L��@�ƭ���2i�]���X�Ir��u}�Fڳo�ӻ		���&t�QF�K�B��#�J�:�Y���c�H[�Q��Q�R(�F�G� �#�W���,�����ڌvXҘT�6�%J7�e�d�g�al**0�(%��$��Ã��ʡ�j��S�������n�蓅[��
����87����pO���e��� �*�b �m�oI)F_b~�\���6&�~�<{�� �����i\Q�|�Ma���gU�}�V���IZӪ�<Ea�����E���Ǳ�>
��>��{�H�:F�1���y�B��_KԯjQ����JC¢�</E�]�T��cP��U�Y��m��bShζs��Zi$E٦-�ϒ��2Py�ԺqvTu��?����9�K6L�ӳ��E�֑�>�gG�]�`}*���]���r�On(��ū�[����H��f�q�9B=R�A��f˳l�죔F�t��q��, `��`�`��<yx�{ ���i�7���w��ҳ�I��m��>XW�L���[���O?�L�u�V���çGװB�#P�H�xom}�R��=L�G�gD����f+�l4pyf��(�;^��;-�⚿'�K�����,\��bZ8�p���s�������&I��1C\��n�
-�AH�-�5B��{�׍+���S��F��9�����]�3:�R�gN,�p���	��Ig��,��79��A����Z��³�z�B�Br����	�%`"dq��,
,\�ϑ�Gh�\rOԞbݚo�W�X��ܕ�kY����}v����Ĩ��n��XeB�������r.k�ʫ�� H��3���v�@� �����F�\�~Aձ.�O@Y�H1"�ؐ�al���Β� O߇,��7�����嶞,x�^<W������7��4�q;mޱ�Ӵ���W�>�~L��>[�N}�j�!�k�m0��H�v|J�P�<)ФdS��I[/��i��ʫ������֊����͂���s��J�T?̫�Y;k����ʍY�]m,���q�+�n 2�u@l��oD ��al��8Ni�F�:I����^�+(��~�-�?|��8�0O۽�⣋���mc"HAj�9B�ׯ>��P�*�K)R4��^��8,)G�����nw7�]��Nu^�Rݥ����׽M���m�p�(��=���}�N�GC��d(��"�؂P�]������3�^hG)+lz%��y�Jמ�`���?�inb 7!_��_�Z���I��v>���R>^��E]<�
��z��t佪9b��R��^ ���/S�t)�������v[m�R��"ڶA��y��	C��I�p�i�,3���5D�y��{߮!Ch  v��Ց��T�JYE ��J.r�$A魷�l`�H�UD�nn��}�x4?��Si��4}�i\Z�UZ�'y�/��$F#Ŏ��Ѫ�6�'��ētcgg7�;{�m����&[Z��}y��-O�����b-uTu���"ZM�(̅C�9g��������Cʾ���쇅_����k�h?� rp��������R/(�F����G�H�eu���ON��!	u�J���þ癉�,Wi�����w�����5+ wiB����[����d�	��1�`�n�:Qy,`e�  a���-�ј�YZ�l�z+q��,p��>�4��U��|��pڼ��?�Ѿ;W����\j'pJ� ���?e�'��4���OR�X!�֓��g�MG}��i�s�-��dܑ��ֳʯ�k������+
�8�} .T�xV�
D��0������ڲ��@�I	��3RlxŊWnA�8�؟�W�����9Y�G^1���my���V� o��� �֭��5@���Z�RT'�1K@$���G�}��Ó�n֍b������ �g+X��yt~�.�Y�lP+Ճ�Ԯ6�oK�j]=���k�����QS���~���i�
=����1k=���m?^6��9L���Ǝ��v���}����<�t�{���;U���z9nk 5}n� e�[���s>�`�k� ׏{_g�k~��u�>���}_�}�X��E�T>�Cϕ+WR���|��I��9��3=��*Ճ_=}<.�����A�2�{���x()5 ;~���_R �d:^���}܎�.c�2��$T�����_����o��ߪ�t�}4 ��P;8g�DWu�9�����v�/^ �Ux�ͷ�o����5��5(k���w�k���>���������	0�`GYF�_<r��dn|��ﬞ�G�!�d�$!i#��{�֍4	��yp0���G�%[$�|�����P��W�l7KƴPDU&�1����FY|pپ~�F��nG �~i�lk_ `Qt��
.�� �E�Ac%�c�E�I����\i�/�Sp�=i)2��S�v�� �z����Ϭ�#vd����sr�E�&X���}Ȳ�@ʓ��9	J�ɯ�k�x+�Yˑ�8K��h�����`�*Y���g�]�GIP�J
	d���7��?���$���-�޳{�O�
�%�U"/P��xk�U�@RJ�=\���jW���,bJ�.Xj
~��F͑R�Y�m�[���.�-pU�؀B�����mA��G�)�b��s�O��A L���x�}˂8��a]��3^AR"�,ň޷m���q0O������_o�<yA5�dN\h�3#-~y]N�)ϨqM�F)�d�V���6�wj?x�d(ŵ�vn��t
��:ט^P��z�}��v>��1�[`�F��"z�v�Rv��`r��kǫx����%�x��N�G�M����G����{t�Mu`��3�c�uc!h��@�����t%I�u�c%�Jh�VNQ�`Q�ʗ9��L���p��Ұ놭W{ͻ�۾k�ڦ�缲E.�2 _~���o��x�?�4J�o_9W�]u��t)|�O��i�i�*��km��1
���Hq����n�,[CN����l^�T��3-��
W����N`�rM,�k���G�@npk�� �d\w�x�ɴ���nni�IQ�q�^�G#!\��w��c�Z嶓��L����I��s�+��p�g�R����7 ���?L`�(��1�/%-KP�45ɯ:�B^��O��Y���|��V��,h�/�_J�1����վ5����=E̴��]�+6���QAzx��\S�XY2�F]{�$8��/w�`Xԩ�G���V8���w���j��V�e��,��`Yf]@�{~o��{�|$��rB���O�)`���?dr��{����w=q�te��h����y ����s�|�^��� �lr��)�To�U��%��v�ԸY+����w7�}��0g0v��2{����[�|yJB��X��W�*�W�+��W^HH�ɳ�;�2�y���n���ۋ�J�QǦ�u^�ж��c֔W�7����d��y�l-J[rҘ���hc=y)ፔ��k�e��w���Ҡ�P?�J�S�i<٭&�j���� �����s�+�~�Ks��;�4�|�X�&Ő�x͕����k�s�\�e=��ӕ�*!��r��]��6��0k�Y[�oG�]u�����w�s����swi)�s�U�(ϗm�la@����b�`�qM�7Z����iZ6�k\�Lq8�N'CD�}gw'నd���Y՗����SRv��#��߲���Y�C+����%��tV��
�����Vsu���XryF�Gs�3�`��Ydƍ�Ur}6�ܚ�;�we p���]�	���2�ٝ
�\�?x��d�z���Oeʮ_�!���k)�&�A� � 0
��OBv (r*����O,��%��b�a
��G�+�4�XDh����Au6&yʲ,@-wEE<��$���С�_����B��)�"͒6i���@�K.��f!+���)?���Q��4��>\/���.�|�tOu�`�w��#���0�<�qD�e��庬wd�8��D!�X"t,O�
�xk%�B����e ����+]�J�[ʔ�����/O�$E��DZ�̺\�o��^1Ҋ�u�� �R�4S�Uz��>��	K�}��X{�5K_���U��Q��j��5S�:o��?�q��s��G�'�';�;.�� poiV���K%�_�Z\d՗w��)Z���%��{?] ػ؞ w�_Rh�����9�慦{�}Z�h�U~C��]�2N{{/�*�qY��r�N��3n�E��22�]�d�qߘ�ϗ��V�恫W`��_���m#�ζ�O��1Hp�:m!��B��Ҽf�����J�A�{��$��nǭ��X��
�Y�H2���Ev\�)=N������! �өକ��WXr/]��\e?� �ʛ����S5��K1`
�9��WP�1�=G�{M_Y}@̾���Fj�tH�Wӈ�D8K�"���p>��X����dq������X�H@+E�e�~\!�&�O�&Lܔ;l��ג�lf�a�҂m{��v�3�H�7<�g��_LiP'�X��Fj�ZS�Z��}���H[N-օT�O��p��J�k�"����� �U~KK( �69��K��Уcx�I�kۢ��2�P|��/�U�@ˀJ �=k�,�O+��*������������m]E���޳�lz�J�j-斬u�$�yp[��1�U&��c+,�v����6�ś
�O	ۺ-�;]�蓺S55 �Y���T��5�c�[ "�K���ReK!�̵O=�Lx���Ӈ��G,�KJ"0��) `�m��]Kl��G XQ��X��-��, �^-� '7��t,���
}���+���6c�^�F��ȺQ�H.2@��"���k�zNS��ߗ�4��GR��Z}M�ޘ�<�O{�R�KOy��UO�����{v��s�'/��k6��R�W���\���2Ӗ�R��G�?�7s�2���i��2��e�,���j}�W��'���J9�S��n%��]{>���(�g�T��3{v�ߓsm��xd���&=��M
�1�b����L�ơ&M�)�>��_������p�E��� ��F#�B����I�h\���b
�@�4�jo)[��"�e�Hr
�Ϥ��o|�$ԥ5U:v�u?+8ZAU���UmF}]���%��[��J��=˟�خ`C�W@�K[��lI��AP� ա(l���Ug��U_6>� D$(���P�����s�F7\uR�#?���<-JBQxoNi��>`n\ ,���w)�����*�U�Y�<s����Ƭ:U_���EϻPK�����%MA�s������wOo�Yx��JV<�6�Q���4@��������n�s~���acs+���׾����/��� ���q�U`�O��s��N�Lr�� ����ȱ��
�e�ֳE <���DSjh-��'}��P��ٖ{�ƃ_����+��Y�xݥs��K�Y�1� ~�F�b�o�7j��,�W)k�u䩍R_k�I_�b:ߛ�ʶ����gh����z����m�%��=)[ �R����.&�6���8�Κ��3 �!����z��-�,����6p���5V1]����� �����1T�
���w=Ӆ!����)[���9�0�]�o6��j���Β�G�T���ܡY��Ux��p�1m�fv�.�N�9��l����Gõn9���r�M��b����B���3�k�����pW%��c%e�ha'm\)|DӒf#dB%�_;�w�T
fc�:g����='I���v ���bSҺ{ AHiX����
�v�=r��T�6
���R^���@O���|��M�<�^?¯��A�%R�Xw���*d����ӳ9�x��u=�}��u���gA��+=-� ۾a�� �N��{6r�?v���~�Q	`���oE?�����.m��xX������t�+�z�#g�T��tn�M�_VަO� ��&��+�Vr������SO>���Ū�|�����< [ �`V���#`���m�+`���p��v~��� ;��x��]c��J��ď����Wx�Q��(�l��&PU�*�8��:�>:0�̼ ���G�ٚ�u2,�>�|fi���s/��H�/c�J��������Y���~�4����ռ+o>�%�{�O�������E���� �%ZqZJr�I���R�/�J}ϟE_>�4O ��k�:gyRm�]-L
�����8��d���$�s#L%�m<2`E:\�`x4�X �a���I���Iz�h�#�i��t�r�x�j��؊ϬG~r�I���5$�[vgȁ�H��jHV������ꫯ�O>�$����o��Fx��/�Z�e�%l�	ks��hT�ȕ�ҷ镨t܄xU^�jm�o��R	 X���h���w���4Q�4m������|˗��B � �fQ��R�z�H�S�-�2Y�ǝ�}�8^��;~m~����7��r�ki,y����q`��=:l$r?�}��r����+��x2^ X����?�X ��޼�]�/��!��&�)T���J'1�F�3z�/j
N8�>L ��|��(��j�͂�T����I�?�O��7�|#���?L��r=���Ȼ/{��}�z���.�V!c�+��@��K���u ��v��X� ����/��*�!{RF��*Z�:��ԯR P����1>���3)Yrp�Toc�gV`�r�Z��*X�}Zu�Z6�y�*�m���m�k��j�.�}��˶9f�f��;A��l�/�wҢb��AX���R�����Ӿ��'˛]���Ji�>v���ԥ�Yy���� �܍� ���O^����K9FB^bgM#jЄ�)Z׺4!�{�67g���9��	z5w}n�G�+7����ڿ.e���|.���v;������N�I�5m��%o&`j;��G8i'��b��~���(��}g( .M�v�X�������k�Li.X�fu�y�I��%PO��Be|t����6�����=���g�5�-�n����U�NR^H�㙁q���ϟ�� ��Vs|B��k=n�E/,�(��R����R=�ŗ�% �r/��V��g;�u� ���RYm�vL[E
J�>��^�`ǰ��iA�[�,?�*σ�FIK<
�i���(s�G�qM���u�Xk��$ ��F��L8F�B^Gs�
+�j3�Ku��Ђe�M�`\j�l���1& ��F��^,�?;�]
?�m�X�S����8�%ZgAC>�Ki�XPTr���X ,^�X��͏�>�����BK�C6�C���8�O�S��5��nd"Ev��2eȍ���a�р~�{�t��њ��'�0�b$٭q�N�^J~���8Ʉ37�t��е{Y�*�j��������������Y����Vyc]���~ԧ<"��ݾ��KF*��Wv_��ï�����܅,;
��i�����|]���K�L�)1_T��#W��t p3ɭ�m��s��1HLt鸞��p�歬��F�O���	�{3#�4�Z9�s^�ۏ@� WVةB�~l&wrn:fv���*~�j��u:jHܝ�yK*٧��-	W:���{��H� L�]ь��mb+@�Mj^P,�/�r����AS�2*/�[@��|~6�. ��g�_{m%�F5W]��'Yv�����ǚ�(�J X��U��&O)m��+D���Q,<\�C��(��B����F�ْ���.�6� ��,�~,��+ϐ�Y������(�����R�f:��O��	���pa~���,f�Q���4m�Aٕ��D����
��l/
Pa׷��(��>]����E���L�p�ƭX��~��\\��knՀ`��[��ڂ�l��$�����Z���޳�q$I���R��J����̚�g�s���s����?p��1=۾��7�n��0�J���JU��F��Df"M�a�܀2���r� `��K��F�����:��0I��5� �₠�P@��B �eH}�,�@]ޘ*2W|�H�0��eȎk���� �oV�bAd����Á�ϖ9�X��+�:�4��h6xL�Iohp�?���!��z��i���"�w���\�4:t�Z�cjLO�5/�qy&�?n��/��`Z�Ǵ[�vO����0Z�ᮻ����]�������oϙeϸ*���ua��M��z�R�"}�`�բϞT�Ĳ��i�^<m]���@E.Z V	��s�$�@@(�^_f�T�3�ěj8��(U����7|!��d{lR�q������$����� ��wee������%���q"a��ڰ���m@]�>�a=�Z�}K�S�"���}�����q��I��	�E|�*
߱&��)��i_�I���Ѐ!Ś�!i.���[2}�����Mڈ�7p>��Js6�&1��T��P�V1{U���괺V3 ���e��d�b}�txpJ��80��E�8(��dM���j������ݚ[��Iz��l�s�뢢MF5�L�~%��`��_��k?����Y������V#m�A�cnS⺛���a�l���B��o�c��[�T3<ЖY7봵��cc}Ռ�
�@,�1�R��7c�Oh����m��:T6϶����ij-����j��(`�Du� ��K��q���\U4HЂ����	��� �I��Kc>��_'��I���H�w讏b�����w�{]��,�O�賋��x�4&��ǅ� �Ų�n���fj�<��+T�����9&�dC��=�꾔�� ��ҠY�$������v1���Si�� l /<�Z���ԧL��@"��#/���9G�>=;���i�%-	t�7�%-��)Yg�@����
� ����8F$�1�e��2b��xا��eH66����:ݻ�Mw�m�c�67W�^�P ��QFp���}z�Dϟ��~|N/_� |L�V��u6������5iW
�Efs��#��$i�G���s���>M����y)
�G��Z���ˠe�@�\b�>�f�.ɰ��7N�P�͸�Vw�1�5V*t��}��zp�|_���5��  .3�Cl]�nH�Gg���������g����h��Q�}�<c��w,_�<�0�Ƭ����������.�hm�0�. ���&�Rk��q�,=��JK��]Pt|��y#�p��\����[������ �
���M"�;��*��Uvȹ�1tI���:�C���;q��1�fϪ�s�i��Ӏ��`��Kn3�W�_�F��D*b%���E �^2�-�����ڴ���H�6���0�h�حT�n�P�@#	2�����eP����z��)��1�>e ����,�&P�	��ITD���O�d�6�,Mo!�{�������8 d������10�Ӑ]t���՗���g��w���ݤ��k��V7{�BD	�(�U�v��{�n�K�V�m��n���)��w؊�`9�,�9�AT� 	�U��Ve�K�%g�����ֺ@�t݅�����h���.�V�ն�)�|a�<�������a9�Z�B;�����C�=�k��}ڻw��6��Zc3h�1v+ ר��5�e���Z���?����C:9=�N�k�L%ߥ�6�.Nc���2��,KK�ߡ���ιefթȵ7���Ŭpǫ��ehA�+|��t�:H�v�G����#w�'4������?������(_���\m���d� ���(w���o҄
 �?W���$(Mu���oi��u{
��=��^td͒b|�̶N��0% �16���2
�Z���a���c��E�&�i�� ]��oIKZ�dψ��[-�W�" F� ��U�+H7��vis-0 c�~��m��������f�5{U�B����4�G����2���5eVWig�z��6=}�O�����קt��ª��2��lmp*XH̴�P�o��i'fYK�}˵x$� ٠c�A�W�J�~L�v�*�
��٠�~��������gwiu~�1���˧�k�iЍ�8-f��u��e���z�^�v������=|x�������'���[v�~�f�|����#_9�o�S�@�4[���Js�j��y����-Y��-󦑫�Sz!�$.������")�YZF��>NĒ$�y��\~�ޱ����eUMӇ���� �`>s$����A4�`+͎�3 ���Y��-B�(�A0*���"�/�%Q�JS M��"�U�l'��D����-)�>�I�%�\Ғ�ts��$����B�ԟ
�#h~#Z])�έu�����w߀�]z�p��5D�X��aǺ�$���t���kՀ�T�������j��)�ӠQ�c�Lb_�P�jM�5����B+�%.��a�t��|�{]̀�,�KxW{�6�.�{�R��I��x��7{�}ã����!g1� �c��o�~D�������]�����sa����MA��{lZ`�̹�±W��&՚k��Z�j�������s�r|�2�(N���]�b��@��h�q�>Ԕ�K:`���M�}����y}�k�y�_p��{g�Ez�h!�&ɧ�ts���������&%��]E�o�� �F	H�X̡A�� ��w�[����g)�ǿX�f]盓E5�Y�fѤ��d]P���<�،���t}RX��Y����@���Y���]d-�� 8��lTg��#0�XE�&��$y����a���ms��Ҫ%-iIKZ��%�8�c0���:���>R��X�:��"j4���ޠ�?�C�����~��]�Xp=6�.|1{tKHY����"�RRN���(H�MQ��<��`svb ���^��I�jL2�Ш~�>�~v�´����3��"���1��Y�ɧ���eM*[���2��N��y��m���P%���HgU
#�\[�/>@�������#�ڨ��sn��#3/��7x��JA��O�C�)��S��������N/e������Uҁ��o*�jд(�E��{�����ߡ�����ty.���h�GGG�	KH���!�+}�,kN��5(,H��^X��]M�K?U�v,L���;w�������'~+9��}�����y{���9�
��Ol�����r�|^J-�Rë�:u���2L ����i���?iY+m��D�ŝ�=p@���8N��O�������!rl�'﹙(Jv�8�`��榏[����L�¥{�bs��_k�&\�0�K��idՓ}$�n��-�s4v.�D *����Ƒ�CՄ���kD��f�I�ݢ�~�G�|}�=X�hpl l�������
�Y�ao��ÁA�Up��ڻ�I�����Cz����N[l� :�бP8��2Ղ95��Q�\���_>-���R��i��ߊ<kr��n������g���</@�$��g5?e��zZ]����m���=���=����uOi883eu��At![Յ`�lNj�#�e�*15�5���N����b3��R�oSV�t��6jͣn�,LvV����X�E�κ���3s��|nӀ�E�;vu}�D����� � �ȱ���n��`��P�9��_�VT>Q�<�^�r�L1 �x�d���,)���I�ϧ���F�;�����Y�����yB�ܿp ��1?
�"��/����� �D3<��$�@W6:4��;�G�D��	��~�X��m&a�� �vK���ȍ�,֕J��R��vA8�n�K�L��C�@s&�H��i�M_|�j">I
\-Vq0Y���?9`�%c����=i�,��/��)��?��t��L�?�a�� o��H@Z��J=Ֆ��k�&U�����y���c���L|��}~ҭ�&ժ�D}��j�Dǰ0�+K��<�q����kg0ܥ�f����>]�cz��]ƶ�	8o�e�7�Ѐ^��)u�\�r�B���H��`є������=i�Җ�ed�^�&O諫�=.��˩<���K��o�-�`�ڥa�g@�:=z|�>�����e��1�'f,v+6`k73,(�X��@�(/c���+�Z
��/�X9���S�7o����C���t{���G����f�n�i��v�uǪ���ɗ#�-�=\�-Q�u@X���H���vJk�� W��4��޽���:<<d���.�_�u��r��
��/ 5 n���uL��`�0���M�s�J�w�g��.��>v�	��Ȭ�����L��N^�⣅`>1�@#E;�����.Dp����03n�;<^0�����CQ���$��z���R�&@�����˷�� 5@����#Q̃Q���RgH�..��џ �J�j
�D�-6�.�E47�&����� {>��Zȗt��2�I��D	����د1��=�$.��'�d;�E�+���?�OrKbj�s����eZ_���{;�wg�u\�5���y����F�t4m�g8C�5]CJ�Z�ĩk*��l��!�0�[�+t��ݻ�E�g����;}6���|����5�<'c�]{�PÔW�{�[�,m�.;H�iB�m�4ZA7��%�e��9$�����2�� < �[]i������6cמ��3�*��v�?����//��xQ�U���UA4�$#�g��6�t�vv��ހ��nӋ��tx�6c��>m^pӾH*"\q���mR�\3��0V�Ã���3 _ ah|�;���b���q��} ا ,��R7��7`��<�pB����X���e|h��z��-�N\a����Y�d=�7^}_��,Z�B�FN4�
���tA��e6�1��4�����F$4�׊$0T�\�א|�ؔ+d�-��%�;���8���4���O�^L���39}�����x�|y�R/Lx� �h{���MfIKZҒ�t�I��4������mр;N����-8A
�����!�=��-�{ך4�-0����[���1���\ZՀ��f�nm�r��F�0��=��o�3�Us>d����)�?����S
�+��c�v��z����P��d��2���|�����t�V��\��"m��w}��4��z��U|}���X	Q2�����0 [������da�W��a�� �����tmz���~z���E}k+u�X����*��ޤ��:��y\�B��f�B�[�|�6c�m���И����<��W�.5X���^���W]G}N_'�������E��9�������7o�x��5�͚�j����R���T�y�g!�R64ˢ���� V��O�>���wvw��ݻt��}ú^y�7���kk��w��JLٳ̣���E�Q��i-$��4���TFL�11�q��DKh�0ghb1���6g�i�_J��:XA� �٘���������������9á�x�������0-�{��IĹQk�f���� �x�-@�<4���Y��P����H��tI�^�ּ8����x�r�g0˂���gY�/'�3������f���j��R�����b��ط����('��g]���m�V̾�(ҫ�Q�Q�"��1�>�j!mm#����S{9^�!����h7��|OY�
���E[{�.�/�j� ��[ֳ�Y��,v���,AB����ި���A�z�y� Zߨ���[t��mn5)t9XZ��Ȇa>������cz���N�zf̴ o����ȌM��רT+q$�th#�7�e�7��5�4H)9@_�ô�)����|��M�-�w�jh-�p>����pj���D�cC@Ήo/x_�:�}��?��B�1~Vq@����J�$�^k�4E>!��!��0�HL�%�.����c��A�� �����YWM�B&�|F=������q{I'��h�}�^���<�����]( �@��dM����,������2̣E�@�9��r2�P>$�I���H���b����O#�c���k{O�Ox⟞���k~�U�,ڐ�#�����v,�+* q�L��^#MkZ��c�{���"��\�[I��:w�:�aN�[.����0�HN�u���_�}N�W5റR��&�º�k���6��< ���O���S:kG�A�� �>�[�Tk�� �r���@��J��i����\7��M=��ʊ�E�$�3@f�0�+���s$��=(֏����EhS��sU�x��i�����ݾ}�>|�uО�a�
 <����i�W_?�{{;f��P��̌���[eDͼˋ��zuB�^���iD��:2��O�6"��is�M�z��fp�ÀM��� 2`�D; om�Q�Z�t�_q_�_%s~�Iƅ�y����i[��W�^ѳg�������@�(��<�՚E�i��]��|��D3-��^�����|�_|A{{{��:P���y����7�4?Mۏ�x8��%"���m~7I�M
����a�otRİ�J87IT�1���a� 
"� ���3� 1�Agk6�#I'i�k?Q�ãC:<�O"۵�'�NI�+� � ôe�$��O��r �Ou���$Ӕk@_şJC������ȻΦ�>q*F��%��	2o/H��<`�<1K��� D����1�9J6h#��0_ܐ��؀�.���tX�~��R�)u��MGg��Q��WRb#Hc���٢G�*��u:=��a�S�LBc���ݻ�X^M5CZS��1�2�y�W��wmQ�j��zFZ���.K3�`�&�Y��o�<x���P ��z�� ��Չ������m�7�`�	h8�V�0896 ���vݒ��B���c�:�w͘���*�i�|��a SVX14�O8NMRG��m��Ǻ�Mgƚ���#n�+m֫�������<�kvrMK��<�n��P��|��M�lJxw� Mh}�ʻp{I����W�־�t����R/h��!� ��	��!i�v��$�2?�z�;�t�7�(3���z=��]��"��i:�,������I����ω�s�ɂg���ٺh�����mm��[e?#��/7J�ۿ���7�����c>av���vL�H;�����_,��?+6�{��)
f �,IN4|�z�_o�%-iZ���!��;ڹL,�M'�d����'��o& �� ����C��/�� ؽ�Z�a�o~hs��T h�¸���0&HmS��Z6x��B�P""�ٯ��>���\��}��Q �{Y��?آ��*=��D�~�`�X ��+���=z��}�q�M�%@i8�5o�MS��e�Y��\&P�к�f1`>k8�|��@M��q�V0�_~�%ݻ{�c��­�f��zf,E�\hs�l����y��>��	.^���f@S�ZPe�(�{��=f,�����X	0�$̶��������Va��6�cR�W�`k�%�<�����~�&
�������[����$����A���	���f�/ 0�3xvX7�J�!���۫M��R�����Bn�%h��ݻ�@���`M0���[�X�0��7YAU�i�Td���^zn�rn�=�:���\5M�Y�p�� I> 0&¨�*�6�W�զÃC�u�˕Q����,ʰ��s����VlC��#NZ�(Y�)�r0���$E^h�8y�s�,��D# �`��Nq����/'L&l0�X q�G � \��K�Y4iQ�=��p��u3��b}!�Th�c�@ĥ�[�J~h�v�,R�ϯ�&�l����'KL��iI��}��Z4X��E�Ba� `����)J�-��q�i��k~��a�ׄooٜ�%��y#��Ṟ�Je�W,�l���˦�[@�Z0��QX2�}\��!`h�a�%��.��'eϥ��ӧl�NQ �5� ��u��Y�f���e�Ou�zJZJd��o'��B#��.���
5{U�{e`S?�	_�!M‭������Ps%�2c���V�a�0�s�hdǀ�<���\��LN;�E�A=�t畫�����Hc���r\͙��Xe]�����PR3�����Д�B��[Rqw�����f��w~��s���upG;%چk����"��y�H�E�W�|�22״����=��^��!��Y�����7�6K�@��?�_~����X�L�T%jw�f���+��[��!G��TZƉܱ�����xD[�L9�.���8��m=J5�p���l6�$� �o�Dy���x���rqqN6(��/@2���br[S�&=��'�<�ZҒn�69?]A|w�A ��_�(�7�j�@U�K��P �یt�F9�>&OK���f�]��W��MvF�?�pG���&�;���h��#����K�Ǳ|�W��0o�H�gX�:� WaP����׋�E �>k�{lT����V�5�sg��Û��&�lJ��==�F�5���;���tp� \uJM����������_�J�ww�J"��L�4�m�����'o�մ��D��J��PG��Y3�YeN���> r���?��O/^��v��+�������g;���>�?�ӗ��SMy�R���l'����{�٥�v�y�
��ȩ����(Q�Y&�%J�!��=:>;����"�η��{��ɟp�C�,p�7�H�>`�/��3bgs�6ס�u��K<W���ĸ��_�Jϟ?gh���
(w0�d���r���Y��i�֮k�=>����@��s�6��7����&���ԥ�`BG �~K�K�\�����ӂae����t� X* I̈��ۻ�t|rF�Ng�q�d>$����sh\_���r�dN$i�pG6eG��xY����H{w�n0���q$Rhp�����S::<2�4a�7:�Z��l�F�����M�w����Z�%-�CQ��_�5�XO8�+$��$O�m�K��&����_��E��!��$�MH�,�bb@���"76c6o9��x�%LL�06ք�F��Ѿ8�^D<z��H���
\��=�/��K'�v��7���������eޗ�h����f���yg���E�΀�F���+柝[+���j��pJ?�%� gf�zm�~�������?���S���1���f��˯��&���=hzS��ߋh��c�e���8y�n��Q��Ε"mv�%���|?��3����t~zf@l�M��sj�V(�6�vh��:�Զ�dx"�ā��\�iU9Bx�QoxJ��V���Ӫ�����z�sVC��k	�3 S_�;�6���@_�(�vFd]ۦZ���5&�Wx�^����rN�%�NL���Tt���5P0 ~���@�+�9�[�[�<�=wN�Z�;��r �D�-m����h�&X�ln�M��"�S��B��,�J��x�� �g���I���`>0 t�X����`f����9$�㷄hʽ./�`X1H6����lǇ��, ��ɵ�D�Cv���t��Y�0����b	�@���{z���M��G���C

@i>�_ }�\��[�=[8�%-�i���H�f!^�`���V:�|�1prʀ�?��0��Q9D�Mx�ph�c}�p�V�t���\`aаf�fN�V6�qr54�R�V{Lt�®�$d+��f'��(���u�\��&�ǔ7vbϧ��  �1��0�`�����|�Ak��Ck���p���y�h�ꆹk�=�4H�G�Z��f�no��=��� W�~�4{V�/�i���k��R����LX�#��м��O�7��`�r���ç%s��Yp���9!X��1b	�n�a�k	����z��-m��h�qT�m�aU��j��o�f֜z�NO;<]4ks�F;��}k��=��1���K�6V��a��]��B���}`e=��7�΢q���ܟ4��`@����1.����/�O����d�S�����y$ʳ�w^u��j������m����~������=�EW�E��B��3�n�;F�x����n�2���p��?+Wq]�	4�����O"*����Y�����>�nwY��v��Mh^W$�`)�X���^V��r�Ȍ:�}�C�4X?) �C���/��� �p�Dkl#?��-��������I��F0,���KZ �T�8�����j.`�M���7�Fl����k�Y�9���ئ���zww�H�!t�m���uL����f����>'�$P0�Nl�M%���B:�K����G��%�3!�ɸd@��a\[�� �{�Ը�|�u,�1'H���Nm��*U�%:ouy
�Lz�Q�u`Ve��������L�֐��Z��݉y�	u;-������}��`X��,���M�^�d֝�Yg��T�&=-a�	�V�?¢w����;��U���T�#�U�����;I��j�L�=�ժ0o�i}���ϥ2b�؊��*�:��2��w���Szp�� ߧ��n{��jq#�^%iM�O��
7�����z��@����GL[!,�>�4A���;4��?�'�
�7��)B�݈�/�G�b���v�~����@���"�t���W��z^���.���r>���"�(��Zx$ќ�;�##��+$.�������ٰd#,�b7����3�p~ݞaf��D��o6t{hZ��Ŗ�h��� �$*}-����ߣs�ا��^�����3~��6���t�	���> ��T?���5�Y��fw�9�5��1�~���J�.K��8`S����߿����gi���PQ��d�b�Ft�G����:2f�v	��;PB1����� �E�u��߲�L`�hU���̺����umD�0��A����,k�|�c?�OlX!�M��![2�|v[}:>�Ћ�tg�I�;���^�{ u���0�r5dFnu�B����@�[7 f��_L���\m�۠~/�ÓSz��=�y}�&����#Ic�y��`8H��Ƕ�����=?ـ�G�D��\l�A��ioiw�I��ޫF��A�U+dg�[]���H��C�
k��+�vl���Nq�FǧCz��}˟<3kKیY*y%Gb���*��u N�v$�hv�[I���/�Ab���5�R��Ǿ���z^B
� ����*�/�\����L�����2\��G�ӵ&�� ��}������߳@Y4��V�|"]�D�G2Vf������ϻ �ṋ"�K��mZ4��O̳���k���0)0T�h��յUW��ty �.έ��:5Y�f,ʆ!;:>�ޠO�n��a^1y����v�Z1 ��Iׇ�TZ[��^������g^���ko���86L �$p�S?8[Hɠq���1�P�G̾��lI�*}�R��^�|�<Y ���C3���iig~)}��t��&a��N+�MK�ʪ��y���Z�u�*�U���r|�X��؈� �rN]��z)PbT�ҩd�0ں��+Pwo�����i�QO��l�Z�V.B�*5��Uh`91ώ66F���Ƿ}1�g��ѓ_^�wF�=�s��0.�Bݨ�7o�[Ĝ��A��0j%	�W����^���}�h��W�B��c�#6#�s�\ �|VJ��nA��0�o�<�e3�ʫ�܀��<��|e��>��?6|�o�|��&���h��j�����iީ��z5��(�)�M����[A�Ƹ~n�H�4�3�]|�"��hFa�#�tE���k�S!�w,E8��簿�/�W�G�}��wӗ5��9}^�?*2��7�Z~��� k����?Y0V�"�w�����I���AO[��Ħ>�� iFdf�q~ʠ����dc9x̀n4��#�a�8gW�����4�m�3�=??���:><��ȚC�]�X���%Bk�+�/&&�����E����M���Ƀ�f���D���&�碚�If\#� M��n�7�^��1�s�+���	`����ڧ���l��kܼ�2�I�$Y��xNVu����#�Xm%
������?Δ�'[p�&`��W�nӛ����3��h�h{�J�:�v�]\#Θ�S��'�u����5��B�+�K+��/���^�w�=7��9�;gE��2�!�|���%}��Aab� ����o��O�T��LBK�w��v���~��!���^;���,\�6�T*7��E@�3��_�П��3�}{lx���+,�q�^�u@)��+��j��l+�|�� ���?��w��h���4D�.�\�?��#�x��U���=���<���H�ry�z�k!���_�F�̽m[xmP�΃%,���U9W;;6F�_8=�1&����y�|�E����_5����Ȫ��_�" ,"�rL21�~��3z��1 ��<2@�܀P� J���L jkD�^̾|�A��14�ŅT��` \K�d�Ke�l>�� >a ��v������Y#�%f#֌:N�$��P@�SÇ��v h$H��r�	x�r���<�upH>	�����0�b�5:oAD���7֔��|�A�UK�E������������,L�����̌]�2PVZ78פ�tP��v�6�?��K}�������)5p>�l0�|��X9��&HL��Ol�� _p� rrvJ/^7���^3@��[tgw�V��W� �d� �k�"�yMr
G�Y�ך��f �5pO2��Oo��^ӋW��nu�v��VI�T���LaáM�Q�&��R�2�|��$�"�	ͤMz�r�ڡ�v��2��uǼ�{1'���}��c�����+��>!|�g�����H���_����Q��n�^5�4(0 ���$�:g�mЭ��0)�T���B�V�3���^ѷ�>5��:?k����R�t��y﶑��3�yti�e|w�����ss�/}�{�n�/
���iww}t�cy�0I[��W � P�D?�_�?|`��P ������_!�O�^W�*>����_�e�z�T�@0��(��h� �s���Ǣ�׬I ��[}�&=KGD��'���K�:��WK,�+$-���F��P���������9�J�2�}M�ͺ�\e �V�M'�'l�\13v�V�(��)?h���)P������D� /(�R&�8X��T#9L����Ǐ�� �g� �	E'I�4��x��4d>�˔���w
�ބE�S���K4d6:%rE�i_��0�����������)w��Ӵ��H��!�@a
��F�x�1�z+�
i����� �ln(9ťk�<K�����3N5��ڷI6Q���9'�����G�o	�x+0&�,R!���-a�qٚ� �A7��WJ�J#R�y�(��%�kA���C��gD��^��� �O�ߡ���.� �X��Y˥:u;!�S|D?��Ҁߗ�Ï��|F0��5���k���� 8䪕�V(nG �Ն��4��Y���Oi�ė�U�c< �k����͑��n�u]�U��:����.3���{���E\��n�3���,`X؃�0(���9��??㔔=T��c��VV�4�_�9o+��eb����e�8<ڧ���_�O�����%��?1�Ԩ���B��6���~�pE��ӂyy}��Իc4�� a�{��[�SAXv�ݱ!�h~��EO�/ !\����dM��v�p/ #,%�;��uݝ?����HƁ�O�^������i�so�Y��Ý`���g�����yXyV+U��]�H�~6o��x_��3�[E,|��:��Ф>�R����dz~�i�|�0(ᇀTG�[�j�LH ���#~	��Dp� &(1�b��u�ӎ�5�t��	p5�s^`N�0��x��T�&���s<ч6�0�E �}��#��`ʍ�B>���A��I�x	TP��9A�>�F�2ţ>��@��[�ޛ|��07�߯q�� 1)�>_�}L��{�~�f���k��:;dF@�e4��F�4uٚau���=n��< "�7k����ؗJ��샹A��׍E�.��c���R���DC �8�w�u�����g���nL�n����H�TfW1g�`9��qHg'z���~��}��z�r߀�S�}���Z��&&��� �l=V�X�w�=�4K�?s��Թ�iZ3�&D�c�zMys?KÒ���������4���X?�$�Y�^u�^�����~��Z����N[�/�CB��f��BEvU�l�k�� 4�Y��p]�'��?��	���+:�?6�G��
�b�Cѥq�����[F֡����c�E��^�%�џ��+=�F��Y�[#��+m�>Ư��J�_��/,%���C+
���fO?����Mz�����u�;���� HF�������6*@2�CK~`���/M�/i�����,�1Kf}և�&��Y�~���0������f̘�;�v������?������1AK5�@$�^2�B�"B~������kw��o8�D�D�Kj������"\��|0r�f���#`LH����?���ϹKZR��i�8O�j�
�R��)�����߬�����{?erA�KW�Љ�Dk�E3�2T�)��e��C0C:4��_�%z�����t�����4ǖٻ�.�4����0x]���������y}BGG�n���B�W�P:���UY��}E�~��]5�k
E.Ya*���
gb��< ��I��2���. �[��0�z��g
����h����/n9���j���79"N%4d�J��
v����tl ����/���!�}������u��mz��.���ZȦ�2���C�����o�:���'tz���j3�+]��"���߁���-�}
�u�t��w���eNȱ����K��A�	���Ϟ�f�N�{u]A |���7I[��c�Ќ~��RҾ�w�`Mn����]L��I�]�~�l�b���hM��E�y��`e|^?�"Bp!=.���Y�u�(I��J@�4�|�T�i���S�Z0&̘Q�յunC�z||DU3�N�$<?���ͬŁ�7HL�P��5]��@����gX�٬9��r���]�!u��Y3�Z�J�+��`<|���/&лwo���ŋ����_�%}x�)�w6R�^�%	>�v��w�W��`WC[����)J��[O�ᘤ5\�$�e��k�=���1`��ٷzfR�}@'�'t`�Wo��`�v�3�_  ����~p�v��{�޾1��s=_Q�Zc�}z	2#T1��!�2�bG��>�ai0�Q����%�| �X]-�f�D� ��w�i�!*������I�R��S�����Y��u�1rY}皇�~m��4%�Pb�L�d1u�=�π����^�4�����;�ԍf����{r|� �uѥ� ��ce8 �0�6��:pux`'m�dq䳉(F�Ѓ�ӘYq��C�+����O������`|n�Y�:�\���D8�6����V��E (�z�`��5���'�^̤%���3|k �?P��7~C��.�_��m���H*((��^�'����O�>e�����"����o���S�u�;����UѼ�-� ��`��߬	>����_���~���[�W��D^�۱���LD�a��S��XvI�!�L%�Q���Ao`�r QՀ߭�m�������X�U5����������{Hᇝ�K��g~��)P�z��ӵd���k�"�ᛵ�_!��x�H���)�'N���n���'����",4缏��g�9��z�n����3चhlȘ����=6u.���
��"3���BS�"�G *��Ӹ
��W����*��\��]����J�c�u�6��$ �E�v���N��� �/�� ����������4B�����)�K�uL�p�%ܾcle� �}1n��NY����)=���e�g.����E�����s�<�T�s����A}����Մ�U �-�c�~���"̟ټw�� V���Xk�dހ��!GA#*~��kW�EZ�(k����/�h~d kWYA�JR$Ah��Gk�<;����;�t�� �����[6�3��X���~�f��h�F��������46[�V��7���RU9��DƉ���9���͕j6p4Si�|%��}���"=��� ^ҧE)���Y��%]�3�Ӄ��:<�v8(x.���r�YإT.N ��۝��تР6��0��.u{:�hsЯ �s8�4�p	"6m�s+e C��"��FJǵV*A�����@�/�jkk�vvn�=��$���<Cf�@�2�Z�,Z���\��O�֤߯hz���(�Ԩ�n��"(�i������s��Čs��$��x	j���`ƊC��j�{=��l0|B�*��$1�f��1�0����O���^H��u �?�߃N~��\�k�>�cږ�%8Ȳ���E�7d�Ck$}e�Q��A�����9t@�z��	��5�A
���]:b9���GM0���`ݦ�t�Q/h~qH�>��U�- ����vh��h7�	<�����Zw9ܽB֫�јg%wr#���,ٓ�ٝ��M���,Ͼ^ �0=v���������f���4�_�5}��W����kz���dRS��EַW&o�n�qR~��;�0+-�X�ך�t{g��ܽÀ��ݻ����/����g��#m��L�������CwI7���#3�[�9�OSv��h'��	i-�d>�R{]�|[�XD�����fNc��.��/���R6n��Y��3J&�d0��S	�%1����e����j�*����� X.��-�?|@�Y�S~�T&�@L:��0�|]mN���i�����Y�)�FNS�2�:z;�%��X1[[!H@e'�F�ͦ�X�j����Q�J�FWO@�)l�{��,��ڎ%_��DS��˵ӂ_Wङv��\ ,����h�.`��*/����xE����ǂ�Cs��P�`<�q�����rb.xO�(>�++)���:A0+��{	ڋ����X���Wk���Bj8K~`dxA�0� Ɓ~�ubn^��y���Ab'H������9$9���{2���>��U�I��i��e�F3Z�s�8?�H�l�e6o���|ek����*�>;;5���9�9����ρ8����DIx~���*fc�q~`IQ�A��f ��m>vͱ���/�؀�ϟӳ��x"���v*%;�A,�&��� �3	o!�k�)o%�k��k����p\0뾋,���ZM>���u���<�)��%)g�[��A�u�,p�Di�[Y#8�M�k�	��l5w�v8J��V�&^J�GRE[�p ��BK{{g�������?cF[c ��nd
��� ���� �4pE�u��q�-_�w5�>��k�O�~���
������J�K)pI�*�#�9J��鯬�-���&��1����l`��9s��e���
��7ig�@�:�D�"��<�%s�r�?}��>K�����"�B`'c
�,�4� m ��`���
Xd�tA�(��(�vU����󬻺]Y��ڋ: �KRh~�DS-eh��?�v@��4�@�h���A�]*JE8i�1���Q�h�\[�� ��^ ,`Ro�����)=y����駟؄g��.Ke���k��7��������<)!�I��u��K8���H�[�[�@rks�՛���&OdL~��'6s�#�L����Dj��H���7�XҒ�(��ML$���U��_1�����K��^'�&�F�Կ�w���M����Ä��w�1"�e�I��M��-�=8�6�>��Y)L���CC;<�U�{��,�T8\5 ��Ƣ�3�%�um��Dk'+��s����_�fk�j���Cأ�֬fH4��Ay�,M�Fy�s��A���X���y��+�W.x ��" �����$}f��ۑ����]��,,��l�� �䳟.�������Z�نH��5�����	����)g��at9ұ4@Z�% ���pF���C�^��������FO�O�R�M|�Q��#�7_,`M^n�w������ߤ_ŲB��˳$��*��+�_�M���uB���º [|�E#�����婧�<c���1-u�����NTs=n܈ы�k��I}��o�s������ ˆ��zz��C�<�x���o������r9�5y�?o� Vh�ۭ6��=>W*�x�,Hqj�:ߋ|��9Ƣ����9o���� pD|�"��&�X�b����󗴤�ȵRH������_ŗ��%]��6�r7�<�$�0IS�GE v�y�=o�L1GN�N�2�|-�R����/m���G'��P�>�(��$kHh��<[_k.���{z����Zah�p���3��j�g-#��E�?��$O#T�Y�5z~ ����V|hd����$���t�dyB�č�y�t,&@W�j�N*ڕnI:}`L��7�'�G�X�@�'�#'�$m�{����40�A�����φo���2}y�} Xʒ�	`�E��#�-e��"��Ȉ�cJ/��5�������Hl/༘��LkR�"Wh�N�{p�\���۫#����ٰ���� W����WA�����胙@�R���I��=��g6��OK�	I�7vHf`���
�4&)^$�:�fB�h��<�v����tr|����߇I%�(��#I.�*�gK�Thl /G󒮟��f�j	|�$�2K�3+�����@ɭ_�f���^M�S�X�P�W�ӓ�FO������Yb��x}Z���I|4
c~`��$�M4B����c-}��&���o����y xR݋h<�2���e�_�_��`�����\u���1q9��#�l���=hM�e�W~1���0i[�4VYm����<*����YQu��|��� �"��Du.��
�1� ����Y.�mb>ڀ?�4���f���h�u2Ɗ�A�����Z��gC �>����m.*�}��k���
��}1��[���*�m^�n��d���A�n:���r\ޣo F-#3i[��;88����&������R��@��I�0�h�|Y}�$}�� ��`���X� ��9Y�{���I��ʮ�<N��VmN�"�%-�R�������]�i �0�?�O�5����f����|Ou�S�w�4���ʔ_ksq�0)�U0}F�,<��A'A�(ӇF���q�p�	�{n��&�؋aY��u����`��"��� ���i���ʘ�vX�����5��%� [A��}���4Z��2F��ϋ�F�#�\�'o��`����_��rލ`��^w4�Q�]h9��@��|r�'���
�����mwQ��½ ~?�D��4�t��f��;���1��Q�߳1�/b�����yegQ��$,T@��a�~���gm�C���6�FW��
�|�]A��#Y��UQ^��L�S,�Z@���� Ӂ��"�t��A�#K�eA)�l�;l���M�c�Ȁ��k��XX�#�밇�u��=S���@V�/8)C%	�)(���ZҒ� ����.�����6�y6rͼM� /��¬�2c*���x��R�$ݽ=����3	xU✯%��2��KDI�!NMC��9>L�X�;T�P�8 |���7������3>;;�Ë ��w|I#>'����0�`���������2@F���(��	pM��J������V%����f$��Gq�e���H��!4�������d��	�|���0)�c1������-g��΃�Gy�\�!H�S%�7>�ǎ ��9x�5M�H���i��v�#.��r?�����ё������s��
��@K=���V\�
�楉k3M_���	��\���0S�d#J8x-y-�b:����,��)���0��������G�}�\/�����������U���k"!���,��&_����8Cj�l��zt�~�=�ȵ�/f��_|�YM�q$�a"�ƳB��ā.q$��Fa�b~R�9[ZU����t��=�����f������Y}�!���I��E�M<�Xx?(�+1�􇜧7���#�ݚ��X���hl��c��|�v5��g�b%�g��7Eƕ6������e�����5������O((����8h=~HE[+y�u�-��{�q�c��Ԛ`�K`��c�7��;�g���y�����L͒�wu�s���(�`�m ���"5�z�ԟWiᤅ����=�4��
�p�}��)�3���8� <�<����jne}(��w��� r�����_	/>�lya0z��_$j�d��e�咖���)a���ˉ��#��I�W�|ݛ�<�����E�j��6�0,��;I.@/�t`��'},eZh[-��/cD�>%��phuʌ��D`�XD�IpH�`�<yBo߾������޼y�P���h� K�{��6o�y���j��kD{���_ӿ�ۿ���,�" +���yC�i�,I��uV3, X�ta*��(��	�G%i%r�~K���c��h�Y$����a0T��Q��6;����o��傇��r�h�-E�_���� ` D�z�5�Ӭ��k�u�SiI���g���.k��>�Xc8��x��=��	΃տXk�aF�˨ �̣yH@�p��y�0i��`���9��M|������.@�W�hӅ���P�:�?�
��5�8�$bpN�N�P-%�d���5N�O&U�y��D����A�X�������7A�3?���ddw�4���㥀h�X�>?��X��E�ބ�J���ޠ,?�i%�g��\��-�����yp�E�X�&�`�)��=Q�W�)�d&�81a�0U�ap�ꈭ�8�I���I�V�8x\���U�=4��uB/^������={�2�n_΢5�Ңfi���I)X�X�̸�|^�|c~fнf��zK�"���G
�Ե+�]���-Q �Z`�"$����p��0�
�A-<N�y�#sƖU2@� BX@ ���x�c�-��z��OE�Sk��8{��TQA���{Ek�}��>��]�wY�t�ݱ�����I�/��"y���5��Uc鮟:�4ʇ&�`< 4�&� a�h�]s�,�{����xJ
��$u�h~v/7�x�ལ/�6N�zn���J�g)O��+iWBZ"}�\7%�p}�u
$)sVZYm����Ϣl\�~y�]�8��C��H��p�J�3G4�!
]�aO�e%�?Krql��F�	i���#I���4b@�o�E�|���<���sK���E��1�q��~�c��H3F>s�yhQ��f��1/]'��sE���{���~$��c��`$p��5�hX�0��~��eU*U��V��\�7�&�#�i��3p�~���D�']�{�&�^����C�2�WQ�\�r����k�LK[����aV�"ZS���Ӵh��(E'cѐ� Sk�Oޏ��� �cy��"���Z��?~���ڰ8Ă`� �2�_�	 ��a�Jf<��e��*���	r`���C�h����Xª�*���Y.O8��>8�y)vנY�p���ɷ��sa0�@�q�
�̷�_�
�ߊZH�V�#Љ����Zd���_���m�ɚ�zdnhshWÙ�.�O��ͯ�=���3���vZk�g%^��X���Ǻ�Ԭ�v��8W��|���:O���5�nt��u�0,�t��]�4���~'E�v]���Z�1�Α�_�έ�0M$��K�ǣ�ċ�������w���EL����%��UG9�r�|�4I�[�\�o�F5���g>��(��{Y���{�_���8H��k�p�����>__���m�J�F�+8�Ԩ��Z�B]�S �J�I�nd�3::i�����C� 3�_�h(R�dO�)c�m�葦�0���i�`eiJ'=a]��0�Y��1暺j��I�X3��0�y��R��IGw-���[Y�a�V�3����mV�^٤f�L��_�
���Q��r,��ڽ>���զ�Vǀ�J2���%B��r�
}hl�j�fz���Yk�X�5Ӛ^}^�&p�:��N�~�z�k�F��iޯ�s�_�`�͙Q�1� Q?+�m����E�h�,��4i��~�2�\�m�����F���<�BE"?%�Z��gA؈�W�-�:7�ϸ���u�=�2"��_�����2�Ղ���g��+@��)�`�a�A!c�FL���' �1>�KZҒ���O�\�����y%��E�]�묙?P
�R�
a�(3�d�R1=�vY˻��J������;�po���n��Z��l���i pX��E�Ooߝ�����'���{Dp�R�0t(��Qz)����J����=L�vW�f&1+ �g_��< *��W��p�<_��p��P��fH�Ff�Z�R��Q����'�2���f�=s]��W�t{k��ݡ���6im�N�b�˕��д�զ��S3��ū}z���O��M�fdꨑ5��z��.H�':]��j�| k��\�!Yy��Ɨ����<Y�.cR�  :�ɤ�`MX�u�-B�����ɳ��/�nAs��,��%�~�kОׯ_��3ڃ��w���g�[�iɮ	6�> }P���[YT�%��`=��9�5N��>�k27!�����O<`A�ٟ��gz��)�i� e�ut�~��KZҒ���1�F*����h�e�nM�����L-.�3N~�0Td�h����0k���5z��.}��}��=ػE�w�h�i�̙E� _�R��݈��l��f�m��	H9:�H�;}U�$�@�6�Mco�b�f W��j�&�9�FO��<��g	@f1M,Ri�vd'�Y�p���j��6���z��}���ܥ;�6 F����e��J ��0Y5���l��l����x���<{G������p�c�B֜^��h��(��Ƭq�ߛ;�|�����qV 0�C�Ҋ��B�E,���n: `h���j�]�`{�#6� ���y��/�/� TW�7h��� ���k�<��,m��.�k�on��"k���H[.i�ckY���1���#������ �!$����s@���u�GK ��%-iIK�,��T�I-�A,������I
������u�a��J�����.��]��6��ߦ�翣o~�Ѐ�ZkF-P����!�qD��l�5Z5��v�B�����z{D?��������/'֯1���m�����~Z�|��G:0���~�y�p$�H��V�����5�>���Т��h��������}���Xr|g�"�]��Yis�������o�����f�V��/ca�5��Z�1�6C���ޥ��ܥ������^�_������_���}�qXf��K4���Qy��ѵ"q��5�V��K��C=G��hK��_�[������[���E�"$�B]�	 ���&ۋ&W@�-&�'X�P"�D�_W���X� �<4��o߶y~����0�*�":�2u@� �gZ�5M� ���I�6���o�N���Y�U�,s�w�{��$sZ����ygg������o��/�L���Ǐ�O����|��n�A��r6gt� /iIKZҒƨ����$��$��cd]M�os/
�]��<4�F�)�(	�ȩg��6�PĦ��4h��T�mm�3������y@_|�C��a@�K�~��A�`�A��i�X!PVV�\� ��I[5�7a����)u�m`��X����/3jI~�T[x�6�tYz��>��A�=��Ƭ�'�<�,�2� �h�v��q�S#�6�j�W���[�ۯ��x�`�j�>���F2c��$����B�������Xߨ��M;99�quz֢n��>���<�o�l�ꑼ�'��j��}����=o��em�B�
�~�W)T�>���("p̖����>F���� ���H�	 �}~�M֚_ d�_�*I�����B���#l��I�t����+o��[���������a�[�n�5+�G���s^��q���KZҒ���1�p.�yy �H]}����0P��KL6H�5Y�j���n n�Q2�������;��oҽ;M*�-j]�R<l1��<����e��a��A۔e I�Nam��Vj������#��暗���w�f���#k-~��=c���asxr]5}}�x��$! �M�S�GխKV=gOR/}��-�g��xX�߹�s!�G��Ѥ���3���N�o5�R�ҠNèm��r�-�J6Z42O���X���W��K�R�>�����;�w߿�v�ĔQ'
��ӚE����ӿ.��@k�Ƃ�D�w��<�I�E��I>������|��ө���oQ��"���B4� %��.@0�8f���� ���ŋh��ý�J��n�u�O�3����U`\�]�P�c���_<�X�]��ub���������w�X�U���C�dC@pH��X�q2�/9o�| 8ȕ�\�vIKZҒ��"ڈ�b��YY�����Иx�u/���]���4��4:f�!�Q<`Qo��ݻ��/���~�>|�*%Ì.h883�6�.���ym�*��2������VWh}m���os� �G�hY_M���A����6�����h>'���@�&�q.h�گ�Q�� �:�e���2eX�O�mȚK�g�~�i�]u�g�3���@`�о=�	�T�����I�v������mZmB+l�C�2���FeQO�9`&f��>���T�4i� �������q5�w���ٵ��)�=+
�&w��gi5�ӀFޥϤ8Ok�S=N3�#�F�P��s� �m/H4� �8���{��=<<L}{%�����lmm1�Κ���H�o��DX� �&�Z9�w@i�iȷ����]�D��F� �+D�ϝf�M��<�-�+�ov��(���y�X���O /�풖��%-�&1��)�� �g�G��4]&tC�o����g`�l�#h���F�m4V������w����:���`He�Z�t<0 � `|�
��a�h�1R��nQ-P�V3eާn7��/߳)"�GQ����pds3�QF��<F�h�$W#�l�~�w,>\.��r�4u�r}��j]�O3�.hv�v�׌�c��428*�H�����T>� ��.�WW�������szx�6��Oͻ�`�_
�d��c�?l�Ǡo#���	����a^Ku���!��/����iπ���i��MY�L�s�>�%tp��f�:���Gc��X+Q�@�)^����zK^bhru�`h�;�� 1�ja�M�[��F�BY��>p糞�V����w���i�'�("�F��S>���ݧ�V�Sl�E�p v̶���y�Eߚ���%�]Ғ���E�$fS�[cW�fՎ�l_%�8P̅�)u�yxYk��c-WJ��ޤ�w���mZ[)S%�Q7�RԀ:��lw��c  s���k���5���{�1H�ʬ�{{��ܦ�����1���,�(�� �H ]��W�ܦ�I~m�������E�I*"��AVD���n58ҟ�ݭ��{�c�9�a�Oa�݉�y���k+u���}�x��6j,T�`c����8v�}��< ����
ՠ�a-M���81c0�sU��ڠ{wn�cی�S���9�o^|}���H�&��4X+\��!����>}����>����J-�O���h��Nk�� �O����Y��=ןS?��1/a���rо�����P�r.�Q������	�&}W�����r����~�+�>r ��%-iIK�J��>w�(O�����(�F�{�P:�B�#�Bܠ���6 >�ad l�K����+U���P8���wg���)]\�ث�V+��j�v�V�޽-j�T�^������&�P�A��^�;����:��P�sN�*m��{p���0<ojf,����f1dn�\���a֠La�W���]�f�\��,� �)e��f�m69=��y������j�6W봳�F��ҽ�M*��}���|�>���1�%}ppJ/���y���6k5�\[���u�C]7�Ѱæ��IGJ.�6k�{{�n��:t���?�݉�����Euu����#�jM��5���⺔�cA��+���:�aP�b��j���|v�]�����f���X�܋�`��p �J��g^W�|�üu��o�zդ��U���_V��I�x�y	:������΃��h	����%-iI���(|hЛ�	p���}��'��̍�`Dׅo�`p�?���a�h}�n@�)�[���"*Q��3�e�^�2 ��	����0 x}�B=SVcu�J�2�e�ۍ�6�M��\c��Q�:]��R752`jh�B� �����;b�c�?��AѴ��sZ{������>��I� �w�,� �x_вh�jU�Ҳ)�y��ww���û���-��^5��u~�V�R�Ӂ/ߞѳ�'tz�e�g ����D�z�<���J!�?��ҕRLk�*���2 x���8�1+O�o4c�j����L�.O�-kͲ��O��t�S�[�;v\���r�/
����֐f=���a_M��I��#��ĵ�&�+�K�D 2+�kˬi���k��]�\�I=�����A>�-�<?�U� /iIKZҒ�t�R�O�S�K�mJ�џ��	�?�+`Vhsc�VWj��O�!�� �vwH�������0����5m ��JD�� ��~� xc�0��3!��5��J�L�=ޣ(�R��n�pה�0W�P����������ݻ���h�|~r3�N�	�$�S�usjO|��9s��\A�����9��F�A>d�q��-j�[lp
!�J�L{�7��/����m�X���B��������x}F�_���Áy�Fj���N16N�_�����G�.��_h�ڤ� ת%ضH�v�>��̠}��>�sai����9[@h���F�:�� � �Z�pi���>V��7���{]rʦB+�ܫ�% ^Ғ~e��ҳ~IK�P
���~sI*pZ5`�f�z��ڻ
rRrHg�q�����a$/�ttԦ��u��A�5�%SV� �J�k@m� �*5M*Wlp����:��ۥj}�V��2�	æ�O��A� x{g�?~�+�ſORhp��3��&�Flv�w��$�:��C]���5\�<�[҄�� ��H�Y�U5 b:�h���9G�=5 i\��;Ԭ����
����Κ�}����)*�DMy%��wh��C�N@�~��Mό�A�C�ʅ���66j��ڠZ� i�eʉaeP���&��������퓼��e,�}�1���bv�y�a��&?�ۭ����3/�T�($c�y~߱N`,�/0>�:	�a̓���Mo�&~�3�Rw-s�k�X~�4�Y��]7e�fRsy:(Y�s��Q�jhs&��% ^Ғ~U�}	|>U���O���W�:<�qj�����o�o̚��#��d��b�9I���Cq~S���Ц��/=���h�w���M[�SnL�^�2��T��?{��%�q�P�}��G3�(je�^��w�;g��w?�'�]�ER�f�c�{�����_$d%P�v�3� k�&��H��u�w���[�Ͼh�0�X LM.w84`�?d��Ç���^�x�L���T���$��</�a�Z����T��� ֦�ڇ͍\�e�����RY�jp�/"�~�����_��z�3�|,E}6O�Cj���)����}#@�(�,�=�2���y��h0��y�Ogg��E����Q4��F����:�M}�����uc.s�
;�2dja�]�������߬�Z���<T%�j��R�0� n766XӋ�#�����9�!�<�$�}��i�����}e�yv/ZV�I����,�r���j�ݵ�*��\]����+�ͷ�	�f xF�.|f��6Ӥ�Iև�YC�jm\���L�B1]U�O5��?A�~�1�e�r%�ei`|գh�u7>�W>.�:-iƶȟϞ�䓘<�����Ξ8H��'L|R�2�F9 ��F�b��~p]�~�>)��C�>�q��G�z:���3��9��l���g�LN�h>3 )K��A
(�hз�ťE����'.M��U�/�W�8�V�Ǫ�|u���������Z��v�!�n�ߣӓ35<���g~��iЎh����U���<0,�k̘ds<��7�n����q=�C�c&��Р<�Z����9��!��Hr�aG<����i�{�������8-2u����%��&������d�M�\%�s��o����������E�+hz��ZM0F�&	�ý�`y�>�؛��}���.[��wvI��
��u����4�_�7�&	�:�����|�`R}f ���e�������{{5�zՁSp\�e���2�E1���&4j3!���	��ĥ��"�!��`�i{4S[��t;���l��y�gɷ�[K�}רRR Lx�#���0�q"y�`�6������sZ#h�a�B;� $��(4�7i����)b\����)jڴ��1���Il��To�Q�٦���z���b����;���Q�>g�kr� �����ۿ��VVWC[#��_�!�ĸ$��>i�F��nJ׬�np^�;�9������u���I��׸�.�[߃������觟~���M3��YkjǑ�;�=\[��_ܧ�~����a�J��72��4Zh�i�ұ�q�&���:h���;���b�;4���ha��{�������6G+�`&f?రETEH���$����O���[��yw�Ӊ οw/E�롵۲�]�����N��H�X z������~�����Y�@W� e\0����40��SZ�_V�I�����<�v�,��X�Y q�#�£KP��M���h<ʺ�S��ْ$�;\�S�\&�K�7̷K����s\��"�4�[��� ��<t;Ό����q�n�����o�fL'E1���LS�MG�tjp�>GH6Gwc�k���c��꣟-�|�o����i�F�3��xU���6��>���/�	(���X�=\Ft~�3�d� b�x��AN0d?�8��`XZ�;G�gC��=]+Ԁ�i�ѡ���$m �B��p��� �Z9_�l��nc�~��9���<����7 �a���0J��9�_�gͮ���n���L�o�T9滿�L�^WE���{�8��Q�r��|�����׏����9���˗/������k:;?cr�@�{���_������JÌ�e����ENjNg42 8��{�l�����9�"���o7���EZ6�kn�IA�B� �{��c�؀! r $ �$���Z��Y4Nr)](?Wq�~��L>�\a�$��GW����}����Ʀ�YWH^PB�� -���c����e���S�	yO�*�&cD�p\#�ʞ]�.Bz�@_����
��q0ݻ(�UIҢ��o�zUFz�����������}�'��h��>����ďSi!'`�&њ�q�2M�� ��f����P���Y��z(��k$�x����(�u3�Mz��Ues�� h?A!���ѹ*%'�0e`��U��n�6k��M^3�Z����}xH���\%;�l���l)U)����v��������Z�����җ_� �@o^��a�}���,.�����.���i|�y�Qir������=���s::8��r6�j��:�й�HIS|�HU�34��@1���
�G�����>��c�|̖f�]��|���N�#u�T���21�D��OX�vxt`�J��P���q��\�[ۏ��}䌎�Qm}FC�ؗ8�_|�����>��Qߔ�<�wW;�f ���<5�x��@3Q� �Nӌ�Ь�Èz���G#�-v��"�k���=�s��!�E�l���/߷~?ET_a���0����hA/JE��_�Xǃ&���޽{���%0��� ��o�g��@�&�o�� �5�\�.}pϸ�<�����u ����[����l�}]��w��������<��|�3��@p������� �ь~F$`�{.�J��J��Ҧb�Y��N-&�E�����y�Ϭ	$nl��l�I�f��2� ��\�o��BE�F�5<Z�+�+H�
��R|%@X���;�l�wyrrL�{����.�=�����7[4�� L�MP��/P�GТ���Q���D69:��2f�75�R�4`��y72������ F�ց(���(�m������`=& �( �t��%������qY��"0*%����
��������X67w��Z���ܧv��b���F#���s`���R� ��;+[�%��X����Qh@��g}�?4 ��0��ħ��mBEI���ķ��~�i��ְ���
{/�"���i��u�� q� x����= ��دp����h�*����]� �� *Y��|�WMz_�`�� ಹ9&��PM�~y!�;n�<Oܘ ?��rE� A���������w[ <��e�����Qk�Unn��>�0Vf xF3�э�^&/-�+M(ʀ��#�i0U�����/"G{���r7>9�r����	6�����ﺫ ������I0|k���L�|tC�["��CNa������iu�.ͷ�p=4 ��Zu�n���i6�o@-
�@2�P�V;d�_as@��[��{Bo�lѫ�[����Z�9��M��1�u�~�F]�|�2&�v��E�	�|��|@����Ǟ�M�1������^����|�f\��ϙuc�¢$MQԧ��>�}�Mk�;���<�{��Ż��*���4c�� ^5�Yu��<`����&��-�u:<����>�y�M�wX�So`l5�>�Ӷ�}7��͜Ϧ�q�[k�ǂ-A��k�}����k�+�Hjmg���d ��	m��y��M����o߾ek E���w�Z;	�W��Hz$"D���1��y1����:5��.�gF�D0�����oi�~�G�w�e�ߤ{��e\��c۩��O�N *��L��o�1�_M�a�ux>��eBz��i���m֙^�z�^��r�8k����/3 <���R��"�����Rh��c� 00-r�-�H��I_����I��`$ܠAr�*��4����{�ް5�
�ǵ6�f߽�sD�Rsg���d��x��df��Č5f�W�7@iуuH�.�E�!S\�Rk�A�"�o�!����2"D�����xH�_�����'��ڣӓ#S�j��u�8�G$3,.�c|��޽�"鿋ꡯ/씑�F@���� NR�p:i�5� �� Ի+M��36:�lI �@��AF�	��6�G���Ј��W`�C���;tvӛ�mz�|�^�ۥ����ز�ӷ�
���O˛]D��]��	F_=j*(���ИZ-?��a�^g:$�4� �8��	Z|CQ�w�2��M���v�|�ם'Xƍ��]k����4<�O�Z�\��(�@���k��4P-�#�q��B'�p�ZD;<<���z��� ح��^� �hF3� 䓘_��wD$�"ل�W��=z��4�v7 ��)�D�O�e,|�H�hm.�r�߿ςHse��Rz����â�{ �]ST�/> ,�c���+�<��Kj�$u��d���'�mZ(0��0��u���Z\�{�3���=��{��9E�>�c�Y�m���i`�F���A5n�`�thw�=��/���|����3���Z�<��+����A!K4Ѥ�C�k���f�&ic��2�P?_��
S��T�����[��zal��@�9�z��
��_f���;��! �Ç�����}h�5�Q��A?1[���P�È�W~d9�l��~Ԥ��}�����wo���:<>1c�e�R�����]v�1 w�*#������_�@ze�d�)+[�.Q��c {��KV��
�׹� �������ڊz`��?�����E��B@2�ٴ����	a뤋Կ�y�2����0�����:�j �"���v�#�__��y ~C�2l���~�4�>.Є_���|��������s:�I��\D3 <���H̅��GC�lwX'���+f�u�ٰ�yAc��L$o+i�L�xٌ|f�E�̈�@���y}�$p��
�u��+����.R����Q��E�% �s��Զ�ռh�k!2�?ءW������>��ݻӡ��p`.�c�s��<"yf`�#�fۀ���lf�����z��-���&�C���3�Ux7V��� {w.�+��n��g�G^�)�7��+)�L���;5�[T�.>���ُ� `�F�Qb	�s�eßw�?���}��Nmd�0=X_0��Q�0G*�,����7T�Z���4��C3�6�����/������ǈ��e4�@���i����{������������6_T�2*�\���6@¼'��9T5jrQ��c�:Ͼ��`��N]ͯ�K�|���M0�4�A�v� ��'�W�U��� ��?��x&��"k�i�[d�PEV��"�e�K�g׺�L_�{!\��ܤo���Ǆ `��}��n��ޣ��R�߸ `[^�zE���9������$����gE�`�u��8�7H�զ���	f�UH��,κLa
ˤǷ���"����D���u��"fep�V���e��i�i���7w�3�z~ȏ�}nk���P������џ�<4L�1����~��c���a:�4��h8 A��^V֙�5�C�͜h�%������/��^һM�/"͑a�;��W1k�P����k�'7����w����
�'�V����e!�׶�:�{�U�E�D+�O��� H��ͻ�'�2����C:<:����u�m #
�㇫ ��3����w�4H���W�:�����hc��������Џ�|O;{'�	0�o�g��� X�\��<J�  ��IDAT&-<�����h��*��}GE�:��U��n��yn@@0޽쁾y�[��9��}�f��G|tEx
�Zt����3��o��\� S ڒB�����+h*��*��o�h�"Zm�O�" (�\�+�NJc����3ɂ�2��T��,���?���򗿤n�}����~� ����<Ӣ!���RVY�� ��f�����e��UY�|�n;S>-]DJ�Ɨ�3�t�� �*MS>o�����W�f�=��2�T�ν�L������Q�%�a�h��"�M�#�o���|y'�w02��is�^�آo���^�zO�HiS3 ��<�\ΚBS�@��'
`F|�NMb檌1��L�}�������h|���k�[����˼�������q�? Tk,��#Q��9`AG�0�}�����kq���Ӟ �kD'g�k�	���5�����逶���?m�w?��/�x����������
��$�6�a˪��I�^X߻􍏢�E���v*oQ��jZ�]�� 
?\	�'tѵ�J�@�6��1kHq\r����O������BȦ� 1�F;q� R����
�B�B�-Ϫ
Fy��}�2�iU�N|J�8�vZ��j�3��v������Dũ8=k�^3ݴh�����	2�h�g4�}Rt���S!͐�n0��P�Y�|�VNF0�`��0�̜���ӷ��nЫ������ߥ�w#�isd�^��3Ø ��hprD?|��^��e-��i�lL�6�(�����W����\��ߋe��*ڑi4�^RL�/�#u(An9 ��.c��0�a��r| ����"y������z��I�٦Z��d�a,>�V��Mf���{pxH��F{�l��,l>�+��
0@�<���ߥ~o�ywvN���-z�n���1 �7;4o����\�H�䇻Y�������1�e�i�gW��
<\f[������Y�z��;b1_���� `h�E�/sR���"��q��SLOQ6�����vp&ψ!y~]��~|��:H9 ����Abv���y�����v���溠��]E�A����>�x��ڸ�TS���~��2
�X���A��iJ�8��\���(ϙˁ�ٓ��Xuߥ��{伮��}4�3�ьn�&0�Be�6��4�4Ŭ)
��qPK� �	����	I������>�ãSz�}D��ӽ{+�0߱ ��3�b�NO���c�5����w���C�'���4׆��F�&�����q��W�6b�V���
�,�N3V��U�(�`�zj�����\�_r5���WI�TKa�$їف�+��_~�5�Q<����n�����-��w�t���_��z甙e���#��� �����^��6 �����Ma݌�ZÚ�Ǚ�T3P�^%�c)	�V�����u��ӌ|ƿ
�2D�$�� ^�> �r#AO2�u�!��7�/̐�$ў��SP��iǻ���`haA �=���ã4�������dA[P_D�_Z\bm3hR���|]<~����ϵV�e� �>~]T&P���$A�K��`��ԭ
� ��f4�%f��i�v�i$�3���R��\��h,&Z�8ј�͡C��uH�aD�'=�wi�����ޣv�i�_�A����3�G@��������6(|3~��Ǭ��K�ؚU�fhE41eZ�I@`�v@|�u�Ia�]�K�0K���Eǋ�^�a͉�Ւ�C:X�u�C��ͻ*���ؗ�$c��o�8�q�7?ztv�`@G��ۥ�7�Ԟۡ�cHyd���Fl�?�M��ܚ�5)@���z��i��Yn�8��\i�!���/��o-l��J� W
�� �	�f��8�%ƃ+��"���)�-h~%������5о,�	��i��stth�Y?]tो����Oݬ/ �K�K����wNhBŀ�G:��$r�pU�m��q���E�̊����>�>(�Ѧi�۟�j��k���hF�\�^�d�
��ߋn3��(}�%����������$ܔ���Kd�����OG���RX0�&bC07�� `����8�f�I�9��-���?�{A�Z˂�j '�����T�n�l0È�^5�zU-��2��_k^�-*�_��@.0��'಺�y]����b
zQ�g��!z3����m�rV���E-qb���Dfl��HWԥ�vY�,�$#������~�3b���Q�øn��C�|�"���6�녈�=��P��U�in.� �\	4Uٛ���H���,�0 � R⓫˞\ �L���j~��p�W�iH洞�b,��8M0��4�!��̜�����:����g\D�h���Q��H�O=�u��I�W���n>��eEk�o}�4g xF3�э�I״�W��	�4�ӑ˨��>8�E�M��$�|3����d3g\��6q���7��r�޴A�BD���+̝a[�w���Z��d��	#D��(�����n�[�Q<��|.y��P�vM�  v-,� ��<O+��
3���VCyq�:a�ܼ�. ���(��'O��VЂ��G�Y��u�Y��F���-�������j��Aa�֔]G�t���0e��id�h`�#�k߷q	��I��0�k��4tU��L�4�����z� �9Q�#@B)i���>��	�ϯ���h������.~}���0��Zh�s��	i�`9wB�A�B��<|P���u�!E�p�YUH'B7hh���j��ˮ�c�2�rt�&Yi�4�WN�p+�S�-0�	.xnF3�<��[�>M��=�͏xz&)�2�\��2�vF��6��ocv7Ut�{�̾(7&}�)��L䮏%s��(P��5�,�A`��I�?�9H�m��� ���x%П�Au�o}�ڝ���ӯ�kf�'�i�<�Hk�ЮP1l�$Zl1 �v�\��v�H9_�`I��d��P~2> 8h�eȭ����Ǐ� �o&4t�zhM}���q��6�zZ������5�<Ht��=$��έ3 ����@��ˠLk�DǕk�4��X	�t2������H�=�}`�p�����֍�kiz�.�l:��;w�}��+4��ܜ�\�]��(Ȣ���C���D�v^t|��J�� s �#�2a�C���t�.X�6��� ��B�C]/_ۮJ�>M9y�;>}QPH���ҧ�|��5��0?�>3�WN�<G֞�����hF7E�����%�$����_Q2�&?�� 5GL	F�D�Ϗ��6��>��W�6���Zo��������[6_��c�En�;WQʏ�X��f�a#�'��3��S0Ϧ@�L�d�7"�z��(�4�ڱ���p:aN�&Z��FA=8<�ã#Z1��޽���?���Pi��n�����h�W�^��=>F_4���D+����}�9�yM���,&%�i֠i�	�W���������Xj7�ٜpƚF�1Dh�Z��c�c��l��D
�A��7���s$�ĸ@A�80XD9A�?�o�Y֦�����������2&�H �s�_�`&9zmTJ�BIj�A��^@]�&�bh�Ӧ�RO��XGƘy��}��WR�[4�e��W���ehM0� .ѵ1�%@����j-�om��K>[���{�6����e�+>ʍ�UƁ\
U�>]��I��o�u��7}��Imq� �N�㞛�+�I/,����$�ьn�d���
]X�����D�+B&�eZ�� �1W�\�i6ʘ�2S���j '��j��O��c��{5�u���|�D���5�Ή�$�8���`'�%�J�@}ү$�4@H������#�� `�жtisc��/-2�f�V37�n��Y\��I�ƊF�S�ɕoyoU p�&�ƺn���|�lyFU�����������۷�����B�D���r_�W,9��z'V5�YA2.���q�D���}�-�� XƝX������}al�洽DyM����(Z�5Й���U=��1��jg�� �����-C��I (�K�gI�}l}�Xu[��|sX|�v TQ?�`��F�%}�\�+O�������chaՂ6Kt�i���)�|�~�2~��7_������?p�GWxTv�$r�E�ve�3 <���FI!av�RB>���q��ۤo]���$�U6�i6(���Iur���3�|��B�%�0�̴��(�ˬ�Ƨ�Z��.�+2�@��q�>aJX�8���yD�_<���Cz��477o��e���$�ET6��$��*���Dy͆�5i�]@[�� ��&^�ͺܓ�c�'��l����G��ꛒ!�0��X����,���Z�Xͯ��%9��K�t�o�&�y-�D�����i?yۤ�[�:�D�N�!��y��2��.����Ǟ={ƚ` 9 E��B��H�'\������u�_�u��"�n��sK���<��G,R�}�f�<w��:�b���v��i���2�X���"`��>��a���|U��w]��D�����{����3 <�����*%�Y���
��<�GG7'��2�:��U�*�����<SG�����K`��j-�����
�U��yͱ�ҹZ�4�����W����p�� �>�j5I4�b����M��Zg��g��h3r�x4.���9�f��:��I����&<2�>-�� ��^�mR&A��z�f^l�����_{g�pӖ�o1��$y�ƒ{��	��A�-p�;g�Cn)$���-�lw�	,�ˑ+ �j�����wƌ�[Z����_����_>��w�XP+�t}��p��L��Q&��x%)��[�[V�o��n �2�a�@{�D�F;$O��?�"
�c�}�>��3�}�pS>��gR۫����o/��Y�X�L]�>��u����]_t� �hF3�dȂ^�|y͓M%Yha�YŜ�c"����|`qZ�nYyӞ�DU7l7(����$�6�ˀ� ��� ���&L�5Ui9;/-�$Tӥ c� ��{ai����)�������o�T~s�niS����F����IoG��"AG��T3pZ���e׌�\�j��Pi�.2��:�91����������~@g�g���8�7G'O@N����q.);|D��~��rL|��c�e|�9�)��R�`N>|��6779]!�=b (>� �ŵ���~�6��s[�_�/7�V���g�C���vw��M�$��1?��������x]-��[Y/���:Wl���k���W��lٴ�HA˴Ⱦ�u��� �ьft�$<�5��(�@��ƌ�j�6#��_�Q*�_���nR$0J�J9~u4%�^䔋�p�P����R`N8���5�/���^¬��� ߵ�5���'��gO���л�w�q�3hg����P�8)�>�{^���mN+߮���j����D���6ż.B���)lӼ����[�Z������Pm���FL��^�m��,���%f�9Z`��/�I��)�ఀ"/�]M<�n�����M*��[����(\~O�:�u>� ��� �A�Ч���}�y�_�����U�_	<�
~t;o���I@.@,�.��� ��[k��7 �@>���~�o������4�����-��T~\���,o0m�����9������<� ��f4��8s��ϕP�qn�sVs�<��4�-���Iz�`�e�\FqR���) ,�0��̄�IDI]�*���Lx.�$q�}�軖� �o����I�t�6�p�^���6ϱ����ۧ?���lv�
��.krM�w���E	c�� ���h��Z�ZW�����Lc-���/�?��?h`�x~�� (�ԓ@U����C&�Ʊho���ǎ�(e��� ����@4�
kK�<o!�t�����t>!��b�!����|q.z\h����I.N���L�/B"��� ���ұ� � ��)���4  @"�)1R�H )��Ԃ�~}sG��X�C[�.����6Z|@?R'����?��?��>��R��h�MZ��Y�]����b,'X��cZ�	��89��hF��%��,��j��|�M�~�V��n���UlD�<�Dk�\p��=>�1�
&o�ya���?��2�Qd�Ϲ�m�\�jt�O(���4��T% .�l��٣4�/R�� �폈,� ��N��8�|�<_jV���%�L$.����+���8�(�2��������n�YO^#�V�X����5[�6��l����>r�w��9⻮@�o<������=5���g�0��E���Lۛ	Rl�����Ќ��0Q-4 ���S�B�)��Uq��9���!ũ@E�����vw
<�����i��"��P�Pŭ����+ө�e��zlB��&���f@Ë9�y*��B8�Wh%�3H��^DXpT�>�.RW�M&h����X����������=�=i<\��W�a�TI(= տ/#ę����ơ�7�"U����hF����z�J����X0��-�2�B{����ڴ��M�
Db�ېݾ�H����Z�2�!���'~� ��3k՚u��X�fR��;������0��V��*����w0��$�����F�Z݀l�Q�ވj�&��zC��Q�q�搅A��6�~o� �4XKH�9k�/f��eH'I���a<���L@"��G��v�l�U�Z��
(\�V�:k�X
�q��kc_�|��53���r���u �H��ۚ�42c`0�(�b~�`7J����]S7�Ȏ�^� Hi��ب�w��c �g��F��ɩ��u�1ޠzh5qSq��U���-�OP��yg۫�|�ٖ�O��������9�\W3ꂧ��'?�����M^+�:S�_���<7��G�~�m��FK�K<Np^�*�����}�#G�:�$���O�^?���c5¡��i`8�X��گ�����0�o�UU��{ݴy���x�]ׄ� �$afU�s��~���H�\���hF�a��6����x�n� ��۝1�"@t7"lڐ�#XL�į�j]}�a��A�a������=oZ��iiu�����5	D��}z��h<٦��#T�O�g<d�Ҩ��iP��b�u~�c���j�-(Y�=f�����)��٠6��j��!
纑1�MI°Cb}�آ,I�"�U'`�:y' ɫ�W^��scPWr4c��(�ܣ5��[ ��Oo�}z�
3�/u�ur?���v�{���k�Y{���}���߬��aϬ�Cj��4�5��cj~�I�m�:l6܃�d���Р�n�g�tpxD�^���w��8
�ڀ����8�'�s�5."�q�����@�IOи\/��f��lm��dp9����n	��X��8�.����`����CG�G,�� U��H� ��}��H�^��`>�6K�c�
#�|�������mE@\��6�M���#�ϟ�5�ƫ�oV,T�>ޭ� �ь>*���a$�A��j�C�n�vv�5�-fl��1���6m�R�w�ү~�+�Y��kz*J^]0���)��T.�e\TSQ�n�����y�iC�$ȉg����:��� ֑i���\�����_�������}��"����s݌�v{� ���ئ�o6���״m����A��?3'�cI����$��S@���LCz� X��*cb]�da��P� x}��$i�f<u{��:� ��z�R,ϏR�� ez�h`ւF�V�:t�ުYo��ޝE�c�Whh4�lU1������6����g�i�����k�4�x0�����:�, �r9�E��ӥ��X�@ =���i!��-��f�u���O\�- ���{�_@P���K�QW @ ?��7����{��  ���^ ���ׯ�8�����E��&i-�����t��ǵp�T?7����4�% �H XV��g���c��3�?3��3<����ŕ,����~�#�N�/�p?Vs3d����Qza�ׅ�3��œn5��A�4��43���0
�Z<h�����<LkʹI��$�~�d�Uf
V���E���EӘݗ�C�Zr�/&҆��f�-��ܡǏ��Çw#w�V���gڎ@G�t�jt���_0@�M�5z�v���Oh���N��h��k[���ũ���MZ@|� �5��^ �7��m~A�$��\%�b�ڨ� ׬?� \K8	#n֟Ĕ7�<C�%�f�WJ�� F��О�ۛ���B�`k݇�2>����`xk�R���B������
}��.��-��W��Z\Zdc�ߥ!k�k��g���u�1�Zn��N2�Nm�� �%��5����A����~�oߵ�9}�]_�g�@@�s|�Xյ��>=�t�7�@#*4�Am郿�	 t��1�O�+ў�n��)h~�<y�p��Xx�k�\����"`wϑ�9�O�w�HٵB.vA�o)ߞ�y�<w���A����_�ɥ}�14	S��B
<�O�돘��a�g,�l�9dm ��x��V��1I� 18:u��Q�7��
H�^<��� �f	�՚.}��5�J��hS-z�4��I��e�ꙕ8���5��qu���Fs�Y}��������~D�.��rӼC)"6��X�?p�@F�Ꝑ�����%=�|��n�ӳ�����?��^�ꍆ�>p�� ��� ���Z�$ �b����<���j��+NMl�{����)&&����u �}�C�gFa�S � �3��Rc�v���ʆ���A
v�F�� +AN�Y��ږ�:V ��U�ܺ�9g�W=��\HOޣ��ǯ�_=�k����2��ʁ@	@y�ϭ7�Q��tg�A����={k�mz�*0@��)2kr��1���E��B�p@��y=���O���v�WZ #뭬�hA�o�ʺ*u�����"'j|�=L@0�����O��� ��b�a��	}!� �v���l��O���>� q�b=�?H�}���z�|���|&`�|TfQ3X���_�	��=��	� ߭�� �(;��[��KW4�s����xaUMg䣘Ҩ8�po�`y	)}�o �=�A@�aHy�G��Q�TG� )Gݚ��"��:�5=
���޹��X�czr͝�ѫ*)�rn�w&�(ҾĢ�
���L�=�^�N�3�˟r�;�y��A��!u�����������봲3�!�g���2P���� �h��&ͷ��/��:G+���mq�I'G�4�і��k�i �����rT�>�E�2&����7�8ѐ�jH�^�W�!B3(�PPs�q䔟�# ��P�&¹�'�U^p�EEC�m��K����%�O@��c�f̘�yWޡo~i�׿|F_}i��JӀ_b��(���U���C^Z�{0
��nН�9Z]�������NC.����3���&�K�^u�3�q��^����ߕ�sg�4H�FI�+���a���H�M�A�8 �8��H�Ʒ�G	dw��x���`Z_�|�6���mH�/�����_'�k�q�IUڗ[-��׍��^�Q��+ۗ'	�'���_=���3 �3�t3���dݷ��W��@}W����NxwS��J����0��� #.|E�	�	W�J�Ö1�[�(53�b�ܨ{g|Qt4÷��ķ��LB\�f�sS"i�2I�.��&3qʳW��ʷ��^�Ʒ��� ���_� *"pq�e����,/-����)���_������`�S��Ā�3Hn��1m���2�(j�2��Ŵ(��2n��b������6�1���<�ӳsP:�;�Tc-���
���A��Fq�|QW˘,!�+^*�RG��<������.��H]�d��I�ȾGG�'Y0$�F��Hq& ۶=N���J�s�,�E�X���4���/�,�j �1�,���K��o>�/��17���9�6 �}S|D��}p��h��Ԭ���Ֆ�O��j��ɹ"Hv�����W8p,�(�9�(YMm>ʸ�����2�������x4���q��'ÑS�*O��	`�S�0
��u�?h ?�@��"}��g����"��T@�$�c"�|wvv�������_�>��Kޑ��t�hM˭7���cB��t��\���'�����WF*f����³�s�]2�f �S��1��!�c�N���	W�yX�{Z*�Nw��r#t]�3ɘ�>>��2mP,���h!�ߏ捲w���<��@��7.�Bbr��R���ۥ)��fM��"�T�/�0v)�t��K��Qs/R��4܈�>f࢚ߪ������>��2��~}�����
��M�Ʋ�%s���tگQq�$�/��\�I+�K��[�o~���z�Nw�jT��09��Q��m^�0�[@đ�REr �kˀ���<}�p�~����;���9��k�\F�cj�*5-�3f?5�T��(ן#����ݕ��t&%=%��;H��̰1�~�k�g�̏U����봶-e�b�a����Ӳd�I����H�������~Z���L;���
8FC�Ū�����~��Ǭ�]�3��p�60�q��`��"$A�#X�����s4�ߡ��@22�i��KŤ�`Z�}ΝI���c֌����r����o����@��@��ȫPnQ�R2Gs��%�0�>;;��[[,�A�C	()����e��QA�`k\ ���}?ҿb�0�_�-y~�
~��r��:J�^�n����+e �I[	H?�c��{����\�{��|��q����w��]R�c[�wN��ƹ� ��ilى�0�h� N���;�4����Z�Ϧ�E�*Y�".]�.C>)�;����]�V��{�@��@E�Ẁ�?�m�:'n��!-��E$@V�?�j3QJ�� �P,��O�%��-����orL8�K����ːo|���H�������}��U��
��9����2O��.���{�(�cv�������'�8�aܣ_�hZ_��`Hw�,��_N�����twf��N���X��%vu^C.kl�?������a��g#��h�֤?���/!m�ۦ�]�(�Kvq���Bq�4f봤�W��뮱E��I�d?�/Ps;��ŶpxceP��R�ܗi�6-H�[�܋���q�ޣ+�}��/bik<V/.��d�H/��Q�ǛݟkG�����S�B�C{]X@�5�t���u~�	��R���1�{]�̠��!�Љ���ߘp�e��=��vz�z�F�Ю�o���\ۢ�3��x��K�(W��[��B���O$}��{��7���	�������s�\L�|�ˈ_	�4X�1h����:s�776���7��,�/�,//3�� �ZH�-�t�Ջ��s5|nn��]��Y���F�h����f�����AE}y��s�.�sF,ܱ����A�ۿ����A4���G_4�(W[�I��f�Ϟ=�W�_�����O�
�@5�k��ng ��D)��	��pԅ�O	�����4��Q��`gʚY�ۈ`��EJ;�E��(�+e��R&�� $��0#��NF�ޕ8_�
q�%���P������1wu�U��N^�bs5�0�P��)�M<.�߄��	��
���h���f�q{�9Z� L�t9em��~��}@���ck�hJ]�L �$#�s�c���	k��4o�u��u��ڡv+�A�g�Ч�fu��(�AoH�����Y�Q��ap�-���X6k�����Ԭ/ѣ�{tt�N��Wi{g���tޅYg�	���(`ag �M�&���"Jw�D0+~�: ����
K���a�;��d����i=<�haY��� �7=i��#����Y���=��8}�߅�i�zo�VH �>V c����;�!�\�2kaތ�����/���/��J̜Ck�<2@��7���!�4��u�k�fٱ�[�o��1G�V�x���-�=8��������F
����UgQ�5x�Ѵ�5�h�������Ʈ��"0q]46��gs��a
 >� 4n��p~K�`��Z����'$�4E��~_@DWC+_|��u��}���G+�`��sT��h��q"sC�=_\К^CA�;�9C��>}������ܸ�X�u(S�`��t�T�9�yx������"�^;�?;���@G�]r~[��I@�$��'��m��l�;t�,RKˈh��_��X��K��䢩�D���aD�� �:�~�< !��>&��S��|��;1W�K�&����|igg�	�(�
ۻbUF�gfR	��9��A��fm,����>���C�M8�O5�}c#��[ɚ�
#��8�Y ~�i�E��0k�"=0 ��
R��P-�т�8�^?2�)mn��I��V�IK���,����ԨQ����3���-.4������}d֔m:�S�i~��	�2d_��G�6k?�� )>��Zm61 ��������+��i=���ƈ�M^��̛ �8��%�&�����$ѡ��nvή��ۏm���H[��7���:���7��~����?�C3lL?�1����Z�?O_~��c�	Kw�N+���֨Q� g��o���7�t|2` �0צ��y���f��f�Ce'>�CN������$��ks���1V��Y?���If�h���!�Jec��:*���4�e�xь�k�E��"4v�+_@t��mF*�0XD*<I��~�V��Q�ݘ.��l>�b`�`[�E4��'�cq@��X__g��]@�4��MR���:H�S�X_y�r�^S�׮I�B��s����-{H��ੑ����^,�:J{$���4�?K��&�kDڙnP~�Y�%���Dy���G��>n�$��~��)/^ �:/��/��2�X� ���0����dQ��d�R\����f�]O�5��Á5���Ʉ��ʌ��{0}3�0���ə����HC���5���ɍ�K5���1l|�`S'���㿜ie*�񉐫���H�s��s����]>(H�.J�Z�U#>�~aa�VWc�B�K�	N >�a=�8m��ـv��hs�^�9��.��j5��ڣ� ����P��®IAhs�v�5���b@�=�?��(2(��f ,ѡ��63(����v�Ƙޫg.�����LH�����B�$�2V�؎M����R��^�X���Q1��[&��4K�'+���CG+��[7-��p
E}�-�cW����n�����H�0��t�y��ԤG�l.��;�@UCN��76?�����sd��� �j���#����)��-�6"u�sP�a��IA �����j ��ʼ�`Z#��MO.HPk5����[���?- ֚�Tc�HWF�
������O0����-��8mNݞ9�7� ���B�r���b1o�1 �9=;e�E��:xG�+�v�w�Ѥn�{����(�� �;.}V
nZ:wN��#�|ɑfcG �ܧ�`��� |�ܹ�� 0�;��֤i���B�.&r����h�N�M2�_�ۘ�Rpc��ew��(�� ��l
�+��������s����ڱ��`|��2��d�E,�0�`<f 8i���O�|��5�f���38�)I�L>�?��b�#��)�W�r ��������j@d�/\�D��#��c�';���\�<Gr;��]ݔD�*��1�!�j�@pqi�0�4o G08�h�c�����!m����.ml��L\���?$j����Օ� BP�pd�y��t��s ߥ�S��-v ����	��?��r{�wr�*���OP�Z�y"�˫�v��Yʨc|���n�by+��h@��x�줘�G����k��>y����y����;���i��|��kt�4|�C�������~��~|�I/_�����λ����3���3�Βk5������	�f� \��ԞC
�y3n�<i�#P�^F�;�j�j���z=>��H� ��i�����Tx2�h��X�<f2��l� L�h�EYI���!zxπ)�f A⢆�"�̝a��oh}ES]�meFWC���~^�|�Q�!(����}���4��Ѝ�	<8rq���ѻ�w�������~��.��»����bg������/$���-��:�k�l��<xH��v�â�O�Db� �}V�o��},�� xs�`�$ڥ���w�>k�=|Dg�6�����sk�d�A����˴$f�̳�����<��ŉ0"H�"i�Q��|Y���a�׾p��q~L�o�,�c{ft�H֗��Y�s13���2��Ɋ�5�Ȱ��f�|�]����7��'��N���7`d��N����cz��#�vYY96�a��� ���9��Ç��Wh��gf&���A�����_��06���NS�\��^06կ�[�_�|I�@1N�.'���T�J�r�J�Ea"+��)��5P�S��[���W�j����3bL2瓖k����(�6�[�6l�/�>��G��9�{�@���>4��F�,���.�͛q�?���bM�;���K[;Gl}ګ�`��V׀�s��m�?�������5�sb����=�m>sf,�Y?Iۂ�ׅ�5���	a�cʴ�zo���em>]�.Z۪�-Ӿ.�Vf> ��. ��b�qM��0@��q|��2�������Y����y�]Sh}�D�O���ٔ�㜌�y�'�. �� ����&��˥�.�y_T��_��Ec�ҝ/�c��3ow�P�w�]L��DY>"@�ih}ͻ���[�,h�����F��_��~܋����
Pf�A�{�{d�?q�l���R&@|M���b슔H$}������}��K|�ki!_��MCb��F=���7��OÀ L+?7�Q?���/���~aA������k��㞐r���l_��)�]]]1}sJ˦޼��I�DQ�O�/�0lj��J��iD<Ϧ��D3�ѧG.���bAlJ�I�&�%�@�gyu����#��YJ8���&L"q���x(���~�PQr�<�Z� �����s|�O���0&���Q�o Lc����1}��*�Esb�, fm4�k�J��y�0(���y��OK�/�����nV�k�0rv3a�9yw�7D�JAG��!�[JA���"S����P�5��m.0�<��r��-#��ܞ=�-�/Ҳ1^V�W���Z��B�M~����W���i�]���0g�T|D磐�&Q4�TZ�!�k�=Po`�ЀSF0
9���ӝ�ݿ�43��  ���3c�N�V�ZmN�=<@��^.e���[��uz΂\�ȏU�q������*�R���A>M�n�>'|���1���Ȕ(�0E�&���X�i���`��G���ן2������������*�߽k��e�7���@�I��s��L�]aDU��^��n�}:���w�[EcvS%��/�LHS�?�%�����w��?��O�sC�������w�}G�~�-�>c��%�74 ϵ�k� �LH��<9"ر��_^�4�ǜh*�g'�k�;0#�/���E�L�c��Bz�������%1;�Z ��lH&a�_dh��d<2�v��=0籑���ԊM�>{ �.,���|N~`ƺ��=�1`s@��ٽ�b� �n0xl��m����i-8���,����)s�M��L2b5��2��p�$�b�ӌ>q�.�e��|��|���eZ"����Lab/æ���!@�ՌE�gH?c�'�.M8[�U�@�a�M��
�L�+b+v4��G9_�$"036adׇК�őM�I^�:pz�(EÁ�c��z�zKgZ3�Gp�7���$ۍ�}'J5�j��wgZB>�AD�`׻�qݸ���Z�ȥ/J�x�䎖��E�l?��_������`��� 0�On����\��z��Je���@-���;��g4J�%�3�c.P�K���r�>C�Z���j�]K�B͐W[�4��3|�uYE ��h�竿6��O=�7-����0�7����O���oC�&���@��E�������������p�>d�H�����<es�&\b�!=/2N|c�"�J�T�}��-����^�_�d����M���+�����?�I����͚_(�~7����Z!� �'O*� ���D�J�g�8c�M�nq�p�Y6 H#	��놆�4W���%ɠM�y˄v�QgM+��j"5�|����"$M �b�Ii�C6'r`���ߣ����_����yvv����'�����������uf��lh��o
0�
`Z�駬��ҿ�1�Q�EA�K��|��[�ϋF�5�6uR(�`��i4t�3|',\��1;7"QU��0��8��O�n�g�}���藮�G��9�H�I�u�P>
t2�� �g� "䅙7��1��$P����&�ㆭ��5�d<aX�/�����-h����D>uHtӢF�α6�_����ӋW{�  �"�}E�\�S�?���f��Q����DkT��,"��n�ѫ��<�<�ٍ��v�K�I`r��j�W�
x�+Q����~v 䯍�;m H�
���/@ʛ7o�ݻΟ�=���L���w�̘��E�=Y�_��>�Y	y��H�!�/8 a� ��р���wY\FE�Ӫ`�}u��Q�7c�1wךf�'::>���S����Q X�'�̥8	x&@����h�yS\� ����i�5`�|�"��.�y�>�:��s���6����*���k7�R�[4����� E�����1 ]	�$�W~��͘�7,lͳ�����Y�Э ��E ��8�}k�hfA�+�eǨ���/���ӧO�_��_�o��� �'�����߳���d�/�/�#L��>���O�3 �3�|���D۞_�$Zf}�0,�S�!/�A�I��j� �����A'#��Q�D�j�!����B�RI\tY�����m��t�'��R�9� �8�$�/,�-vT`��a�����f���f4�AC���x�ʦ��1w�g��Q&��a\\�W �6mp���"9�jF���;�S�w��{�{F�6���������l�D���`W '5D*"�*r~��|�#��6�����lHp��`0�t|:��#���F`�!�ɼY��3��g��$^[!D�wG$�����A�~����\3�:�)�z���0����C�[�v��������W��ڔ\0���K��K��� 5��+J8���~���L��='�Oʑ�"��n(5� :��I1��xo���.E��@�~zI�'�4��0��O�Վi�~��@/�EԬ/S�f�k`E��?sf�ܿ�b�L�OL��l��4�:mNqtou�SnAP
Mo�4�֘3�An�g�U���Y��p5������'�P"zg�:^�]k�����i�� Y�-���@�E �쑁Bܾ�I�h���릟r� ^h��O�/� �Qo�V"lI����6!I���_�0�����?�H�nY���A{�w	���W_�����#���X�9=@����w�ހ�w�ޱ����������-�i�g4F�'p�����"eFh��">�[d��3Ȋl�J(9����G������INEѪ5x�.�dWLY�� �`���ٳ紷��Nh|�,���[��l�{�{��#G&+�p�%�!3�0�Ib��7u��w��uM?Fؼ����:�%�?�Tb�R�]M�����Q,Გ�s]��L�;����7Y#QI&c9�
�{�9x;�Eq��h{{�]2z�9j�1@~�~��0㭍8z��?��Y�޼�5@��Z�v�F�u�w������\���R$0 �^k@ܧ��}z�f�� �~��ԧn��,%�[M:>:����t�1�sg��&�.-��-A��#1����P�[�$�R�%XU�&��9	x��YTy�)e �ސ��KI������ �̅:�_m�۠��8:����[�ƈNN`m5�/?�CwV�>���G���ڥ�}�d͌)�-5�m�kP�Q�53��<X5 yɌ�����"6˯�[o-���F�0@)̙��v}�D�FZ��e��6�uǮ�a�:�y�>�Y�����C�;��O��-x�u�M��&�@��!�x)��o�Z����5u�D $���$��6��s淎��c!m�c&�>���*L�5�t�z�&�(k!�����������?�{!L�����gcc�-&�o[R���ϊ�2�3 �)��<�N(1+d�šA����$e�M�B%��T���:[�DjD��6���"*��)"����ǾRY�?Rǲ&T�ܓ]O�͙Lrfͦ��bs-h�9��&>H�t||����(H�����A����ˬ��0��FH��yom�=�0�`��Ijz繛R��T�� ����A�M��;r�
2*P��x�k2���|�{�'C�я�P�~I4�ZU�X�03��c9��������㐎,��Yk�u��e;�����/����0�� ��v���ԡՕ�?u���a��s�5:;���{�]إ���OL��V�zԭ�}������̈d_��o�f<&���t������jy'<Ki{���z��}|o��:ż�H�l�zzb3+�s��TD!��u�=?�ha�e �.=�צ��<u�5��z��f@�V�A����" x��"�7�SF�X�!�~݌e\�3n�tx��=`����vڤ}�O�U�7����li�[�3���-��{] ,�5��{䢏lզ�B>���(j�R�Dѵ�Z�?>��#��/2���_]���TPݿc�<�Rv ��=b�|��|���` ݝ�mx��.4��&p]�d�����e��/�}��_�f ��'g�����B�p9̀�ͨh��sw�~��Kw[fS�s�*�Պg�*J�Y1���4֚�إ������:>�/���!$��r����aZ3�Z�2�T��.3���$���u�D��S�l��Ȯ�&i;+���лH��Vh}m�=�d�K��%�N��'/+ 	�u/G��C��}�}��Nφ������xCg��Z��j1��0�.F���*3���>����GsZ�y��@}���K����0�/�U}4�isk�v ~�r�#�=6�FC^{���.�b'��~<���Y ր[	�?�����6}ppF[���;0�[�<;d�Mh��dO�oh���S�U�}Jo���2`-w�c�`Xb�{��w��z�֡w�!n��(�3���kB�ۢ����y�n�k��nR�Qc�j�/�wGT��ѣ�yFoD;;������:�Ok9�g��όn��Hk���.�}����}�Y�ύ�]$��\'T�-��
]�9e_���T�����~���ӯ~�+6y��Z~D��7�1[8Q������b�3@�5�g<��hק� ��)�j�^�x���(���p���gq�M_~q��~�Ns��a�l4PD�)���X�\�,x�Z㐁e�j�y��>aM��i�����=�T;V}�*�t����<�f�%� ���O/1)�K�q̻�1}9d���Ľ�-,>f�}����<}��=���ӝՆad���L?!�7Ƃ��7�7L��w��2�d@�=f��m���%�l�U.h[��s|Ӄ��`4�~��6��c��3��^�b�͛-zp�C��-Ҽ�A���H�tF�ύ�Mo�l�٘���+슆���|o��D=s��z�j�������Sq�.HA�@e��:�+�.�Ik?�ع�ן����D�wm�OAE��M��p����g���g�{�G��}��DKM�@p@`��� �v+�V��{?L���&]�bN���_f������C�����ն����1����ȺybSSr�(lі-7(�O#Y��,+�=�c���'��r��4��W-d�i�%��GL�9��ڬ�:�X���+�,��+tJ�"�>#�3R�B��
M.��A�����r��K �PDAc�C_�L�gt	�iǉ�o�U��W�_�Q�M�Glep�,�eq���d���:��m���֡��F��4��&���j�)�ғ�^LV�Y��\4֚�^gf���`��4�T��C�7����a���:���2=�b���7i�op|�Rz~$y�D����K�|m��`�>G�~@;�]:<�r4�k'W�;�}r��uq���t���4eC��v�����@�]�N�IK����h�kn�sÚ'�56�0k㢄�B� �,s�A�:<9�������_�����X+ȆA��e�"�{VK`��l�p}��5U-I�$�W�H����/E����� �Z(��~-I�G�ֆm��n��|�Nא�a��jw]<�=æM�(L��̙�]�w6{dB�5[+�?�ѳ���~���i�vw��=�� ��
�H� �\��Dhͽ���=^ D��T\ׄ�狩S�M2�t�IyeW�Lן��g�㚁�4r�:]N�)�&__V���$Z�l�4���	4���Ox�G�/N�� �[�}=i u���qI���<��߾Msk�4���\�j�eD�F� Ҿ�Z3菂�b�5=.G9��bd�X�`��׮��B�l� �1K{!�e�0�	�����{�~\o�4��"$�-������q���>b�@Y�)-t�Qf~c#+�8�����D(f� �;b�� `8��bտ���E^�ns���	.���4#2?���]n�Xu����K	�� �>�p�h�����"�E�M�}Cj�a�����̷����D\v��	�*u����c/������u�����em��/*�{%�7i�|b���X+�KF��y�]��ݦ�f����+^s�~�F�f^�EsM�Lz���o���6�eD�� �_~�`�N�Zp~h�ɫ]��o���M��?��sô6C^?�t���8�d�4i3[�XUf�5#V4�q�5Y�l���/3�cЮ؅�s�bْt��
 [���3T{L��-ڻ҇��k˘T;�4 L|�ɺo�z[4���w���^�k��� ޿�U7��f#cr&��/�_��V���ev�y�=�ӫ7�_Ӌo��:3�+4�a��E��h���N3���5�o='iz������qC���>�.��T�������{X+n=����w|u��g�4Q܎0H�[F��=�=�^+}�K�Fh ��U2�.hi_�|��^���*��r��T4�Rg�=ヹ��䎫i�/h�o�nX�'�1p�&�9�vB�f�A�{��??���!E3�#�"& 8I+a��F	�5��}Ȑ��\[k���%�`���L�d�͙k6xS�3w7U��8��O�MG����.���`J3	��d!�ˤ�&��36�o��͏���~a�D�L?������m�c���e�a�H1期u�h��D�`�V7h��V�=FhMYU���4~��2s'W�kT)���i�:��z\�q�ĤLzv&�'a/����ʘݾ���:�Ra���2��'�GU�ۍhk{���_?���9�X~��Ǵ��B��V�5y#�wS�9X��L�����hJ��o��t������/�������]:5�%2u��)l���ȃ�1�#�&#ZE6�I��-#�'e��^'�W������&�'ҥkڱ�g$�Z���(st���;d}��(�)���ܜ,O�#����ֲ��(��3(��R����ptk�����,�a���;���_}MGg������A0Ř�>�7�7bW�8q���G&� B�6���~����/ikk�M�[�ql�X��ٻ��c5i�tl��L�>/�5��ej R���帠L�v�+��� �{)�\���Kr�"T�ˀ�"p��eW�GS�ه&�ZK*� �5���#�Y[θ�Ѡ�� 4�;�cS���Gf|Z�2� ���seh�u�*����q笀Z�`Z̨���
� ��҇��	����\�&��X�ٱi&����M�	"��F}b�'��Alˏ א����T��E#L����h|"�k����vc*q�DAƌ�o�f"��'	�̄f�H���ƨ��X�0̞'2�(.�@��#DY�����J�!���yW���a�����0D�� �=����ţ"���i��)���g��q�1�e$�i�FMb�o�Fy[h�ٔ{�Uh���r�2���"�X���"@��3+�����̑���u� �@��{�֬�pO���~D�ݥջ6�;�M���b=�!B�]���1�&bw�^��3��5={���p���e{�歃v�aR��m��D������S�Uƌ;d�xAZ.@�GoTZ>�s��S[�t������se�����쇭~��.����j�XOYw�Z�j���A��^'����W^L IȦ��� ��?�4`!H����f������I����9��A$x/��#$G��ß�_���v�kG(,K�LI)$qc��9���eUVe�T�{�$3�Guu]��̬�k��hb���oq�A��ڠGC�ʲ��w-��t:���ᔶw�Ӄ�_�O_!��s��ET�5NӇ�S�"A��l � �r,����e�\�崝ϯ��%WѶ��z�������A}:�Ч.�3.�sOB����^VN��7�6W�h~���xQ��: V��4G40.ʀ�vg{�ǵ ���e�����޲O�a�=<u�$dD�G���q뭮�!X�'�(am�B ��9�� �1�g�S�\���g�<�OEA`8k�a��f�O��*���4G��g�{'��Q��<X�!�T�eV�*��{�6�W�g�C�K���F�����|*,�\����
֖+��+���~�E�?_��t0�Ӳ��ԁ��t4��7�~O��Cw�M�ߺN�=�֌J<��ztp8��O���_�_�q �����z�|�^�ءQ�-�p��<�\79ShVkxeRnK�uS�"�|KM.ܵ���Ԛ�^!E_���d%�.kI��3@���M��NJj��	���CIp�ց���F�FR����L���s<r���s����������ߤw�IoݺF7��8��d�U9�v���'�?�}��cz�xρ�CWޘ��X)�+oJJ�ܒ�I�i�֩��R��'�%�Z�Ϩq,��GBI��f�,Y�  ��={� H[�`=+���� qQz�Mƞl�_(?=z���� u2���	��/?�J�@`1Q����u��fP��6u��vY{�c������ �Q����\�����4�@֪�I5#a������)0�����Ma`�0���Vկ(�,A��	�e�� X,��Qב(�W��ɞ��ɘ�%V!]V�PDu������3;�{��GS�-Jh!Wm�B%Lp]����xe�=:���U�y�gm�u�H	���6�k�͎����R��5����ҋ�mz�s@?<ݡ��[oߠ�k\� �t����pL?8�����g��r0������qx���������[-B�L�`�da���_��ױ\�b9�xIYぽd*������UU�l����5yi����J o����Ϩ�!X�����3
j�Ⱥ��.��V�C�Hm&����|���1M�@�����O��zo��z�&ݼ�I}�N�G#ޣ>�s0�v>|B��k��Gn|��q(V6�s���G���V
, ���$������&�Gn����.� @?��ݹs�#�jW�^6y�+�<�Ǒ�w�EV���Ǐy����z��ț�>-Y����Ҙl� �*#_���z_��GI��)�2�-���&]�!5\�/X�tJ�huiΏ)kCҊ[�qq��7�A"8ΙVIio�_�>MD��*� ��CM
���^�������ח�\H@<5J}���.��*b!��f�7�+��ӧ�]��;z�PP��~�ɶ��`��tB��;t�t�v�1 ��_����!m�8rtm�J�S���i��-u��#�!�@yl�����-�O��&�R�o{;��Bp���)��z�J��B���У-p���7��m��MU
��!�"�TV]W�m�U�w�5؊�vӚ�[QXv���DKt�{4�Y~�3�	{
H�YK�R~i �H����w� 9�x���/�4:~JϞ��_�yJ�67�:�a�w�s�h:�A��GGcV�����~u���pq���-�_�e��ǲ�?�. ��HyZ$�����������K��^!]���\�f����m���>}J�ӟ��͛�m �及����"�bI�� x���k������B#V掞�]��\��ʞ�2$�3��Q��fQ�gӞ\\'��U9/���堣^� V�UW�#������ƍ|�MC��l��yt���l0R���ƯL����fwuZO�h�s�I�Z�MF�n|����"�oU%w����Ӫ�j�k�-�H�wf��g�%=�j�s���ߙkNX�dU�*��n�N��U鼀�I�� ~A��\r�8���o�n`+Z�j�5r �9�Ǉ�r�������������j�?������1��Z�|�gvE�kg�S�m8Ae�U �g]7��� `m
�"H���,sA ��3U�Tޅ��di��D�&�ӆE�$ŀW��Z}P� f���U@����8�.ʦ��u�~<g�EYeeE �6F}LL"��o����"���v_�pcf�,[����9��|Z�����6��.�7�Q������f؟m���*�]:�UwYg�r�Y�r��3�J��w�@�>}��W���P�g%��}e�4�g���װ�~����?��ݠ�2ϊ|8�[���=O�䊤|^�{������(v>�����ﾧgϟq; K��i�����g������?���O�䞄��� ��3��&;XIÜ����+ݹX*u�t+D2�d�O��jO��TYyI�H��^�j��MVn��=�W���_ Yǔ��b��QYm^SZ֝銖�60|��7��ew$�=�,V��>����p[��1���O�������5'(��"�����#�'UՏ�z,���R�t�/��(mmH[[�N��M���\���|��A� |A"46���^�%^CZ���.��@�S����~��m T��d2UB�j ���ʼ~�:m�~`�`v<�ã�`�I X�ƾ-��U�����G\G��Qύ��?_�s:_�A�����$`�e >���ԏX܉�������<����VƲn�Mкx���_�eD�����}��=��ڈ{2��].ҖU| � ����?�����J����@A�es!^��PPŕ\��ڛ�b<t���~��G�/��/���?�����~�;���kr�uº��'����������7* �s����
 _��1!7�H)�3��6�H�	m>�&b�Iw�%���v��+����Wi���V�(�:k���+�i��<-��P2(k�ٓ��"ձ�Oq�v3~���-���h�Ņ��ai�y~�ӗ��nXm��a}�LH�<���g �J;Ñ�{!o9���எ�5�r��	��=[�k�̸����I3Z:��|���{�.����w�y����z�����L� �A�Fq-[��4a\��ا��rMX�l�O۬����>ڝQ �/@F�������-���o�O>��n:�q��j~&�i� K�,�X�>��5D�p�EKX�;M�LUpg�!��A {!�[J-U����۱�YJ�߫(�Js������w�����c�������-��x��w�K�v�W�+:{*)�J}���7gX~�� �����>/���c�����Ǉ��W�y�i���I��Jjq��g,����~�� .�p��T�^X�1���/�����<�),��/,�/�!o�R軮 ��EW2��,l	�snI1�O�r`�EICbC�&y�h��g�&��e�^y�-B�:��	�΄3�?GŎ���C@��ٸzALS	#�<3����hS���F�b�M`�y\/���׼�"����Ezq������r�}I�X�m��"m��r�T�]�F&��秵�ޅk�0ν�!�U���~���� ��V�,.�(�O�\z��O����w?�O?��>�w���C3��X��0�7~�+��#��D,2�E�-hm�#-ϝ� י�6�Q�="������Z���<��+��5�/���/[>��o8����w���q?0�����Xݫ|� T'�vz�p�-� ~gEQ�[׍�^���C�X�^Jwm��"���6`:oݛ�����u ���o^^~���X���3ƾ����'��'���o�(I>Y7].�Wtv��RP>�eW��y���nާ��:O��e�M>W�r ��e���1r��])W"C�:���`���/E��^���eI����/����gk2��0x�A�Ҏ�9ZRdE��x�
 _����kR*�H�h�]��b9���D��#�r^�"��@�zHÝ*|�E[*A@,Ƥ��0�"���X�0Ԩ����/1�=�-�&dxF$�h#>���|�.-���C�y�[@�b���'y4�}��-fE��:���L�kM�������A~����.�����bo�x�Xe��_jF܇��ѦM��2� l@y��)}��Z[[�q���ϭ3e��t��|�6��K�*c=�P��ߦ&MO��QL�<����"�������H�\̩�J�{{��_~I���������Á��S!�����2al�� ��l'N+��X
������:%���y϶��s4�Y��G�y�mV�6�2J֧EH`� K�W  I Űc}��(晶��z@\�y�ȃ&�i�]���C�!�3�x�������|,��"����YD�Z��m�v��5t	|�9�����nܸ�c�����9hS\�� �\�!��\�������+ |EjB��HF�XRd�V~$c�������$N��^fA}:?+��}R� �Cz�#�!-Lᾮܜ�I���#����r#B�k?����?�۷��e~?����f�h����)܄|t�+�$��z�HG���}
�\��\�`5x����9f���^Kzݐ� |��yG�YZ���=m��7��'��{�_+�u���"��B�-�R��
 H
��ڂ#�swS�KŠW�z�Xs\�� -5�Y �Ixe";��8G����й���)��vm}-�f�5����oK�`a��R��c�j�+<T}�Qh�gڳԯzO���kk��G����Z+KJ�6�,cA�2����[z��[ʥ7o����k���Ξ��5
��_����J|K�'(1��XW��f_��# R,��/��%�_r�v��y��pux��׵�^�M�H�#��Z-�u\�'��bu5�.+��')g�L�Q��J����|n�M~�]�Ӡ8�U��` ��ݛ�$� F�X��~�6���]黩S��Z��P���?�ca��;[
�	��6���wߡ�w�V�m>{:�j��& X�N�pEݤ�P�\ =���8�d��`��X��� s�n
Q��3�s�
��^�,k�Ӝ�����N�{�nМ6.XFX�( `_��m ��]ip�+mi�I �+dOj8وl�5���[�� 5A#ڰ��Y�����Y���� �4�������끶��!��y�wLAR���6��LsY�v+լz��/SԪ�L� ei7#� ٣.���"�Lۨb�2ʨ����\/��Ѷ�� Y�O�s�����}�X�%]������IƉ(W���`���C��@M ���?W���e���sO�]di��{@���~i=�Õ�MM���p�����c��. ���y\h(��ꛢg�n��J��|�c�R��r�n.`8fs��!�I@��H�aO�b��	8�ަU�Ir#�V�^���!(ί�}���F�i>V,&����`�7�Ν;E��:9�L�-Wk����Sr|9�\�Z_L�9�1���]���2����ׯ�6�w����W��EL�?� T��1'��*/�vҷ�� u����2�$Bf��47���m�L>�q��2p�$i��/�����!�Sfaւs�� ������=�pqW{�QJIe�ۏ��3mXg����\����8��ZK���;�_i������ڿ�����Y����/����P�ʸ ��h��u�j�?_��Gm���J�	�\������U"ٟ��Z�`#�ۯ�k��</
�X�1����_�2�l��h8���\Ĥz]����[�LY��SkF_�,�֨��ҳ�ZI���GzBINJ
L-�BP�$I�!IT�߉�7�+sf��x4�u���\�����͘�)x���aEbN�*�Я�o�$�uEv&����y�F�/��b�b���u��s�V-T;� ��Q��<�벮��m'���6������J���mO���Ig0�tS����&"���)`H��� �F�M<�\K�b�=5��.k��
��[M���2e뀏>,��-!&(mg�L8���[l �P�͸ۉ%�HO��R�$�M������q�_ kkw�^r��p���F%5����~��s�b�F�`����n(>�"3*d�q��j�+{�,�a8Y��Ά�h�ln�k����̉�u�w��s�F斮Ӡ.�Y�˶Gb%��h��=��O��Ki��[p�~�[|K�V�'�N���!D���9S��Ϊ�ʆwsc�4��a��'O #�D#�� 0�?���m6���߿���|���gr �]�/�nܳX�΋��� ��e$�����e���|�5ZӂV,W�!ÿk�$�����H�b�8�9(� ���ۧU���
(�şt�/��֑#�P"��,�qьG��[+:��l�>�Cp�aAM暅��qM���h�=��d]�lTqj�=aa�FI��X7�Ҹ�:[r,i�{�$��¬5@� ���B���hcK�	��~T%P��D�ؼ�Q?(�*��>�f��v��o\��h.E9]����`�O�ߒ˶b�P��;r�����R��k
 ����֦�=3���EZ�����\�{�|���#*�^��&��/�g�EѤ}�X��[@��Ɓ���2Q�٢��,�Qd�֦v'I�d�c��u{�@Cu4�5�4���R'�8��q�2��)Y�[ ��hS�\��C%k�>&}%c6�^��|\P���<)�k�d��빾>w���9�]e�
ܜ���o��o|/r �|ٲ�F8�g�d5�����y�H�(�O�� �,�m���q��BK	���?o0G��L|���r��ڵ-'���0c��pDb���^AǴ�Jpt|�2&����zn�������U�ǻ,�jʌך��H�_�*Uhծ�Iݣ��;���N�2���ҋ�7�[՟����-���Iv��֖�z}���1�!�xA�do)ބ�����N�@i�����(.nb��| �&|��`-����,�7u���v�OU7ŹVki��^�,�D�'�-&P_�R�{�y�s���VeՅrцw=���YfI)I���l<�Ⱥe\�d- R��euť6*ո���K*SU~5�kw� ���Qx��i��k���N��/ky@����L�����&��|o��3�
ei�ղT��I�<
kOeIRW���K& ir[[��������&�o��:Y��;��&�]�o�F1�4s�jw��q g��-�|�6_om|'(.[-�����aж��9)�$T�eK�x�({�E"_���u�6�R
�����+)����'�o�5��h�#:��%� � `H���U��}�����G+T�,�;��+� do5ʇ9�]kA�+ �X*,Q�ڢ�-Z��g	�e���K,�y�N��Yyf2Xе�kt���t��t�ƍ�x(}�{�}2E:WN�g��r{��>|@/�?�	EIH#����j�ݿ�O ���[���es^�i�5K�)�Н�t����S[�2oKʲ&}�
�yM~[�I�0�F�%AրQP/�mM����)���M�0�7���%�	=�C��j�!��g*8����{��;��>>j�BԹ�_=��F�X	c�/�%�X��U)
 b��2�|ĹҼulp&tY��(6O��k���Ih�J	3�ur^}�qK�ys�(�v��23[@g_"�v#���+�x�)�U�<�\�P�������Ǘp�流'���Pc��ڰފ@!��؃4��x�~����-�.�[��v��]�Ƀ��"H��ǻ�	P�I*�� �T�V��4�)�s.�kN��	��>�c& ]�U�MH��C�Mz���_I[7�����`������x�TZD)o!�>Ԫ�l��a�.���y,�R�c:P��>����W�(�1�����\��SIA�
>G�uM+�����3�-R?m��1���L��K�f|$�b~������@�,[@�U\"d�C/�㋿�q�X��=�6�n��Ѕ��.Ah��KĴe�Q8ΒdCG#�W��ߢ䵷�nnl�[�ߢ{�>���SΫ���M�јzfvO�W�I=� �𚣽�#~�X����%	{K���G������Ѝ�ޡ��c��~L�0U�� |�zw/&�+p��@PQ���aP �x�ҍoݮm���x\[J8���h͋3�Q��6��O:κ�\N,��GJ�E��x����u�[XF5������N�p���Vj��`-F�Bo��8a����h��C�,��i(��f�r���RB�	��qS��$�)��G@Qh��첀�.���
v���y̿�|J�`m��/kU�v��� ��6*.m��]%�����jب���ɮ��f�iQ:ť5,c�W�.�����'P�ZxDY�^��"�z��n��݃F�*��j?�?�����?�,�j� $�:j]I<�"�P ��S�>���0�ٳG��s؛\I��B�!p*<�LlOÀ}F���i�!��ra��`��ѕ�~bC/�Qyp5%j��|�֨�#�v~�eX#�����=3j�\s��Db����.�� �6��,��<V�6�k�r���Lc� 5�iW��%:v�~���a_/"<#��E0ɗ,u��Ms*��R��1���[[{��h4JW��%�Dg!�{70o�G�zt@0��g��`� �޽���N?��g���ӗ�t��P��7�
�7{}l�Ys*���5�q�&���������|C��OXF�3�2Mܻ�iwoD�_9U����Y"���*���O��aK��� ʝO�h<��=��On�S��m�6������[���I�^�хb�.2k�������J9����c$eOi�pL/���:SO���6Z9�	�dy,a|M��0Sw��{p��ƨ�M�şJ,�Ya�5��"���V/��"�J�>�	�Ab��7i�{����'��|%���cI���@̋ʣ�/YR㺪�pu����
{S-���9��Ҳ@\�eh,�ta(��)D��-��V�h�-)G���^i���+�gJ1M u/
D����Ӭ���A�T�eg�Y��<�J�E`��(�*ͥ\ߗ��l�K~��_Y{/���"� t��&݇Z�=+��ג[�v,V^���tC$�n�"��x�OZ^`�� ��g�}F?��O�{���n'x?
HS���OZc'���8 0"��,M��߮��T��a/.@/��=,f�4"K=:�bp^,�����ݼ��@-B�:^'���@!!��:�	��Nm��`�������M���r��h�Gw����5�&�v����O��}�|��ʥٯc����W�~˖^Cp�ؠ��Kz��<y��1���IH��'��d[~K���Ղ�Ʉ����Y��pL�B��z�_�Դ�{Hx�Ɔ��O]�L��g� 8�Y	� m���7uo���ܢe\y�����txt��֗�G��ď�����Tb�9�t�9۾H X֢��[�����D���� �Y�e�7�<��j�V��% ����M9~��2NlHм�/���2yD��}*�o,J��X�m����冚�[&>@�W���,
�:0���q�X�h=��U������(3+D7�I��q�XB��@��G�aBv.G]��q��-8�^��Q	�.��h����ˌ���p�|@o���Wo�� XJ啞�I�fA�o�����石�4�_-�n9@�����s%�AJZ����[�良�2T�J*����6^@��&-N)�_Y ��X`�G7�4��䎎h�-�[[���I7��Ӻ���	���!��i����.^����v_���xB="w��L-�|��~�K_�uHFޙ�������Nh�]�7���b{ρ�}:v@ʷYpݒ�#��6>�*�2%�S��Dem�	�`R�=�Mp/YTA�4I(	��f��Gz����#����!FH��bU�<@��Űrc����v�i��� Dӥ�d��ĕ�����=�U���w	1������2�y�)������� 26�r��l�3n�ME�/����X�W&Sy���V	h& ~����?˭�TݸI�8��-����J6�@��LqZ'Y�mE1�sį��X@n���\_[�-�f,Ȅf�G��6����x��EzC,Q2!�C^���ιC~%��\�,�E p�� ��Ҽu �[�OB����/8� �֭[�[�k��I�!��<��͛l���m��H<@�!e.,��H�c]�r��l�噛ܥI��]rr�fa'��b�֒n��	M'#�66����No�ڢ�uD��0s��po�+���&��ޅ��`JGG���������3� vm��s���"q��A
��d+����"0V��su��iLc҂���:l��Y�&h�O�	d��Q�L�"��c�<3�Q��06���ǋ��Px�h{��w��vM�ʿ�����9"�Fѐ���{,g�GS�S<��۱^��9�u �ϗ@�nt���u�d6]v۩�����~����.�S4�-E!>�_o�{��g�+n�J�/
�P�H�xϭ���8�@��I9��������s�ZU�[:�hc�eb�MX{�}��;�!��̛ʹ��a
���eP�e�yw�SK�X~���#G�'�A|�gZ	��Z_�ԴW�� ���Hz��}�k�+��ߗa]���p�4MW@��H����湢��J��ӻ��+����osÎ����8��G"-�5:ER	�u�@�q�XE�'|$���W-c��`���Q����+�2���],�H��l������TN2��L�T[c��#@��v0�[��p�@�a�歭��QҼ�B�<L<7�8-λ��yB�^H�m�A񒃾/o�� ����X�O���zj���7��@sv��b7�E�Pk̂�T1�X����Ra�q��&�Y31�.���,���C�{<�Ǯ���c��`�QAAMK��R�M�:h�H�{�Z���=�~h��5�|����Tڳյ�k���sk�2$���x���g�;
g5��[0��y �דp�/��.���.ƕ�cpC�ϔ�ˢr�/�bmu���reh;���-D>�2�"a�Gf�!:�r\�K�N���h͠��(׎���
JJ�d�P���rA�Rn ����ި�n�yMl�/2�ݢ�U�g��b5�,��s���pe.�
<�s;� ���� _j� ��X����\������H�����l�m��ދ�dem�?�����Z���9��5���*��/ �J�� r�ui��-~�Ɵ�����v���%�4_��oٔ�0�H���T���9������}wm�@\"����窿� �[��IbErYup�"�.{��~�T����
;
�3栗��)U�
��˚�ݐsT`{Mx��h���V�E'30��k�b��MU�n�s�Ό�[	iRN��IO��rQE�	�z�ERZD��d����6� Hqڑm\�<��-GW���q;���.�!+㘶�[�JLfQW�+�N�,�5��s<�9��=]n߳U�v���E\���T9��g�+�{%�q��n�V����dm�aN���&&�)��l\���8�C����ϧ�r��,���V�	�$G1�Tl�c�a�5�q�_w�q����5S?D��ǒ���}2	16��8�,J�r�ٰ���Y�p���Q�&���`���,�Di�u޾�\<Ѻ�Ǵ%�9�s�<M���f!��Wy��_,����|~��]�gUZ kwfg6�%Y��w�|���<��E-�:p�@��v���K^�B'N�t^4�
��F���./��Ԟ�.�bBaq�y�f�Ȭ��z?�L��@H�:k�k���ݧ�����w_��A�Z�t�z�j�?����t��-z��w�t�v�� �4������1@4^aPy��x�'8/{}v�RniK�A�S�SNԑM
�$��Ca1
u��]�:&��u�1�(7�� u�QnJ�c�����k�hK)�,�ߖ�xAM�p4�A�\_J>7mi�R���˶����W��$�\�P�S��MI@cT/��E�VE�1K��I�mIj0�L}E��< <���	"�,��E�����x���^�X�����k�� ���>-Rr��^�mm���:�ߐ1 %N�gj�a��㽾�y ���X��2�˰��ځC(V�a�v٨�M��" ����1W�y@b���*�����(n�1e�4�I^6z��6p�-Vװ����գ`
��&g:�; ||<�-.GG#�R0�\X�Ŀ��`i�~�����pc�P<��)�J�p0O����+���R�]�����A� k�Uc0�� �]���������=J�k��s	�I��w���r\<*�R)�
{pۀi�@�nIg��(���y�U̗����_�6�z~��R�}�:���li�ր��vr�Rh����_�أ��^����$*��A2"Cpe������5�8n�ֵu�Аߟe��@�
 ��ܹ5'����������L�@%H/$	������Q�������G�1êDz0-`K��:#k� �
SO��"��%4�k���A�K�)��-�O�o�hcc脭M�v��6Q?����Q����ð[< rt<���}7�&�����V"��Mݳ�g���o�>t����۠���rח�eJ��y�X��יJ�U4�]}��W�W��3�{�Y@;�z���L�<�j�ܸF��6�u�]�6��!f'bA@�:e0Lbq�9t��j�Lu��O�������|��YX��0H�Rl��gD�4_&N4�z��Qa�~��q�j�Vy���5���7��{��߽E�7�Ɂ���o2�{㼫�i�͸��=pyH/����o��
cVf������sjuU�� [4 �zY�-�4y�=u_��j��)���횦 ����V(m]�眖��r�Ů{z��忒g�>w�/����t~�2ڮi �,��w>7��"Ts=Խm
�e(��%P[��́U�ua�׍V�։BI3(Z�O����ߵuh�hĩh�������5"�c�m�`w2�h$���֦o��h�>��c��Z�SA;�߈�]�F�w�n������J����s a��ې���� ���3�=���O_г�����3�,�[����LsX�9��}/u��h����Mz���t����gy�8	wyQ��%DQ�)�����i/^��Ç�\���`�!�.E{Y�1�|>c/0G�E4#0y��:Zʥ�T�E�{ e �_�`�ө
���4��㚜S�8X�\[YmǺ΁.Z?+*YC�q�;�׷苟}F���C�}{�6���t�>G�3
`���|�F�鎘�`��9��O������s����oh���G~߇UJT
 ���1�v�n
M��%,��|I��f<ѱ�qkktmk�>��}��_��>x��'Gn�� �N��Q�nV�|5tx����1����;�m�ww���tm�S�I��IJ��#�Ģ���]��V�b��~D��$ѱ<(�#!^2 �|ztY�`������$�sb���u�`j����.�OW��໢�|=/y�����e�v��6kn�b޽%*=[�X�Qgm�͕1�XzK���I��s��sĺ��WU
̣�,_m�����μ|��:yǔ&L�"������\XQ+<{�,��v�7�yǁ�5z��uZ_2���^#<	��ǎ��ݠ��ڢ���S\0���z<}%������AEם����w����9��gYH1���Aw� �!�Vy�9�)!@�&={qH�S��egw��Ga�7q 
����<5S>2M�wd�Q����H�����qr7��t��5������Oߥ[o��n�����=afv�F046'���	
���}��	=�M>����7G �^���[+��j*Y�=Nf�ߨ��L��K`�޶
���.����������*�(��<a�2Ϊ��1I�.[��;o���C�s��6�;w� ��	�������V�p���x ���`�&����uw�"/`�ح�G��cE1��K�X�7Q
/�
߸�4��~���b^س�s��ݿw�>��-��VZG0�uؒԬ�^��ֈ[��t�k�!|cMƴ�/����%����FA�a��L�
.�f�"�9H�����~�&���z�E}�$�
�e���a�9���/ �V���k�*F�+:}j㷹�O�����Z#[�L��z��L]c\ϋ�zپ�c�U:W��:��1߉fe��2}�"��EȻ�:�=o���}�O�Z�x�&=��[:	�I��|�Mz��x���ӳgO�����&�;����Kfn�5h���r�_�u�ό����Mtxt�{��G#f@W&�COFN����!A������K�(���9u�>��.}�������}���B5r�z�5-L��6.g���}�!��A�ߡ��}z��%��3�k��Im�D
�Z��^�4��ݚ4��̙
6��s�FE��7h㵵å��olxa�{o��}�:7it��@����z���BxNȂ�w�cp}ߠ�cK�^�����A�/���,zQ#��C�����O+f��63� _^a�ċՒVù&V(wZd}�r����Zg!w	�'�N������h�.��x_@iZ���cVC�>�=�Ͼ��'n���^Y�r����f�Ϸ�C�)��c��e���q��a߯��9��@���eh�����XS����`_��=��}����=wν+M��}���h�S���f����z���ĵ��8�k�GWxw�yM�#~7A �	F�����k|�+Bf�hNVⴲ%�GT$�o��
��$�Y��D?��ɓ'���K'����:�n���.�N ��{�wIA{R ��ans '/R�!"��ITz�U��s��Z�;l�w�zh�e�T��uV����./�YY��m����L�wZ�[�T(���;:����@,���� ߾}��z�-��Gg�����#z�������N��.��}��7�}7��a ᾵5��W �/_�����ޥ=�wݱ����=�f�X�a��+T���u����� ��4��t�e=�� �cKS�	������Ox8����3��:���h�d��O�r��z4��M��I�N�2�N}ן��}��}{��}k��!`�Xt�[`Xd�~te�z���ѧkC�6���B~��������k#�(�~��[��`g�͡�<��{ l� 2���"M�:c���]u�V�c��a�@�8X�rW�.!�m]j���6aEG�os	x�<��.�w�g��B��2h��XX;'���)[�:�,�eXr���8q�0�~G����)���cˎ(��z��خش��4�;@
�eex�0�U��!٩��t�U���j@Ac�>n���` x3p��T���1���j�Kϯ��㠕Qio���+:ӫd�kTZ��1�>R����ƣ�V�U�R}��\�<�8��)����;��ox����`MW �դ6 �)_���*<^�A^�2�C� ��{�.ݺu+�L�c��-[wm��>~|�uM���� X'� ;�Z��s�Y��ӳWq㴙��c(+�D$.v�_�΃9�p��74��_�|�@�1Gk~��!���҇��ѯ~�K���G���'3#8��^�Qb{g�<��}ғgOigo���]�Ϟ���!��Ş��y��[��E��Em|��wG�G4����BZ��Ĩ}�o�9U�e�}��Ak���?pB��;wL���HeX;��"�~��U� V��%�#/�ښ����X����N 8�d��	N�+���#�0�ɀ��w���}���	���9�։Kʇ3� �`4�^�]���oio�67��6� ���I���6XRв�,r�{֋��~��Ս7��T�J�Qc?���^	X�;�_�"���j�^X��� `Xiǜ����h�|Dk��5��0�1��װ�D6l�a[��>!���l��U��!w��8�}���**i	�u5�Qzm����W*��Ha��u���S�PxQ�U߿�o�o���]�',�L������+�J�>�3���#y4�c\w(��R���KU��wl�p��YBJd���Z�����Jۂ ?AX��_�B���o����l��.��bN~��#=_�@_^��� ��(�ݥD�ycx ֊ �	�s�����B��?�y/]�Vr�B����3e�TKgA� �
% ��ش7U{����L������z0쁰g�X��� �-�Z?��C'����e,���n�"��ԝ���������A�ό�����������u��Tx�~��u���1p~��1���>qN��Zp�@^�����+��YX�d
-�U,�P�JI`��S�����,����&��) /!�Rm�+pbM9��i�/��o��OJ7,�pvd��<d���;�{�Y�ou},&�j����y��r�+䪄d	���?(C��QMg�q�Թ<�⚇Eu���O�8 ���Q`��i��ţ�c�������/ʴk׶{!�������gLX�L�z}�y����e�t�"��|�����h�sТn�R۞�V9��_��<J�x�5:^�գ�>r�t��aN�Q^?��ƍ�.3�0�ъj�^��ҋV_��DQ)�yE���+�y�d>��Ӡ�����	�P�2�������<C9lm��Z榭����Ԏ��y�̉�k��z���Rm5
��W@��Vr�D�I�QAy56�"�$�7��Id&j^�縍�w�+���<��+
A������#v��%{���VhX���ԟ;	 )�ˮ<��FK+q\TZ�4?��m ��\zF�2�e-�������:�vK�,�h�v��W��r��[<����70g���ƫJm�Ӳ������Z���{yf�yO�H�nF�|�������Vd��V�GY4)(��\}%7]�����3 ���Oy��cJ���{z����/�&#�Ql��Պ�I�.����tG �~G'Arb���g `�O�1��&ɚi�@R�I4�[����&޻��+��MÞ#��pO�W$&�1;�������=r ���PM��'c��=�nb�$�h&�'�X�D���B��6bz��VآU�y��>��OI��S�}�c��VfWbo�lz7��-�
� ���T�ΓԂx���[�"E������4i^G�i��A˻% �*������[+��c=���%����kQ4�t�UP)vA*�)��~���jik|�u��	�7��w�*~��fUՌ��&"��~X��G�E:��1(���~y��Kh�]r�M[��)'��R�c��z����	���q����<䆽�Xa�6�$��V{h�SE.󝼲5xI�\%(�E�c���:�
��������P>![0ѷh���C(�����q�ܿu�����\	����>�y�k�{2��ǵ�τ𩌚}�䦮�� p�,Vޣ���˖�c�КxҊ�.�f>���e�L֟F;��h��2�\�Wq	��e-���cn�����M_��	���O�gz��Y�7UofN��|,�ϯ�gh%*����w��}��׌K�� ƥ>zr���1xG�_�^) �)X�ɻ2AP��HV>���｡��`��� �:<��c97-��&g���54��t~��[�|z�\X�x�|3H�{�>*3/�l�s�S�B��	�Y��"��rU~��"���B�����s���~�c_/��� ���7icO@U�k��u9�[b���(I@I�`+��`Wg���g���� 颢]̐�Q�H�W��d�j�͛.��� /X�L�g����ޓП>*)�U�h`B��r�������<�(�<C�
�N!(]��t�Н9*�)��b�9c�4�������9�����^y	�1��Xc$6�t:F��eU3(��#�Y,�K ����>�3_9~�͚�)�
9]`�`u��M�)]3+��5ք1����<��-7P�5�Ϟ�|��)�����&~^�QQ)�z�D���W(0c�I��!r<%� �E�DUC#�KP�(RE�D!z1�Y�+��Y���jU2�"��c}�Z��O��(U�����j��g�$��x�苳v��c/�����4�k���|��o�A ������Y�/��R"��]��_&j�rѼ)O$�ͣ��|~柘1�e�	 �Azn��z^An�AF>��� �g)K���4��+�����߻��{��޺�Iׯ�hs{b ҰϑYy��5�~�A�GSz�t�^����5�ĕd|��Z[�+6b�����r���c�����y߯����>��n\� ���A�t��/��� ��O����غ;�R�D�Zi0ȵ���ܰ�4����X��N���_7VP�J��<$ G�ƓD�ט �dK@�MTC-���:H��Y,�u�����l�-��E���t�)y���ٿ[��\��	y�ќMzeI7���M�P�� /�R����C%Ͽ�L,X��Z\��3�?A+�<C�M�CQ��e��ka�����E`�r�X^W�R~D���.�H[�䣃��6i�s�f�[�$>�Q�J�U%X/!�sV�h
�� VM�\j��ű 0�� Xe���R����`�ژuѱ?B@.ig#���-�L���ע<��I�)5]R��e7�7-�PC�gX!��uC�0)c�Dz�� R+]�y�y~_}^��*Y���G�=���N
��{���D���MI�����w)
/�B��J| T�v�qLTߗ{~�C��G/^�9�1 ȼ�H�����m����h�.�揸���v�e� �>���ڤ7o�ѵ͚�4,�6�_X�j���?�9�������1MUj��������ҋ���{z����$*4�a��-@�d<�oC��5��v���z��ݖ8��+��k�Òߋd�phC�`�Z��W�Y	2V|�����,�ܺ��2��M;N�bN��zr���<hX����R�g�����o+e��m�'	K�^����^m2z���cCх�|_������
��<� q�\Wްn������,�\o�����z���ٲ4��5W@�GU<X��+0�Y�JV�y���.�hq��iM|X��2����w	Hr���{З�~�v�k���b�����S��*��-H֝���%�O���q��X�_̮�$�!��#l�<� W�RԯiohCy���M�&��ƽ�6d��D�R.k˳�(}Az]�� p���ξ3�-`֯�2\*e��^%b+|>����d�K�揭|�V�.ʕg��6�_��<��7��O��e猾�4�Ĝ��~����5����wY�p�8�ݐ5�� �!KH�_�%�0�I���\\�TL��c���-��{D1�V�e��Z��������i�`c��7�ҝ�䭍hЯ���Q$�`�7�3��1���bh�hD���Em2�5i�B�߫�� ����0@z��`5�8~px�x�ߛ��5,��/��Y���:�X8H�͛7��kt����M�s�Ǟ�TO�u�`��EK����)��҂b�pv���j7k��<i75�)4͔��-?�ݕM!)�R��˹�^�dK��1
�����܈�.�"�۩��z	��C| �/���>��c^�@�������ݺ��`\�ӟx�R���8=�݊)�^��`z���
�iԮ�>�~��Ik�5P0���%��Wj�˔�unQ!`�k��@��l)A9Vܞ��NF:3�	je"��fs-�0��،�Q9F4��¶�|�/�e��Ē-��J�%*�Զߧ��+Z����R.\Vp�-���Q\����?�9� /�����_��=� 'D/2d�qH�Q��g|d������?����qRƞfJ�K�۵�|V.�le���s xП����z�l�o�#o������BAnMm �� ���;���G�>m����0`EGCӁ�oXe��> �x��׷����7��;o�����t��8���r����5��֛tp�CZ�X�m'���0� ����#��*�G�\��$8��4�ga6y!0d۴B��!�,f� �c��)�N��Ϙ=��Z�}��1q��+�4���]/
����?JV���a�������Ν;�����0�+ ,!� �7R������iL ����{�4�ZlA9`�`z8&��y��@����E�H'%�0ɏu��v��:=��O�6�.j�O��,m��5��x�Z�s��VΨ����B+aKe�5̷#E�(�1�����%��%��o�	�Z#��y����xq�I4e!?�w�9��ac���#@�Og���gmhX�{5��@��L���{iL�c���=z�%�z[��)���wP���F��"�k��i~�(����)�h*�Ӹ�|���E��i�U���kI��9�sm�+���_�'�ِ���k��+ڭ�l��� �"W�\�Q��ɴ
0�T XhF����������QX{����1�כґ��WtXzT#U@5�h��i�FD��|��G0lI�r��@��@�Ā���~ƹ<���� a��{�!�w�}��w���w�q��&ܽ�m3 �z�����c�#��ޣ�o�b�������C��/_�����a��=�p>B .��%�Ε�OE�^-��4?�iPA��^�8���g�Ϗ���ƬU����|Ap�k�_��=����a
��b��H<T�F�«5�:�֞Q�W��e��)�p���ŹI�x&�� � �LJ��H�����������+�:k�{���v�D:ߩ���^��-�O\P�;ja�U�	P蕿K�*Ņ޽>������C�X��v�/s��>���v��i��*x�H��Z����*�����\�4O�˽R��Q����o.�p�Cq���^����[
����}2���Y~���IƱN�İ�j��&Q��=�������׸I�=�zQʁ���2wOB%˜���� n�\qX�O!k�V�.3NJʠ��']ʮ|��B�_����_������y����8��
_�y~�d``�:x��-q?���+-�U�����D+/��N`dC���z�V̑CnA�,���|�g��9�KE>2.����4����(� �@h;��W�<km�p:B ~,߿�>�w�676�=����m�|F�A��꡾p��(�T��C��۷ߠoܠ��NA��[�U�We~�\���aO�I[�d�-�ό�5[z[��i.8��+ؙ���]�x�Q��\ �Ϛ)J������8�k�A˞���ߜW�N%we�E�ߡw� �g��S֮>�l�r�ˀ�=�Ķ��r�H[!5��n��B:7���o���0<00��i#��E���a�fb=�{����c��D�`�VЋ���룒ƨ-/b�EM���=�%Kx�N��etk�еJI�M���ʹ>fM�����pKEb]lٲaC�wx������9PH'^2ZxUY�2�Ȇ�Ed��ޖ-�������J5��Z��*��=����cF�6��z���eymS�t��E�}�{cY�8��t�d��k�3����_���D_����V ��(L�!__�g�e�ByM:��zyw�]Xp�����?�o�fO0(�E���㘗rpL������x��{����_~�� x�/C� �/'��w+����{��-u@�ߡF�G��k��g�g��?�?04n}�v
�=��R�����Çcp�C�KV���4��;o�ݻ�; |���/��5%p���Z<�xz����ڐn�z��}x߁�-Z�X�ͭ͸����ƓiR�`a�?8-�99�aP�U��3EU0�@�?���5�Kz�D�C!I�v��J e�L��nK�܆�o
e���z��*J�?Bߋ����_i�gϧ�����.�W5��P6���&�E��W'L:�ҩD��KS� �y����I���o���1��-X��,�b1���8'�G�@K0�%"ʅwͻ�K�7�JC�"��aO�y�@wQ�����,o��� ^�oQ ���
Qru����4�ϝ+hk�A!ŵQt�ރX!e�o�j ���t���n^�:��6�c����6�a��r)m4S��VZ �᯿ת����I������4U�$�K$�p<�j�}�6K�x��(�)m�Ep��(�*��6�S~��oR'�����:'�%:�ܻ�П+�.�z�H[���0V�璀b����˽�}�[��s�~̠��=���� ����������?2���Xo�Q�W� � �r��?��?qL��?�����/ɜ��T��o�K��d"S ,�"���7��:ȑf��m�=K)"A��o�v�Qk�=�4�¤H��HL���:���7���[�<�������nӳg?��^ �~S�`�ڧ�wp_tt�����w�������'
E�S���[>2tвG5��Z!}���gF��� ��
]#����2rI�Y�E:���?�_�jL;s�L!�Pn��&�H�[4@8E,LyEj����bp�������/��$]I=ki��G�tyZ$|C�Z�-�n�kX9w��=��:Y�P��x�h ��iJ~ADև+��]��A��EQ��)��v���wh��~����.:oD��v0���WL���f�b��J�c����rF�ؼ�P���_���͆d<�g���4��#ߪUk�-t�g�ҳq��+���G�c@]��� `���D�=����s�+9 ^K���<_��E�����V���z�>�1�g0x`�,hP޼q�����O��Թu~
�y�J�W���I���	9���E+�xE�*n�ڋJӢJ�Ӣ�2HAA:�m���ׯѝ��0��<� V�
�o��-Lh'�����0/��O���y�J����6m/�6}�"Pŋ��]�>����V4��I,� �đ"�8#�[���'�#!7���8ѻi&���&�	�R�?��Fh�6������l�fTO�V|�7Pz>�k]�9`Vs��l(,�#7O'�����D
&|x�%�R-J3�xkc+4u�Ji����'aZ�����^#:OY�[�Np�����Ewg:�k��(c���^<Y�'!gpN��s�,#�KY7�,(�L�b�~����z`�G)0��F�\�,W�����Bک���y���:�}���7���Q�B)
te�����Q��vҊL:��5��E,�g�8���o�:)�'�u~��"սm���n�׊��4O��-m4��a^�]��Gˇ~H�|�	[�����9p���=���	�J4X��'��=�/ �V(a��Aj@ b#O�U�g����m+��Ef�^d�f���Ǟ�����A�ݦ�y����ӵ7�Y�0�t �D���1�s �A���&c�&=��}w~�|hWl���A����5 �Ʊ�W`
�f �b('d��Tq� �B-�B:�m����^�;[����{o�r�{�92��a��OkdzCZ۸N7n�Ak�C�J,���	�ge�U�p[����åW���l����3U�m�x���UG���DI��쩾��v���ytq�Z��	{���]�����\|pL`Z:��( ��>R��[`䂪����x�O�S��i�ϒ�{��m��w�i���܉��5I��6����`��m1[C3�ϙ�bik�������Y�]j���7,I3���?b��t�`-'����<�(��Η�/2~�]��{���8�=~��o����G}��&5��u���&ުk˕��d$c��]�'(0�}˥X*��8��m-����9�<;�EHmwe��w��!����(�V�K��#h��Uρ_Kc�����]v�o����=Zs@�v�Z���'D�C�9�ka����4:v�y:r����;�����|N��	�P+	�*���K`�`o0ܣ��=u�Q��� ~�7駟L��۴1��z2>r��82WǪ��Y�j��~o����s=:���p�F.�8�j��
@��;��S^�]] �7�����������9����D�W(��fCT���+:)�=�r�@@U��X�^�@�����A��"���b�\���Y3/nS�% ��6���\���Q�v����Y�2�	��/�!����S\�#U�ա�*B�e>�g�S�J��7	�eO�@W��sgM��r�޶�Si����c��"����|��o��oy�$��-��Z'��
 _��S� W�/x�g�ƐmA4�ȭ�g�O����v�"V`W<��q��n�k�}$h�����tipN�΋��[[���yxhi{gB��@�p�/���p{��ݽ1��ܽ��am;|�8accCc//�2DL�uB6|�uǡ5��(�N����PX�oܸ��ݸ�s�:>�w �����w��&ZwB��{ߊ��'tp(�xՀ�}�Gn^��8X��۬������k��:Z��HH?�67lm�c���d�-�~�YuhE�fXC'�A�m���D�ԡ��d,���
�ٲ��w�^��x���>#��i��{�ԧ
n�&Z�/�Hyv�n�h�B�~T�.#��v? �/�
���^U@s�:	�o��T%wȠƘ���ш����8�{\�}꼋�|��Yh��Y����sIm���8���ךG+J�ޘ�w����fv����^�f���Ȏ��H���F��E�i`�6���6wD�}U���N,�H9�H�]cċM�E&OB��P�9�\��Q}}SӬV�Ӹƨ���m�<���tO~~ 0��b%�����>_|���r!@� �X�چt}):��t�OFEo)��x���4��3D/F�B9����+>yV�E�nױ.w�/K�_	��u��~p��,���e�q�� `P��Jǌ����iL�D������F�0��Ood��St�������?ۧ�/0t�:�h�	SiP4�LlK�t$@��/9�3\^��8������k�w'��$��O���#��k4 &N��������ģфF���k8o�Ǯ�:Т�'���-��{�Z��a�<X�b*"�k���� X�����}ܐ�=��U���"c��ZK�.փ�x�3zJ$u��Mm�� ���diS �A����7t�����cQ�tK|��~���k�c%���@;]����z��\ϻ~�9_��퉋����ȯ4>oj��3q�������g�kuX���ȹu��TkX���D�q>��.�Kݮg	���=o��<_��]�X��)8(G	���?B��#�n_����K5�,pgw��^<��R+ �-�A�$٫�ߡ�<�l\��r��*���+x(�������o��r(����X�d
�Ѡ��X�U|�/�6ėF+cRW&���v�.k�''��".�zL�%���9�?7�"Y���a� (���/�� �zԽ1���%��W�=�u!����xz_/���7ady�������<I�+�_��3-�&��ȶ�;dN���0~~ȍ�p��W_}ņ���4�^I��~/��Y����I�A� �ց� 0C�+i�?���5��1����6���]�7��;�Į��
��Z��1�r,jx����C�e8�9-��z� �u�HJY��˴w��>��d߁ZL$��SX�}.`o�uy/����x���1�j��%h�:�?��vy
B��h� Є6� j9��\�Vl��FY>�[^x�V^XW�v��1��8g/M� k
���⤮�V.�����My!k4_���k@8޶���għZ�'��&$�V���ܧ����I G�,��Lhw��r�^U�*�����5E-ߒ^��u�JjN�ѐd
�V %$`��@@�W&�_�8�A�"��(��&�?ud#�cxt�6��O�VIS�z�1.
y��
��t- ��L�;䢂RɅ//���5ϊ�f�c�����	��c���^������M"�!�v����������	���2���1.fxv���s3*Q�c�K�2-��=P���7�ヽip�+{�H�٠����-(�k�����l}�Y��%8�v�g�d��B5x���*3c�F���uƿ^&\��$�:r��+�� k.����[���kk��
��>~��J�@)CK����/m�W�/]0�cW[�u��E��-���DP(|� 3*;���u�ǇJ 8?�]��tP0�z#��;��J�3�z��v�<�wC K(HK�[��Ze=y5 0H@D�D[n���u��QM�cz�:��kDEh��bwg������w5���L4�w"P�ojq]��=C+��Њ��ѱX���籇 a
��`��7y�����ݷ�ѧ>�V�
P�.���G��^絵-7(������ֿ�OY ��-½M��~��N�̫�k�c��1G�� 8��L+.�C��N�#b���c�
��,°�s���^꽖�e@G�V<� d�6���/�ϟ-K�-b���4�22^�W:������i�c��=o�5��kb� b� Vyc�X�}y� �ؚ�m�\�{�}��<�r����i*�_}�_�LX+K�>?m %�Ư�J�$%~�N'!�o�] ��o��F���N/��˭ݓ`i���*��i~��~f@fo8�\��z�=�ZH���E��"@`�
��l�i^��J"��?X���֒���r<�7�;��c!z�VNǴ���4��ZP��96��9 ����
�%�2�-����8���h�8������o���"�m����~-����#������Co��AQ��߻����31�F�;��2�l%eI��Y򊀶v;=��ܭ�����B?[?S��8~���}��=C&��bs�b�:aV���fNJ��@�]P�0`����ȅ0��P�w�Xi�]�����J��bH�9���k��'?�	[r?��S�p�W?�� �A� ���?�ßp��8�f%/��>�ӫ�A��O��"�d\�Ѥ�����=rs 	q����r]��u�c0f��W�l�\�,�`�` `���>�</�e2���z���y�6���)��w>��V�J���
�d�S�{p����,;r�8Y�R�����k]���hJ�?ڡ���tm�r8ȵ�����$ �\�|��x{W30n�m9�[У�;��Ea�{�EH���Yi�s!(��}"����(!���6W}�0����{f/U�%�WF=�6�km�4�;[ \�w������ۧn�[�����J����!�&�	�����M�І-�?z��ۈʡE^j��r�C�xd���y ����xQX���	^4,�[al2�8���Q�%H�MuE�M �DA%�N�I�����(���:�k��iX�K�E�\�:,#p� �	��hh����A�OO*ƈ�F�!+h��ٯA�5�x����à�3��p�az`��=ן�|�R��Լ�w�k��H���5<j�:b+�ᑥ�#⠜�r����b[��u����4�=:��h������Z�RRR�.�����g7熍�1�z#�b�E���x/���XҮ���}m^�_t~����m�k려t��+�C���`I�ŪU���.u)$r�(2�%r=r<�#�!�����9z9�?�R/Mm�[Xj����{��c�c�ϛ_8�.�U�?yL���o���R/_��)d��d���^) ,���%&ԣ�7-,�3M���'0�k,��Hr�����ڡ�O�:�����a��w	������o�z���7�_w��h}�3\t���7~�����TSn���r����c���OB��>�\_�n [z�|�~��?����>�,�0�^�`D`iȞUP&x��`��!�N��m7Av�	XA�ɝ�.t��$!j��;��@4��6�� SKQxт�Y��D���}z����b��mmT4z|��G�zGKb�U����p�&���=}�O/������9�^�[ �F�V�5���j�P��W�Lqo9�3,���������%W�*�KRVU~-�*�ofN5� ��7���<(N+�/IgBs�6�P��4DP�#Þ�%!��x�]o�Y�E������t=8����ȭ+}��T��{��� ػ�� �'�٣�۩;3��ۇP�9.�x�����4��6�����ш��&��� ��[��������PTJU�bK��z�	�N9�'g ��Wx����:��2�}z��|��ϕ$5��Fa�:xy(Ս:�'����_*�C,k���6?��uY�}��߸G����FD�|���e���KZ�I,�j}��[���*,�`��R��Ӣ�C�횮�1��|����K~?| �u@�6��%�;�`~���[���f%������+����X��]���7���d�.Pr�bQ<G�&��Y��V�Ǐ�� 27o�����T�*.�� �o b,���{�r- 4��������k7����;�G��w�v�#����W���9��5 �>����r8;�vȖ��(�M���i���� h�O���F^8+����m��h�v�$���A z�b�}ӎ[8�������((&T�F{L( L^9��o����񈅹��:�.��ה�k��=֩p�?�:�gz�G�����;��uE����/�W����5�����9�
�IV��a�#��!��i���\���UK��K�rr�!Y��@���b�`s'ݚ��g�W����TRո���/���JǢ��a8P���)�4,������1 �J\g��]WW`w��Xě�@m ����#��������Mwk�tf�%���W�
lzk _�GO����:BnM�clcv�D6W�����;$��U��U&o�!������Rͷ�.���h�s�N�mT�3����<:�:�b+/,� �� �Y>�\�ï�˽_@2��2>> �=�a��\�W-��ů\>�I0�` X���܇�pP|���lQF�b�=��ye �'����NVb��b�<_Kȷ	G^v���p��}(��Ggc�`Q�����,�<�8�A�,�v�$�:i:HG���Y�$�q.�Y[wϾ�� ���P&��5Ӌ^$����,3�Az�i�%�� 0f�^k͸�y�GzFEfU�����Tu��៯��(���Ф`��,0=ު9��9�����1��]�r :X�E�.�ϒ�#����OVC�=���n�n�d�@�|�B/a��BX��@�k��A0��hL����X+Z��y�֛�/C�PQ��1�7�Y��M(��O���ʋ�Zp줎�x��7
}�Y�9�J�q�>�Lř���'��+����s�0K�3s��a����81>я�(9K�����[n��X���9�k�/b��r]E�p#�_ϩ���`I�/�[������6���W�@��{(T���鋯�:aЃ!(t++k	x����kx�GG3z���ִ)+V���ǚ*uy{#�>{����+V�0��]`�{��k�={���z� ,-oJ9 �=*zV�z�C�o�=��QxY��7���5���ƕ
/gx%���4UxƲ�#J��2�љ`�ha��Z�o�� ����6 C��29��A]�/R�^�b��}:��y��`-w��9��j��. - Zp
,Ȓ�������b �6���Lx� � ���1�I�+�`y�#>X,�؏�q>H��5Z��@^�n�$�Oу;Bm�昪
�Â x1]�ص	�� /$�L��Mu
������|���8�$NZÛ��"�'J��'��Gg<b��(�@��t6a���O2eI���.�gx�0ˊ�PQ�B��EF��N׹(ϏΦo��ʆ$�,���0��.���(أ��w~NsB>��P�P���e�`�8��p�%�B7�띆�K��OE>*\��Y[D�H�`��va>�]��tK*;���ɷ�_�˗7){����JQd�&�0��J �=��{�XS��#��4�&�p��'�N��]���:��K;��=�2����.�8�?�q�3?c_T^)����
��P�"�d�2�_���5�"�.��X�����X͟V�1�ޛ�m�u�:�T�b!�<=��Ȇq �q��R�sm��nR
r��	���rL���Y��8ǭ�+�-�r� X�-X��!��Y&q�����: ��M�u_��W _]�E�/ ���c�`@���?&��᪌��5�2@��v�ݬ��E����t�n�s�F[��R ޵QFR����_�KS/��	��5?�{����E�>q&C��[a:������+��^&�Q�-6$Z��մ!��`]XDa� u��-�A�;_���90�_r-[��IK���F�>y�0�����͝�?	pՃ\�0ۑ+I�0S�ؒc"�G����s�<oa/���+̀��J�"��9��)�A�V-qEju��.�m�u�MV�O��\�����5]n�Y�:4S��x/�;�О�O��x[N@�W��s'�������V_	����A�X�K�<��&u��<����͇<�,����l�8�'�����vI����) ���+�P|�GSʁ�O֬��&<go�y���]�]b�%�2+TȀ�*Ʊ�M]�=���Da%!j�&m=��ꚮ����6��8����J�^�{
�W��<-��z@������9G�7��2����Z_~�%�C�Qp�g[E� x��Ojd!���ӧ<0�ď}��l��K�E09Hk�e�hf�j#5 �`S��"�xa������l���X �HTrs�A�>���'��B�N�m���"Xk|�>��@"�7x�'�)d���4 �P�Qނ�k�ok:��AЏ"�U�ks����>�7�$��_3N(��(�f����^A>��h��pY_"&��� ��+������ >�A��am�L	?�����b/1p����m��XBWjQ�ev|͜7x{�ŌF#K�#�Q@��2dq����Q��P^���sv�"��Dm+C\�S� K��գ�Z jX�l3I��`錺r��6w��}�9N�n����H�C�E�$�ʲP�^%c��E����x�Ⴖ��Y6Χu������ �D�-K�?/���L�[��M���Y�!� �q]a��2�=��I�|�A�a!}k}�e����AFY�})�f��� ��i5 ޟ��V7G�+sT��R&w�A��=�����a���ʠĵ�ˠ9'r��׵�M�>F�ժ!����E�I�W�������'}o�?NCm� ��cG[P�3	V��9��ζ�Ѳ�1�{��������\�Upp��O§�.�6�(��P aQ���d����u@�5 ^EJ�2g����ʌ�p���tJ
��0fB(��.,�|�0!�o���_�EL�!���vΉF��N���V� ǳ9gx�}�AA7nm��;�hks���9��X,`��'��Q+2Is\1>�Y���tA�w�igw����;6�g�⮻׋��ծN���w!ê�kPX� ��_���w�����^?�Mc�69��-&4�hk%�t����KW!�j,�*v0�@`!�]��_d���b�`�1|f{���ͬ͞��Tt�XF'��X�ڻ�oLf�����R\�+�Xx�"���Xy�v2��oYB ��`ا���t�	� �-�쫬�NtGR��`���X�3�M5w�l:s�񐎎i:AB��R'�q�l��[!9R!��z��#^$�F�ӂQj5�}�#H����P:N��o��H
����,���S�h���ٵ%2�O�M�G"�<#cf_#F��{��Q�F��p�\���c���Oj�Y��V\s��ڠ����c��K��X�<��ay=-�K������|����C�~����ߘWX�u�|/UԵjE}��޿���A��R�6!�?��bi&�6����x�a[U=�e�B� ���H�2�R�}����u��jiR#8��f��@iQ��y�=Lr���s���X�@H�ji��Th4�vmn�e5m�U�L�W�1�hH��"�M)�. N�~9C�np{�����+��/~A}��AK}d��� ��u5���Ju����H�$��N?^�$ya����$�joo�ӥI&OZl=ǰk�2�b@`ʹ�EN[��-���Kp��޼A}�.=xp�F��"N!��+ϩ� \߷bC#���8���E1p x��������}��M8i?�0�f��h���|n��*��q������m�ogE;Dxi�N��#&lHw�ܢw߹E�w�n�@����^Q���Lr�|T�~d\-�>�F7�����=}���������K�Cu����p���X��8�_��-�
�� � ~���hh��Û�g<r��=����w�Э��`��eR�"c�2W xAXf?x#�RxBSPĻ@-ꝝ=�}Լ~��G����9{;�2Vp7�rj����ۑ3�箙�,�,�]V������J�a��3ׂ��Q4D���|���֋&�'61HCm6 ^[[Re��%���Ed����m�2�/�nr 8��X�b	����F\+��d7�+�K�M3�����b�:��Z,l���{r���Ғ����ZG�i�aV�o�=>t�T�G�T��kb�	#�@k�%���&1�<����:ߴ�'�4u&��P@���^vϥv��y6�^a�y���i���5r�I\ŵ,���Ɨ��x�)��:|�
a�k�W?O:648�g��%�����a�Cd�x`�FТ�/��s�9��q�d��� KH�V����t\�z�k |I(���I�ķ�R7!Bo珃U���Vܣ��V����*'�,tΧ�qP�w �&������.��r���_5���B��'�1k]K�~��]�	��-z��'�A9���1Mf�X�	����� ��NM
��Ex[u��y]w�N%�I��4�ԩHī l�4� X��9 r�~����g?}�����DH$�/�!Sj8'$n	�y2�W�qe���4���>����g�����٫��QZ��Mc�Nn#��w`^f�$	���d�z��(T�m������?�=zا�hC�w�m���|e�L_&ͻ�s`�؟��~"��'�)���f��y��^	�ɜ������}N_>yN�|ח�� �P��r}����.XD�=s	�ͳ&-8
?�X��m��ߛ�7YkP���K.\�9�b kQ_(�PsX*b�-mA�uƬ|ۭAomI��)�~�UV%�����Ϡ����Ͳ��
 7�\A[D1ַ�(��2om�$��l��F��[��mj%�jY�6̑*�n��c29rs��!1>����alf��D[[�9(*�B�5�
J0o�&���{���#�T٭�g�`\%�2L�+��(���E���/�>���;���oR de�phQ�\��=�VqO�\2�ęΧl�Æ�郵[�vPh��.�t�~*�]��B%9,��P�J�(q3��<�mY�S�y��Md_��r�y���MQA�B1*�چ9����{»C��_��_�/�Kv�FX����߱�����\	���������q��$Xܣ���Jgy���v��]5�  N_����$���t���ex���V�����b�]>Wb�{}��a��y�k�o��b�Q�8��cvݿ�I�=�M�n4�;��˴��Ր��_Z����x�Ly��}��mn8fV���Ը��������S�?
m�>JK���)��$�Vw��-˃,$lm������޻�蝇�4�s�q��P���+[Mz,42 ��ht�f�nn���4��S�&Z~Z�6t%��npM�B��`N	�<�g�%Nx��A1�7
�����7K���ss�G��P��Cp�\O*,�W�U�Jp����-�U=�q��	�n9�m�捑�|Eov�qp��0�*̂|�2ڏkw�W�Rj��vYLr�o�X���*8Y�5���s� �L�����v=_- ?|�+~)�ԢD�����G�y �!~�p-���|rpُ�.�ajU�����y��k��Ͼ��^l�0	8h��J��0!���7�����h�7A�Y_�" _�U�o���>�?����N�zM�A���"|�ƇlMC��Fz��/$m4�$��m}�3�z���JF��m���sk%��*&R�`�[�	 ��+��:�Y,wF�	�� .� ���O�_���2�: 2g��:�,Hǧ�C]�A�72�p������������v�w�7���˿��@¸����	�>���{�����뉢C���E,�8n�o�t�QH�Қ���MM�R�]C��9��t� �KD�6A�M;4�����>��O�_A��a�K�}���� /��h�����7�N8�����X�����P�4����A�N���-�y \�	��ݠT�WM����C�Fˮؘh��G^���"��m� aO&��8����Յ��A�Q]ڏ�CȌ���O'X���ń����H�>��֖���j� xz0��d�-�!��$m��m(Q�����_=�X<�	2��������xY.��3f��VB�]��N'pO�;!g���d<����]��޽����"�B1���W�lmܦw��ߏ�ޯ>����^��a���µ�W �	ev*��ѝ^���$TE�� � W�����h����}(�W��
� �D�)=�{��L�/�ߌp����Ju�)X��Eˑ��[�=3���c\)5��s�S�RvI� ��z���AQ�9���Ic���OT&e���DW����C��J����k�$@F@H,{ � (;;;���o�_]�S,����t�c��"�4i+%� @$.� X� ��Ac}Y�<��e%�t������w��������O?���ƖX�e��e�>���L�LW���R�oCEh=��6�۷�$�-X������! ���wc�n0j-�,��l�*<��)8��⯎�G�K7�$5
�X�\���9 E�C��zl��mSgG�Q��>6�	��8��6:��@��G�ULj����~�V.j������z<o�yMM��R�$ X~��:�s���e|ĿI�U��V��9�x��0s�s��w`�Ti�k q��8�n.|b��
~��C�g�� S�s��"_3�0���m� �bK���V9XJGՔ������,��;d0�90E|��ϧ^�Ʈ����/�.�9ڢ;wnР }������Y�5<וi�[��gO:�P��i�n�uS�Ϲ���6��i���k��Й"���|˳�P�*��3|,[�H��Rk�P�+�;��{>�ൊݟ��vP�O@t�Df�T{-�LX�: 8�'K�^C,�;q�ٚ�7���S Xmb9�M�!����tB���Bw��łQ^	���r��=9�����
j���$c����w<�lcKbgźM�5+�A��Qvl_���Z_3�m�%M��̏Ģ*m���C{��za�� k��zŢ+.� ����`�qV�y���$ý ��6��`���S�{Y(ǋ�/�;�y��zޤ��������xoR����?��ݞ����3b|?��3��}��ATp����˼���P�΅�mj<�}rpJ�V�q��dt�
u�*�b᪊��]����>������O~�&�m�M��y�ecY(��q����9d��h6���<�_����TH�u�<��*h�q�.�l�9�r�TN�, �H�z�,�l��e�����d+����J�%��Ě������R~��O�â���<D�R���,[�{n��[x�� n��� <R���� ����f!��k���6�ӱ�\m�(���5[��5n����N(�; ZR�L�p(FG�"�ߦ�9�~u����S�ލ��рn߾��������0C%��l�w�S��*:b���}���p�������^�6�������"R?U�bJfL�6^���I�����g?�>��667���Q1��X����m��:	Vm���Rh�'k� `|���0핰��ۣ��`�]����K�#��P���K�����{,��j���5S��60���=z��9��?��+N�'c�/�|�]3�J����W1����'-���2B��p���{���P����a����A-�G L��,m:ɼ� sO��-�`���[\X���
��oxy��J5�{��OqM֮�97�6(��A������-�1P�ݻw�>|ȵe��6�?:�5�/�f|�F�L[�;iŲ_�) ���<rH"i)W������c9W�y��rm}����_q ,���������b��[�kh�AkS׀n"A�ˏ �~*�6Sz��}������??�;�o����cc*J�K~p�
�	 ��Y!���XL�-�`��w�p�єb��uZ��c�`A)M�^��( X=?f
+�>�I����o�z�i���j�d����̷�����zQ��
�l�Ӧ��l�Ɣ�?1�O�����x�l��o�J��y��?|��g�^yL�B(�w!%����q��d��k����Lw�����௼v��RxO�5/�Gsg��m�<, ����*X�\�p� �[�&3Ko�L��o��.\�*v�o@��G�f�p~���ݠa���%{�XV�qK8�ќ˻�4��w���������Lð�ʠ�UCg�zr
�Uʻ��۳���Y��-��b��xp�J�}����r]��l�  W�6)��X�,!&��N~U�'i��S[ؼ���2�Q�b��Y$���!��ݪ]��_�všyNYu������M�d�]	>zH�ѐ�~�5�|���7�,be�tKb�ɵ!v��C7I�k��_g*�˂^���㴊WԀ�&�z��qŊ��K�����ۼ(t9�u��EP�]_�ETE��rc�:x
"y�� �ڥYܒ�) XS[_vy� ��b��	~��4�)��h�ݻw�;-x��'��2۞[:y�� ���eM�"���9�7��X{�����Sxo?8�����_ΓB��~�+���b&���P�AŨƨ�d��Z����_^x��'c^m�U:�;�H����,h����w�u�Ϊ:>r���;a��5{!�b�[�b�0 6V���6Ǔ#��D]^�1*��ӅE�����'ӲXDB�^N�U��*��Y��(�B��j���m^y�\�Kt��� ��6H���S�e�D�1-{ûf��D�M.��-��P�����{�"���G�����Ms,����>�x-hQmɯ�A�4��Q�R��T,3^C?_8f���f���v7�i��s�
�v��x��������m�v+��N��h�̊H,�7?�1�h~���#�	�p�0�UT�X���dL���>=}�KO������� �>_�����>m�i��}��������^Y7��(X9�x�.+�s{�����ή�޸��.4�ՂպB�y
��RQ�(�Gؑ�ڎ��C8�������=������ڳ��Wl+ ��.WI�-��w����q�����Z>h^�4j�柹�V���~���-n;Oa� 旎���x��Bd�F.(�����}��oҍ��	z��44>;�����@3�rh!�)��˘J?D�T�����<P]Z%"�������`�R�8��/6���y�oT�K9%���� H>{�����kNJ��9���*\W1�u�b��W�����Fm��9b	�{��	n���@`m|�w8�0�����)p�~x�����9%���Z�3����q@��u�#�3b�a��� �OX�E���X,�P|��(?ڔ�Y�R�� 8�����5O[>i?-���E��(7��Y6$�
i����
�!`|���n��!�ڭ!� XY_GVbku��9S�	4��"θD�#X�X(	� �+hhM��>�4�cq(���O�OuO�œ]�ǫ�Ҋ��֝�Z�f��W����b�͞�>Њ���(���,�t�q��|��F	��7����G|Lb��>�KNEwU\��V-H�_?�t���P���;+��B�I��/���gO�n�z<ί�;��IC� ���ZޕO����K���"x���Ƈ3���g{�����9>V��#�G,��{t����������ܿ����,S�#\��7�t�F������<^�H!��i)g^E��v�u�ۦp��Zn �@������mh� Zm�0��e>E�E:՛^�M�|�ڹ�_N	b΢��DS�ṫ���,� lq�E�[�dB\v9���~m��/��._��}�{p�<P��]�wb�U�����k�`����?��_j�캬W��>c� X��
�9����uE	��I� ^�]�`�c�.nш�����RZ����$��X��O�7��@���$��6k�_j��HJ�.R��
>���dg��z���e9������������&�u(H%�J
���>����Ĵ|M�26){t� pp�4���eAkdt�� �T��:/k�OC��+H��+İ?`���q[\ϯ�8�����}w.j����Ν������g9���8��I�T��1u���
p#�5�Z	8�e"�
a>�jA<M�B��	�I�Ô��b�KJ�������0�l�C�p�e<H�W]�8>k��l����F�Yq������EQ�[(;bDȅ�����������C�o�L�:�'��Dl������=��M���1�0NnXU�U��f7���΀�6or��t@��#>e:��]%�1�q n�VY��f#��Xh ���zl?��DQ��Z�����D�<�i,	�=N�|�mɒ�ckBV�BbMg,(��Ht���V�H6(�J���j�S�Kj���ME�����T]�=���m$�Y��8u��U��',?&n�����:I}Uo�DD�� ����_�kEb:���石��} I�0y�8d�"cTS�Vf�r���é�{�u �x~�ӟ�E<��:� �
:oe�0��B���݉5_bmu�Ĳ�z
�� �%�ЧO��-��1����MLn��K=�������_��_�2.�w�}�����/��r)X�{R������!�`�JZ�c�.9nk���E2� gȴ|�܂�h�,�
�ʂ�ax��;j1�ˁwo���<���(�99���D\��6�ˮ��E��mt��˺�é��#,2'�S�%�38b��;�7���&"-*����<x�
��	i���WiB��E[���P#�/!�-�=(����c6s��ڱ�ټ��	���S�WN1}�������kt�����#�ۆ�fh,e��2<[��R����`&
;3$� ?--�;׾kt�*��k� ���&�W���s*2ɵl{�*A��%q�d��n��5�l�k �qu�`J�J-��9ks�7Y��=�#ײ&�ݨq��Q�*�M����ù�6ݸ�U�X$s?7��7�(����'O�����$��c{C|�(�NC��`�C�W` £A�ςgPB<����񱋦.tޔ���%<��ko�{S���Y8�����O���g�(��}��|��3�� t16�� �q]�����1^�6��~Ex�q�����v�CFI)���jƩU�6��[XNK�M�R�[����u�f�o%�J_[nH�р�+o� >c�v�@{Ƅ,����y%A�DB ���`F,p�*y�x�ZXЖ�N�n����������Es9n벒~��S>6*g�M۰�գ A��=_�qv��n(2�1��1�ץl�Ow)0���W�L3���E�"��g������~�F2�����;q�@��z:�eᖠ
)���� Q�e�8w�,j��ВO�k�"!� �\\3C	�����^�7/�����6/�iZe�ls���i=G�\��ծ��`|Z ����ymm��h|��{(�«�&?�%;���k�C�� h��"�#
�ӑ����C������ԇ�m�}8���Ut���ٸf��2�m ������ ��ӧ\���+�u776}X�b�|���ۣ�`E4�h�����a��3��W��,�?��O����g��dK�|	o��}�����seP�|<m�ʱ9J]���K�?��?�%V^X}�eY�{y��@=��x�0)�<����x���2Kևf��������/��%w�-c��Ԣ��s����0�@K ��!(͉��(����� ��f�mm: ���! 02�Vֳ���s<�hx�66�P�w˵b�a��_=�0:�X+�ʁ���>Q���ª~��B�Ő��b��\t-u�Ϩ�s׫�%'��<�o9�[�Zˮ��Yа����6wZ{�'���A�d�qz�T�,��:����R'�B�4,t���a�ʞ�.���l���p�n��a���G}2����|">#eSD9C2��G\Nو��ŕ��(ghK�rZ��J:�e�i�i�yV���1���>�|9��$�A�ey�.���'�>�����f��Ӓ+�4�i[��T7��k��Kr��0�r��.���8���1����eBi� ���E�m�'� l������4��#�T��K��8�1�f�=��
�������p�ƻ�K��K�EZ.K�)���Pl���Y�)W 3),bŲ!��5tI�|�8�{}�ڥ���/?�q�I/��(�.{��OHL��d���g߲�
�9$�`MU`<�ux�f�>��sz����p��?#�3kgl]����[�����;�4�(B'����1�`-B��B�v�K�^Akt��K�p�X�"闋bD�rE����&�4�5��eZK������(���h�mbٓ�^�/������v�[D����c�&�M�mX��܇K�Cx�+�*[p���E��!����VIwn�o��ˑ;�y��xX�+�ܲ>���0.��ft8��0a��Rl�w.��s�)���2�q���m����
����[�����%�[��kH��.E�C�t�,2�s�w��rɞ��J�T,�EHX'���1>������G��2$I*#��mƳ�����{&ԡ��gdy����/� �����.�\P2�
!.�� ���C�cY����aՆA	���`<����F���mҙ{�d(}Fvq/{��U���R�A��~Ÿ��3��O@�s��)I�$St[O�.% ^~� TY�-u"��Em�0ۦ`ߔ���rC���� ֔�g*�Ѡ��YM5�)IJwLNhA��N�1d��އG���J�%kz/L�"Q�>gW]pAx�<xl�I��s�y�����QQ���w�d�i�	��:h��(I���m̙e�o���y�O86��ii�w]���S7�mj�廵2!m�ɚ���ڈn�@��N�kq�h;jcj+��MxwV�������\hƊ^uj�������=G���ٽ��O�Fb�	6_�������ά	!�"�z���Ɛ>�I����9��8o�c�43�@�w{D�o��;#���
5�ty�$�����͘>�O���%��,�EzE��\���%�ő��ڑ���vm}�tzL�9W��r�v�j��Y:�ֵ�ȻH߉�������o`  ��IDATD/���,���⢟k	��K����oq�)B��by<e�i(�,s2�؏��� C�c��@A�ܗ�4���/Z#�{�۳X~S	OC�^� ��;E��>
'�K�Ѡ�5��O�5I�j��t�_�9ɖZ�&��!H�Ǩ�Zs~�9�Y>S���)I|�1( �g�_v�址m�۔�v��2|/ ΁ߦ�M�9���YDg'x����ў��#�>5Z�W��.H��h9	C���I��C���X8��`�Ec6�6���G��c$}A]Lb�+� ��ݾ�>����:�8kj�gB�Q��_Ȉ������y��=t��i��{a9u�_!^��~�BL!�0�8�����YW�*���Uي�y��r�5�D��m�����@8��3B�B������~���0�� /6�J��A��������2T[�k˯�%ձ������D�ҩ�����,�*�g���~��q@�r�P�OXYg`�){4���[����?�φn��wo�~�Ǐ6���';��hv-��n����o��wn��}l�_����1z���m�wm�=p{���6���.�'�J��`I.�k:>���QL_��߰��묝)�kf+^�ޛ
s���%����c���Iu��g�7�R^h�=+�%�4��*ebt{�����c��^��V�>�6c��������3gci��R '�~��"/�)FV�+=N���S�Sjx�Y[+NH9%�����)2#��׿f�9��8F,k�1o�eT�~m�K�r�j^���^R�X2Y㹥��d?��	��4���#���I/ޓ�"��uP�5#7�5[x��)Y�U�=��;��h��oU�cip�`ٲ�N.���P�i�8ֺ��j����(h�dR¤�I)Z)�F� ~��(?{��,+��ݣ��_R�����=z�>���cm@�E���?W�` T-���p��u6���iwo��UYu=`���������<(��0�_k`'�!�h��B�&�X�t��r%n�9k�j�C�(�b��}fN�\=�@srIS�B��E%wP��dk�fx�jHz�����`�uͫJKj�KH&���g-i������L����,��+J�8YT�-|	� 8c.���hT�� FCǇ
����`�5ʇ�>ݺ���;����m�`��Xz�F�8AV��X �����w�ͦ=��;p<��'�m��Ka|��?��4��)'���c�V�%�[��q�����VФ��U�Q���z��;�kNpO�\74֙�k��3��\�T��h�u?�
ZM:lH�NDK�j���E"��-���ci��#E�Ӿ��9��~Q�J[�����V_��"�C� tq[���
p\�1⸤8)��3�yAp�7p��DY��\�>*�]��:t"��Z��ȍ���s[ێ���$��K���[J �E���;[��ڼ5�\�Pt�l]�2
�����p�,�ep��~+���z����f}ԓ��I��	鿱�; /&)�ǡ04
س�j�}��M���8@��{��'?��� Ȭ:�8�b��n�x|Ě.���Ǝ	loӋ�;��g�}��O*�
z���f�˖Tq�K���2��B�k�s9k�U�V�s@��u��I��i`��,&�D54mLD='�^�S0rZPu�ޑQ!�s(���O�����y~%�� a�{�"(�a�5}�R�7��}���&P*��r����7̎��*�j�X���!ݽ3s�j�\v8����dρ_h�g~��r&g�B�W���lЍ��4[�ioB�^�g�?s�������JǇ�	����VYhץ@�)<sVf�).��V�a���Lj`�Ҙ�%��r�2t�%-�z_�eA�}��)0�T+ݵV���W������
B6Z<�V	����#����|�Qc�x�XpqO�y�'�����LH]�B���ӵ�q>d���Έt,;�#�XaxB,��~��,k��
���>�2mǠ���%)����j���3�û�s���s~�����zg�� �f���-|��.=��/�+y�j+C<�� ��X\�������:��֌��0�4�S\4$�8�-�1I1�0�����4&&�*�����	u���=\8`�����焻�yi������9�g?Ҿc~��6��8&���}�ZZ;���k��s��3`a�����dhE�n��nA0�z�|8���7�>a�ﶙC�M�c[��;3N^���A�9$��F_ J~[E��M��w�2�j#Q��fW�
{yo!�ҿ�"⟦U��F��g��e�k#�&�A息�D�8�Sl:�2u��GE)֞�+f F����ŵ-ݺ	@��0�8�<�p�0ő;�->�5�
��4Cw����ٝ��xN�~���|��]g�-�XѶ��I'���{>/:+˨P�����ڍWi����N~���f��I�焰U ":N�sΓ.�����%M��d����5�6��7f}�������
��s΂���C�D	X;Q�퀵n�RZ
�&>�$��H�/K��uH��yr.H�C���.ޗxn�_$�}�t� 8g|J����w�i��*Z����3�oi���$m ,�|��~�ҍ-7�o���V������mC6�\"	To��aE/_�ӛ�3����%�	X��,��>�����~�����$n
�t2�I����|`�{���|M���a�q�����b��"� ��=���?������񌦓ͦ��/8q1�AW�����4�r;_X�����u=$������$�Z�+N���S��6��/3#�'�U��m&'C�u:���_�X'�u��Xz�Ow�E�BI�x[�7 c%^�-�xoo���kW�=�4�]}��S�ƨ���]u������mA)	%��9^\�>>!P� ��XfÍ�+�x�ⷊ�%�m�mC,� /� +}v}><�@�K�~����W�C_~�������M��S�9�܄��ב���.`�&��+"D�M:n��^���Z�q2�Sg�a�wC���� �e>��{�� �/�ð
(��c@ �$ɵ/øYEx~���J������#�5�A9 �W��$]�\�����>9] �X��Yo�- 9aikT����t��ݺ�#x4 �
B|? .G\c0(��vH/_Ru ?�9�ӠPò�&��|z��Ĥ ��pE�	f�	�4�ֳo�9�A�yw����hwo�K$���h�C�ˢ𭞹}��{���K���_|�1x�@{��
�E��

\�yY���u]'}���%���4,�ņۆl��e�X`�!�K�sQT��o�/�Q4,�6�Ge���{�W��r��խn֙���b�?n�#Y��K��X�X���:�@�h|��oN4ǖ�fr��}���8�n���.�|u��ސ��������� �!�JK[������3�^�E
X~1gʞakpQX�6�������,i>CfIx�ҫ��۾�������|儺W�ܢ��|'����4]��(����#@�P�����Kr�UWma�.�9���C�V3}���$�Y$��ێ��-�����Q���\�b�$�Ok^6����(�|F��{͍CZ�?��.�Uo�7^ȗϞ=��Pv�_ ]i�</�
K��B�$I��^vwh��!	�p+	��� ��<ߋ/X	���q��!��M�{},�M������:i>~�}q���K��"�>#��?�tkk@�߹M�l���R�7g�"X���
�ኻ9u y8��c%��M,M�8�@�N��iN9'0�1�y�������a�ű �qqf��ͻ~�[�X�zp��43D� ���՗()�u676�`��2��6�Nh�B�U ��z��o��P���r�n�����S��ay�~q)z�T�ռ�������׷ܻ�h��!=u.@|�L)2{q��k?h#.xK'�E8E�ݧ�xK|�]*1��{���k��»��;���̻�I`,�T��S�s �yӝw�zU��[�=�]����U'+B��>�2�Ø0��v���!�ۯ���y��k���@���Cbj~"�_�?��:�̙o�Z�E�^ o&�����
{-X�ЩM&��=␎o��������/vhg�5�}(kz\�gd�G��]^��v���uy��.���)`M�* ,1�m�9��=��׀ʄuu��� �p����m���"}O�%u���c]�Ǧ��5���N��q�O�xe�� "O]��֒h�L$ ��>��s����!�� �!�Ub�!g�"�O �Om)�0��)c+U]&��[��x���g)�4g��w�c����_l��o/�~J!�-ߵ��n�{[{s��$��ŗ�}ma��Х�Y7�z''����sR����߽9�A9�,	\i6�칿L�O~>��8��|��
+Z��)�'a���������T����--��MP�b��B9l����c��y@�i����I��z+l5�Ǔ�^����%��`����\r�XZ' ��`*朥Y^Mii�Qҳ���1�Ù�X�Z𨭧��\ن��]k�N���q���QT�D���@�t2	8^g������MA+��"!ZE�Sz����<}�~1;t�&~^yw��o�z�0�
�DR�^߸q`�ʶ�s�J��<�Ԕk:w��l�Ӵ.8��N7-3�xR�K@/B���Sz�?�O>��>��sv{����{oh��* `�(�42�Lf����D+|�_o	^�z�+1 WHҲ���z�j�^�|㶗�����]ks���p��a�ge��'>_z`�,)t����V	�]V��� ���vY*4hN�����y+�$J���� �w�W��J��o
����:�暷��}-l�W�d�M=��8OK㎯]��W�b�/��6���ij��T��fO���_Ȕ � u�=%�Sx�d����k�D �Ӗ.g�;O���T�<@��=��� <3 0\�%ɬ(��L���o`-�R������o;ɳ�y�Ǽ-J�O�\��6�k����Ϧ㪋g��֘{-�}ip����m�pT8���<�U�P9�i���ݠ���g���*�mH�S�|�dPcB-I~al@�����ҍߎG`8������~�� L`d��lt��_|�}��	k�^M^Ep�ς�ʝ᭿pu-C�M�^�Ё����A~ptH�;~P�lѠ"��2����lF��fB��������10E�͌����2�BY��A�F���3�/���v�h�n҃�k��a>�{휲��U��s�I�׫s}~D���}o�4\B	V�z�w���EA�_�v��ͩ8�=��}��m��xB/_!&�K�����~��K�c����m�(d�4u���pFO�y���x�L�]:m�Ҏ��'�Z�j��8��b�
��[)�+.���%������4��	ѷ/��'/�=q��s�M~���]����T�lH� ^.~q��{e�����8v �Y�o9��i�bޙ��<������딛�����֦4�O��w�5M�]B���ݖ�T𲢥l����KW�� �	�cNp���k����-C���������~�B�"*�E�Ϥ�9T������3�pc:-5������� ��eA����,URH�ݳ&���a�D���~��l�a�d ߻����e�`�b�1@Q���������y�_�k�/څ���pe��1��!K���[�#�y������9�õ����_��G=�.���I}=>��]���x[nۮ�����M�Z X�����oE%@-,���Sw(��r�v�R.� L�c���p	���ш��Ʃ��	B�I�T�b��
m�2�����p0҂�>�Q��M���-fJ��J����Kr�M�M�q�6ݹ{�ݡ��)�&�g( ����3�]p2��f��%���w`��R�����_� �" ��c:s�d�r��L��7���ER���c����~:
�M��y�+�^�u��ڤLf� ՉvM]��hB;;{<����oؒfx�^�e�u����jA\Cz׍������Q�����u;~=�E*$G�S8_F�	�Xͻ|��>g~��R2[�t4u��!ὃC���d� [��/�㇃��̈Ǘ�& {,x�*�<�c߈ цǄ�W�9���P�H��χ]�@��yҒ򄚠��{�p�ʪ�޿�{�γ��1r\j����je�;W�r}<��+]�r�H��8_jOR�YX����.4JNh�@>��q���[��?�zY�S��$���ڏ��(����Ȕ 1`%�  �TɁ|ȑ>�*9�l���ٍX�µ����$yv�xN��E3~�/6��d8�w��8^�b���R���ϗ�w�1��y�E9�Vn�6�):�iw���:}�FmJ�u����T[	D"3�$[�<��!�����b 9P�$�(���$����tb�d��3�-b4����{ _LXLHLf�c�}��L�ѐ�y�ݻw����%[SD��a޽x6�u�n9����4w fk�&�n�:&�K;��7�0x�E�[b+��-�������{�9��Vv�	��OV:������aMi:����v)����*ꨭ��5�&�ޜpV��U�ՙѤ�`-4��e7��ȿ���x�z������`��z��nB+sD�1Qc���8����#���H�J�/�&c܊ �{�!#8'��q��x�vE�r̗�\֏y��W'p9�C��E��� �E�Ja!<n\�&؁9�@�4�b�õ��'�+����|jJ-[�[NH:I�T��IM]��5���Q
`�ʩ%0���ɜ�e��Zo�S'[J�CyhY<�EK?��QGp���͋�/^��~z�
.|�n�y�B�H٠�Zy�DX����1 ��_XBa����u��y�����k��ׄ��ѣG���w\_���v^@N�#lRU�L����n�⺭���tk �A� �u ��5@}� �<�O�C��wȳ�@$o�ry���|p���4�w�k�[ڷW
 'S�PxF���/�iNJ��/���8�f^O �g#8a �i�&�� �$(F�&⮛�HRF�	z�m���~� u����f�5-fc��"4}N�9 {px�O|ׁg�۷n������g�����0�v��Ig�������K��9�m�h����`����*���
Y\��m.��n6&(z;�j��oYZ��'_:Ъc���:�[a�Y�Xov������?GGS:O�ئ�a�>�ӿy ���ʻ���{bl�$M<?Vt��6�K����j����$&$�+�\d%�V�p:��J�NU�&�Ե����-6��d6=x��+�f Wv��ǉ�L�|9��	 ���Ut=צԲ���i}�.g1H-���CX\X���b���T�ͭc�Xs���.�w@�*�EH�K��浄���������d>WB]�<��Zo�N���C� ���(Ʋ�"
  (������EU��J�h��<]@.Chܖ�Z��gƦ���צ$BI}`�i��M�g�><�3���:Oj���+J�u="Re�EQ�J�FW
 {
���~[�q9����ؔP�������>��U����q�&��V:�H&.&!j�!==��نI-.���'��|�qÏ�{�zN��~���|��q ���i�o�z���"	�Ё�>x���]z��K[��s�^�z���4��v�h�
���+桜ʀ�� � ׬��uy�RqE�1%��(0�6��u)S�(�(E�f$
çd:��11fڂ���o�:].e�	��V��xEE�j��-����U��.�x�/,�Xo���T�7��K�x\�F�	őc�-��EPƇ�.^^��PՃ]_ne��_�g�O'4�,����pG�}�.�RLy��l�wm�)�0Ǖ�OUU���çg�Lp����ySwoå�B�E!_]�ː�!�
]әSS@���k:{���4۫����Z�Nٚ�識�Z��sw����:iPp�
�	dG��a�\VZ��X�$�
���L
a�KmR+`^Ar�$���m��7�8glxf��@��}A�'~GA6�,.�(�$J��\Og@�.RX$_5�R 8�x��p�r �"�q�#'e�!��x�gr �������@��1����N$ u1 @����"!��mç���J<r�h~����;��<z���q������+�{�M;��R8s'��������`���}@w���[�is0���fn�'�[�"�~��\�^�O�|2�I�Ϯ�w����%��s҂�*\���I, L ���F#:Y��H��h�Q���"��{u�U��'i�(��;�-ߥX��ɀ�ƻ4� g������>��D�OQ|����.�G �����bJv>ew�;�_x@k!D�},0־�$��+W�9a8�o�/�e��� ��:�|O qkk%�.���}�F%vjy����k��f]G�=���Z����v�v�V�u��Z:�\Hm��ے������|�s���ߛ�i�����o�5�� �~�� wv�Y���0s���9��)ȍ��	�@�|'q��G���E��k+-΢(��d���,��VZ�}�`�7�UNK����\����א2� �z�"��<Xڼ7΋�£�Rvi[��m�9�2 �ٖ��׃VN�d�U�Ґ-K�X� f<X� ��m�P؁Md�xf�<-�ә�`L@���ӟ��~����pY�(����W��<e�c�� M��}I�~��z����`�snv�	�'���D��wާ[nb���x�'=���1,���Tk��yc�hOr�		Ьς�aQ���q�����ڍ9#G&X��`lm5q�� s���c�����	�7MA^bO�#U��B��{��D�2@��4s���Y�
�1��/�g൶��ϡ�����l����m��Zx�U�1 L?�|�9$!�j����J<�$���x���ݻ/������w��ir�B�l�=���2�9~8��·����ܵ�!f��ܹ3��PqJ7P��M�&z�����vp�.u�m�z�j���S!V�mo�v}�.�~`�T}ϓ�d���K�b���Y��\V��䷋���w�y�����ơiI�t9F@�: C���)��ϰ��&e|�"�8ח�*�`\ {{Ǘ
Kp�k������ ���2p��8h#�(%w��'��K_�xN;xfIF+����<�hK�70���� ��xf�P��=��V}��H�x_ ,E�[� ����d<���7��ь67 �zl��q_�qz,��j�:;�1���E�X�M',�l"�8�Ѫ$I4Y��ЮIZvh���	ȵ�H�I,`4�AYѨo��:��ä�d��I�
/�����o�X\�:/�P?��=��@y�h&W�.�F@p}��t�A9X��B��L��7���������k ����|MBB����}����w������̍�J�4�q��� *˫F� ��_NG��{��>����W��s�.�E�l�_��쳺��޽K=�g��i�7@%�[y������L�O�~�9��,���&dm��|/>>��5Q5'�ANP]�lWǗ�Y�-u�&�Ϳk�������k�/�^�����{7�7q<B566�4����
.
�Qρ06E9UZ�[�m c<�"���	~3O���HζG��t8��Ԁ����֜״>u��hK���\�.9����6�ں���6	��~�� N�u܆��mr��9���������E�°u~�̙]O��WC�j�c�����;�k�[�Ԩ���ZR�gۘi���ƭT�ȑ��	C
 �v�=��� �ÃC�s9C4H�� T*�Ցm�|w��BR���_������t��ͥ2Si���S��tVh�� ���d�|�Z��y�uxH*�^ �J�6�L鱬�e���,�8��u@����M 5���	TP�� �d��=�R{���a� 0�';�oi�Lg0/���t�����
�Flk����F!�C �^$&�u����ʙ�%^�c?��C�	���A��ۿ�Ѡg���-�����}X��1�`���;��Bs���l�\�Q2����n�s.���Pv����T �`5�4�E#�I��4�%1�,�Vb�������vv���;w��{��chP@x���'lkw`Ǭ�67�q���m�F�*�)�<x ��CO p ��z\��WU�ٷ�q�"C7"hN W>��h�����I5 nvw�M�f�������
��܍I���c��:Aײ�;�W���R�lS�A�YW��J#�e��1����A��dLx��C?����<#�w�����j��e!N�Lc��0�<s�Q�%�X|�����=����2G��}��5rsnĮi�V��U���^��3�cXIT�Bl-�@����[g� �Λ}�۟:\��;���O�����z��eYX�%\��^�����tvd�+�0$�J�%�E]�㪿�~ρ�Ԓ�*X��9����u	w�6��Y<���1x�糽���m�K{�p���D	���NJ�מy٭X�[�ri�l���냏ԕ<��	����W��/�B ��3v��(%|p�I p����"��7���`�Y����)+��,��*��U����Z��-	� JA��}����5l����5@I�0H�L�0�����E�rⅥ����s��)7�u���P�ą\��i�PZo��q:�RET�{��� X��j Jn0`�9[^�>b ��h�����N�
1�>�(�����̝ 5w`��8`���a92�<6��6wL6/��p�5Wz �q;���̧��]c�A�?~��I���
<�Д�ā1\ſ7]W�r�7�3n���M{V$�Ae��	I�F���C2&�E�.~��gl	�^>��s5 ~� jÁ�p��	p?���	a^,�E���/�R(�Fl1�,]"��,�e��p�-�W(�ʻ�v����c�qa�~!9p}���ۯ�i2�n�*;y�V��۲t�Yf!�S�h�ny������?C�]�:��f���&���	�W��в��J	��iR��Sb�x�/g�m9������ߣ�w,�����hc�����Y���B`�������U�4���� �aVP�''�ݢ�����^��u�А>��}��s��> ��Ap,l�H�t�����δ�
[�`�F9!M߿�8�{��-� �ϗ�n䮟>G�s��1��c��{��g����.Z�YV��g����V�N�A��O&�����rYc� ���j��R��'�g�g��*
+%���]��_��@dq/ƽ`��ۏ�l�<9 ��N�q�Rb��׸7�.ؒ��M� �����������bU_�}(���ߟ�&m���A�����Q(Y�����<^�����6���K:֗���� ������'g�:ķp�v<�қ�*Q��<��(F@�� TUAsl�67�+h�����L�[SP7�,y BP=�
~��_r,0@+�	��`���W<��� � �����>7�������l�s�1
��{�����{�QigwFo��T����LN�:�'��E��Mt��aH��T���=4�����;}��O����l)XG;�/���z���.ď�}�.4Z��X��#���h����4�(��s��xC,HGG����s�����w�z	���a|��]�i��B��y�"�kǍ��P�@��R�,�O	+#�R3÷�}ͳE|uK+��,x�P��޽&A�zE� f��ZҲ�u�Lm��}�/���f�>��=�WQϠ���~ߚ�mL����\����S�W���7��sB�s�Wh�˳��7o�N(q๿E�ߡ����~�������_�ŗϸ�]H�� ��3]�qH���ڦ"Pi��..��`��J͜�ZQ��XdWY_s��ka��v��Wlc
Hs�w=Cڞ���Br.��m�x$�jSZ��]J�?ʁ���RT�N��s-�e���ڦ��}��!��E
xo=�T�N0�:+3�8�i�� Py>��\x�B!�2���O������"��Y`yF���������i�JD�yf��cG�$<�q�]�K��=�9b�ZGF?	i��n��D˧�<���*T�`=�:�� ��Bɐ�e2�q ĺ	�8��e��¼w�\0@�۳O��IsR-����酧��[��&Iv9�:CÄ�&/M'3`y��-���Lg>�����D�1�U5c�(^�)-Ao7�-h����\Ɇ��/�-��q���^|Պ�����{�#�_�������d��+d��If�d��*��t���n���I^ˉ����$Lb��2��"����-b6� O&c�������/_����.�`�U^?V ���C���=d���满�	=_f ��!zZ$���9�O^����9��&��k��o~O�7k�B�JL-����rss�.ܸ\L�"	�bή� �8�,zl�_��b����L�u�-=�К�0����9��H��u�`��&�p�zK�{�	e��y�ڵ���sw}.�d1���6ڵ2�Z�*b=�>qQL�wX��aZ��b�sr��ͅx��b�߫�vS	�M�6�+��khu�� ��V2{vV��]�����16�����s��$Z p�2"7V��(�� �� DR��b0$ i����_�0 �H�hk��Fh��5�:ɻ��� ������[sV���穨J��) �^^�J�6>����5��f}?ݶt��V�7��
 `Չ�v/tI�r�_[�pvh��Ć���_x9!��/��3�m�JGi�$�M���"���dB0�<��W�bp�\L<X&�Q���m��'���o�`�GwoÝw�@��x�]{{� �8��?xC�Eρ�;.������T[~����1�4����"���_�[�K��<�d�cx umk��	e�h�C׿\�m�g����]�(�~E=���{�K���˪d�Jo-��)�1��:����l�=��j�����]ӗ�<�*��9��&�f�����f@p�P+��6�}rjdMb����!��MܪK[g����h^%t�3���NKM�w �#�Mvi|��
��٠��r�=�j�zdBp���ʯ��fn^B���2b�������`S�y+��yŔ��'���&���oV����q��`������6�y���<	<	��1�,H\� ��U(�T��m`*|�����oi)�N�{�Z˼���YwS �hW���i�\9ު�I�΂�r$g��[g)���*�q����2P�kA�gmH��١�[܃P�myӖ�U�E�:�b��� �F#�� �z��%	 F_��x6<#��R�)�9����x[�R_§�w`l�M�n\��u�Q�Ա�z�׼ @�L��  J�}��!�Td�H^0��Ja.�@`!��k��S[�M��A�ϴ�+&���d��Ϙ�Ϟ=#)ƍI.q=����3 X�� < Mt�7a��p���p� �M�-ߦt�_p�c���zCI�d�Kf:��٧�-5�����,x��Z�,��L�Ȅ�g	}E,B�-\��PBR0[����V�*<��5`��9_מ�D�tB![�ocH���i�5W� 0���B��TU�ӛ��u�(+�ف��4C4z�߯i=��7�p��-����|�E������x�v���u� �ێ܆��^��;�>[q��9������"�3 ��՛�C��s�6j�#1���mh��;��Zϯ-2�O��{ ��=zx�f�N8;��=����%�\���5�&m5�n�"�b�Bb�X� ��ڛ9ˉ��k�����*��1m��v��N۾�x�
��,K]��ܷ�s��*��y��]�4��|U2� �K(� ؆�Ds�1�6V�9z�J&�y�hKZzip'�1�I,�8OJ�B6�.����z�g��&�s��'���X6(���{�F>FM^"�ʛ�w�x��Z ��/~��O����ϟ��H�����Վ+�A	��.�����V�Bp?��K,zӗ7T�O5�����bA(����K/~�$�@����ѣG<�	C�\Ľ��'4�i0�t@v��n�s/߻w�a%)�` z}�b�x�u<t�yH7o�=f@���� ��ik��N@Kt&@'$���[x�"3R�w/�mL;�m����h4t�ޏ��2X($yD��,|�u?˽l(��As��Ƴ�\>F�ONb������#����po�v���E�K��e�=C@{N��u�y��JQ=���3�+�cŃ%@��n��θ.p�1�NP�P�usc<]p���/��W��9v ����PL�F=z�����m�����+Y�+s�����痮�j�
'$���������O;o�����9^�h�x�tM�'�<E�Ԕ�^�&����2v�����믿fA��B]BjΪ�v���J}���e"g����f���i_�u��*��#�"�߳�?��g$�F��ƿ���b�_z:s�p�(��XgM�q
�|��3 3����M���}R� ���7,� $h��Vܔe���N��MI��ªp���\%���2d�:oK�ϲ|��.�3⺸'����Uʪ��yzj4�b��5w�pK��M����? ���>���?��?��c��]�C�$^Dȏ������駟��,����6�X+��b �jˤ��2C5�9�F�`^��9+Q�S�w�_�I�[ѭB�:c�A�WL2��߰������6=���`w8	֛�#����v����� ȪZQ`Y0����1�	�+���
�mo�"v���҃P���d��Uqڵ��҂��n�0�!eQ��d�ELO����Â�ݭm�{���|�p����_���ZHQ�5F��lT�$��c߹_������kn����C��򓤛J�r��['mk�Ӽ���� {ҫ�)��t���֡�Z��KOU?sB��9����7Vg7~�
�*�Hېx�ߨ��X��ѷ�w���=��ٞ����S���U�`:�����{}�6�\Z0�-LWa^������I����x�>��F��]J��M�eps;)i$��]���=�.�/��"d�?�����s�>����,�����M�V�޹����}i{��_���s�g����ڒ-���uǦ^����r��<�ڜ�c��[���#��p���U(}������ǅ�cI��`����I]\Ȍ\&�ڨ�O�P��Y�V)ud�`~K�/�7]�kA=eX��?�<�}"�׀�+	=�B�/x
x�<�$�J��Y`1���6�k��B�o���4�P���=�!Q���3�;��"���9�����{�g�g��������Y�YH)P�`�`�A��M�d��+�X��� �I�s�/5��J�6��M�0�����Ms��sM2�Ⅱ|,�p� �Z�?�����sr��!O�<��ј�_�8���نQ؈�����a>s�0N�ƶc2n�,���* ���P���]��Z �y��A��T9�x��\8�@{A��|lx�ʆ,��g�k�7ઝ�DQ�;W,\�g(�;�f���ص����ņ�J��Z��NU�v��XG�hmN��qkN�׈j"���ߣt�Ң2��T����2��X������]hJ��ۺ��F�����krns���L�9 �52�LU���	�b_U��P�hw����z�m{�whhZ���w��+N��:�}���׻t�<6n҃����f%��Ex
��W ��*|��MO6�p^��GI�x_�5�-�T�Y
Xr-#����9-P� ���l	�R����=�_ �s�N�pma��Ӥ'��Z�ڡ���8���w�����O��n��@pW�׍�ӂ�s���Frr����Ӷ{g�省��}�h%��<�F�(�"lU��
���KQSѦ����ߍ�� ��v�$�]*�I��:�~=/u�q)> u����o�%�3�0���I��.u��-��j�O{b�%x0%�)
����f�
��� Ck���V��c�����!B�$��Ⴧ���}�>���L�l`��7�α/���?�L�Xs0�G��h]�Om�v p�R�c��4�j�`�i����`�yMB���A�IML�x������I�e�	 #.����=�� �b���w��5,AxU�������������{��1��H'ٖ������W�%Ҥ�c��w�q�o?�]�B0awf�i���,�ѡPOE�6�U=<4��fC�'�'��������g�Pu�x	-��[�gS1�嘂־���m�Ne��>T�M�B��LK�A�6g�6�1-�����lJ[(�S%�	PY��P6�0�4PU(^�߹��Ὑ޷Jj��ylލ�Y�Yt��8��z��W�� K[�?�uEnߟ��4&�
z�f@o��4�[�v	��9�z��e���ɀ^�9�;{��ݹ�%�L9q[ �TY�)����=w���Db���s�����6�I���hM��JW	|A����6��NCC���N�u��O?e��
������y���x�y
�tӾ�P���tH�۶�Eu�&�Z�C�N��!4%$�i��'��3�Ƕ�&�3}��H+�m<ǐ~Φ�Oϧz������EFm��.5ߴ�t�yF|�9��X7�i��
�H����4�VH)u$ɼĲWZ)u$@H�^��Y�mZ�  ���.Щ�t�{_&5���J�*�DQ&Ϗ��G\�D�ܵ&&3�	�TI�� �Q��J91���G�H�
�gS˴L>���f���a�N�p�e��Z0�\h.�:��E��3��g>#pF%,�cz�G����X&�B���4�����U�����A5�ù/Ff����Ib���~�� E�&M;Ủcz3ͨ2��|��ɂ%,�q9� �	��3�x����鋔g\:�.b9ν�^��T�Z=]� �ܴ�ث�,Mu��9�U�A��"F\���#����$�.ꄢy
���~�O-�9>u|�
�w8�k��ب6a= ����������iwg�[ �J)�����Ь��pI��1x���"���_��E{��l�<���I�e�E���Zz�^ik�,�US��;���KnMP����` �v��S�@�V�#<`��o]TY��|[�Q�VP��X?��sUي5��i�6/����C�u$�s ��rK0�h����W�1@�X~�j,e�����xԥ5�WM�n�~ sR�4�\�H�ڰ. ���!)ߨ�斵}��A�.��0�?��9�z��i���O�/ź��])���"B6������c����_���o��$A�(�6�L=_:n( n�͝:5l���*�f��3F�--o���@�%"i�APyq3$9x<�C�y7��?NY�X�*K�	�K�pJK�ϝ�t1Ғ�i����4�њM�>�_aQ�Zs%XD-62�e	���X���d�n$&�0\���A]{�Q�]T+~���-��bZ1�-ރK�_t���.O`���Ҭ�� �
� \�>c�g ��Ge>c:^l���N�y%>�k�R�
����P�;k|�nquy� =)B飰F�~�
F��FK�<�̗�;��V���8b�j���R�L���e��<��6�y��=���1��u��
,�u�/uw���Qjq���y����|Sˠ|k��_ ׁ��]���7�P4��H�>��0릺��D�W|���8T9�c�TBA�>�l���~�l�J�M��, ���
 ����|�~o��X' �v6�k���(��:�|���9�8 �{�<(C����O.�H{1ס\E�5�^����3�?����jݔ�KӍ�"����o�_�.�d��4kZ(A�Ab�^bA�$���F����B�g��JLb��j��Ĕ�֬��v���x� �^Ft������q�T1-Ƞ�!F%��(3g�-U��亾R�La8r)��3Ԏ�dc��|b���3Ro��1f����m�g�^�h��Pٖ����J�c�JI�����ҕR�zÜ�)�v��gB>�ߐ�*'���8@+1�,L(G�n���ii0и���n�Qa��[�����I�?�G��3.� �MP�� Í�`oQvK�^�9����	X�N�Ox�/����C�"�^L��
�A�Y�5�n�o���-ˀL,^�����w�<u^�%2-@ ,ָXv�@R'��7�", ��$P���=Z�.�M�*���]��c�x�y�����~Yʋ��`�2�f�������+��)����qrD��?�3��k�����k��������
�-�q��H��n ^5���U�뛩���',��v�6�SW'���+���*��(�Qn��
��6����3�۲o5��`ͱ��@$.ːXLD�����|	$,.��N�î�y'�l���j��rH�%�,$	<����7w�m'��E�p\�y�KhZ�sr��j�;ʊ{J�k)õZ�R�!Z0��}�
�L�j�+_��t�@d�^!gԜ���0� �x��鼵ѥ�v�u��P�{���	u=���.��ߦw�hw�k��(_�� ��66�~�s�R����14�Dg�!7��	Қ������	L�R�t^z=(�
�?�\�+�FXfI�RkXZ�ޖ�>��k,c��c�(-\Vv���=	�	r��,����c�$�M���wqE���@b	�e$�ؤ�h��G�>(�`����X��RpsY�)��^vΧל������v�-ᷔQmK��\<�+0,���g�kH���=�o��P��#	�a������ϰ�C!�ϛ��mt� ���63�e)���>}!i��-�Čل)�@*�s��J��-�ԭl7곕�_��Ub$q�9.R�$��OH4���[�n�$������1�\�q��>�!��qC����]�wi©��8d!f[�GM��%���]�E{<:F�u�h�^B/S�7y�	3y��[�TSZ�m��^Κ�� �6�a��nql�s�wg��ԣ��m���W�Oh8*|VzSЖ[��n��vig������p�*�c�+������m%'�B��-�؞�c:9;�kh��
�}wݢ����VC��%.����A��W��KZ"��� ���
��[��u�`=톫�# X���"��}���,�����ʎ����bnL�m�3[^X�?�+�.z�*�I�8?����=�t�
�H)�Zi���̆w��l�{pj��*+���k.,��o������c��a�e����g�LԜ�iU�*���u{�4�媯�ג��Z�dU&T�b�_b��D��#@i[�!s���g�}F��/��Q- .�xO�XKI,Xy����;�ߟ��=�pq����k���q�i1�aщ�ЛR��C��?��I'�9U�l �Yp��$P��"`X��6��S�lm}��	��7�����`�H�&f�E�]�A��Lk���t_F@��d� ����v����q±�W�v{~3%$�b�kڱ��/ ���rW;�n}� cb�5��צ>�,�~t��ߍl�僜`yF�����[z���\׮�M��YZs��%�I�ⴊ�i~�s���~���{�=2�Vi5�� �,fK���}٭!dy�6w ���G <�6X�w�{n�m���e��^NǧH�a�������p��{�C�86����38�o���E�uėn�u�,����+z��z/X�)���wcr_	i�)�r�u �K=zD<��$���}Ͳ ˵��� �	L	��g�g��k�@�,��wL��V����}��?����>NM�jKec��As�'}�Y�!�ˤZ_M�_C	���E��"4*wM\h�UQ[��n��K���+|!������{��o�ėP�}�&�o��q���;HB:e�dJVo�������K���Gv}F�$�+`�I�/���pyF�/_�]^��bT����\��= &KK�ss;�
xDӋL�Sk_k.�6��ez��Je[��:����/jۺ�LF�a���Ip��g��Q���	B���h�^�6�������X���o���?g7,&�UH�mG��Q[��� �@����٦���nllz-*�C���Z�������m�%'�SYd��I|��vh�-��C
��؟�k��j�������v�4��W_�����;.o��/�a���,�o��4�]F9�Z)����X����9��L.��|�Q��_�-��v�(s3o�za���+�z��@ �:�fp���6�=��pw�����[�76`1�����7��Q�a�] l������9�[Гg��������G~AY�	�<�W3��5)��/6�_8x`�AI?�s�p9�������\F�o���
[D��G�� �y�����&�ۓZlS ��u,�l����?���]�V���b��f��X���|E�J���~--3�40����U�/��Z�I�ba��~��_��<-յ��\%IokZ�u��US��/����5�u�d�O=H���8�%@
X{a����~G��կX�xa��Hr��?������+���\�Y�J� �tn��6?���/���.O>jb4���D�f��&K�	�;���
.7'�"Ԝ�y%���!�?�*����u�dp� ���[o�k`9��ߪ�&��pE�+6,�$���K��eQ�ǀ���=X<�61�p�2��"tm�֘��GN��iYi��~F�}R-|�][��>k�/��q�D��J �� .�	�.�;�|��>�I<�b
d�K��י�Xm����r���Ҽ�WG`פ�����X'���^�ݲ���x	!\ �ww��Ջ���ľ�[Ʈ�NV�w2=���������q�^�X˝�6��� �9iVf�5Jo��:<���^�7�>��~��;w��Wr}A��d�.��SZ��x���!	M ~q,�ؠ��p#Bd��q��2Bb��Y`��\�,�վy@�?�d믷q�5�M1�iY�x���,��[�Y���/mH-Jm�L�z���9d��Vx�|N�[T�$��E�m�� �/B��[C�.���[2�X���5Y �����"�z�
h�L�˒�bm��M�Wj>����$�_lPt�� ��kvy�u}!�$,�pu�q�RZO,��G:�]�{���� �D�T���7�ޝ�N�x��67<�BbC2
�>�`8� |*'�鰠	�?����^�zI�Go}}`�3)/�2n�5H��.�0����+��_���RL]^"���)2F��zK���F,�{��ӣGp�ދBPƉ�:,,�n�ƾ,��˚��03 �I� ��=���g��W�ϟq|nQL�r!7J 7�]^ɋ�Y^��8܆������|��M7��Y�o�VE���:����2��˳eϑ>�6�y�x��	:��>v�xB^��+�;j��ɩ�ahw�d��=�;�Z�. 4 ,8e8��ݤ��Aݬ�֜q�wD?����������۟��󷴻�еͰX|�t~�T��
e�����'V`ª�wzz���"��K�#��M�Ԁ�<$���\O'�i��e�oMb��-(�kЦV�Y�P������O�6kNs�((lWoIL�<���O�8��TB�Eȿ?�vy��+c�&hEq^=��Sc��	��T��k� ���kW������6d��~��1����BĆ
8��(Y���2Oq��7�nǼ����_F��<���:Ӽ��w�Y�e�I0�c<���෿�-˪ �P���C��
s�'��������������s����P�|�1�JF�&�����[ ɐĬ]5�V`�6{t������_~����v@��K���#�&df \���O���&[ON ~�������#_�����5������nk1��1�� ��� ٖ�d�41��HC��ڸ��M��s�׻[B Ł_��9��[d�n�39w�gG@0I��h
=*� x�)�����/,?�}<����au��f,�p*���rtc�駟�}�^遗M��nb����tK���~�W>��Y$^>L �w2q�gP������Yѓg}�v��-9�����Uڽ�
�Vddn����� ٢�Po8���6ŕ��k+�tY5q�������۟���=y����6�p<M	k�S�zK�*=�v�6�-h��� ؀���^�(S+�y�ɲ�vMN�>A�L/k��g�j:g!��^)�m��΍��9��vɽ[��ݦ��ڬb�I}6��y��U[w�Q#���h�	����B��)�%� p�%�Wdtpк� }������*)]CMkJd���.�WY�9��m1����3������f��A1~�q ���|%)b|����o���M��|�}�Q$V_�!!J>��y�Ƀ�D� �v9�iMsQ��.��p)�Ȼb௻w���F�w_�?��?���<����	��`�	w B��rr�<�t@n�]��	}�������n{F��|g!�4\�|���4��t77{,8�K���K����/�6-y�{Iy�
�ّ-����!3�	��Ҟ�[�z���^r���>��0 ����\ЖY]ȗjlZ`I�;h��J���M�R1�h#��յ]� ��*�%C��,�e�O&'�$B�;�����������g��j{�m�=NvŖ[C���e4��V�y���\�U��{��%5��lȱ������'�ӓ���k:����v�y��u٭���6�yIx���,�� Т^#�Ԇ-�>W��&�,����
�:[��g$�NjE��k�m��<�xѶ���V��䝹��Hr����Cm��6��j�?�M�D�gi����k�+9��֮�%���uW�m���^C:�X�z\&I�`U˯�j�A�'6YSW$<���P����:��:-�B��4 �sS�w�$�{�Ϙ���k��E��=��x�Z�A�k/�����˾O�����yOO$���'��0���Z�|?�ƿ�bO���;L)�f輮= �s~;�TM������.�<7E'��NL�nR|�����nB�@���Pú�8&���,���b�6�5��2]N3v���������b��d�_�`&�޾:���]���U���&\���8>	[���� T�c�>���@�s$�kƈ|m����k���(��K%٤OӾ�=����Fi|� �x ��6zX����H۴�eӞ�w����J�3�����Z�>8s 3��o���o~v/�hk�� �۶7X9SZ� 	��$b��������Bt��y5'E@ HGtt4�7o�����������)���{���5���29��{c�n�<Z������X�M>%��,���,���aYJ��"Vɶ����v5��6+���e=����c���U�I���ݫ��k�^��_�*��l����W��|N]Q5Ѐ�*��OĽY�_ G�"�L@$���r<x�$=Պ�����媺L�K1�k��lS8���B`����_��3�<��Y�A�j�ʌICN��ң�r��"eP�|ƹ�#�@6h�/��F�Zr��t���Z�Ey�Sئ�
��]2��_�f�;O
�7`�=�'�Xu���&�0�뭥��l6���^�p�]9�V����ǖ����Yr�WN�,�b�����j`K?ū����=�g���:Ī ɮ@M�>��_�̰B�j1V�^��bc���:ѵ6�s�����%���[M�l[����K����ۨ�Z'˰�M��Q�\e�W�.�߻�w���M����~[�w���E5n7��R�;�}`�E���s�^�ٞ9�|a��ѐ���)��/߆�ݺ��>D#��Z��TL|V{ΡG���"U��k����Uw4,_�����	���1&��Y�ym�W(�|'��I��
�zb5>�]�$+���|�Y�R�m�p�fqm;O�+1��I���}R����gM-ߩ���Z҅ΛF�~�,�~����;\'����I���g�5�~8i�g�
7<IY����~^���Ε��<�R��e���bC{$9@xx� J�`<�gP�IX�&�Iʗ�\�ު�Y4�� �;	��eח��r�c�Z�����Ή� |%�[��\����Y�;� �j,��A�.���A���7�|�Y��m�y �v����v�w 'O��ob5��d�%��&���<C[h�R1�u-���j���?�o��(�b��²���u ��Yְu8S4g2�����7�	<��-+J17G����mѝ�{���q�q,�cU'�Ī�M�M �wߒNNQ��3�L�5�u�}��][A��MuC��U�#<.^����� Π53qy`m9�	/��(�PbC���Ck��E�f�^g�>����ފ\�*i����l�`"{�[����	Ӻ�,��3U�M��K~A�~}��pH7�l��%\�/$]��m�5�s�������-�����r<�+:9�����ŋͯ'�f`>��s[�<��T�L�N�P��A�#۽_��㑥�ȫ��=�.�{�H-~4��k�I�A�7~L/�4`kHʯ����6�.U���gY����K�D��z�5S����Jy��%�MʁYV�����d�>^��ݼmj�������R��������`ų�����5̔��sו�^��1�Z�KJ_���b���wc$��S��uST���/� E,s؏�O�e�E��M�`���$>��(�R7m�h��oq�뢀����F�Lfy���Di)sh/�"X��7��-����+�ۿ�[s1fڛӘ*��+�2��9y��ޔe]���=8Л�o�����m^b� %7�v �"�AIfB�&V�`||��g82
ų��rrӬ����H���]%�
�D��b�o�[p�g�ݗ�d{y���l��u�����	��qIZJ�6
��Zo��I���}��_��>����r=�r2��dz��e���A��]$��������۟�ǟ�9A��#�u�5Lz]�:��/�Tc&U��O�Sm��E,�|L�U@8ܿ����G�
��`U�6�6�I�=�/�E�Ld��>^�U�]
LtE��Ib�ţ�ߧ?|@�~�����n܆n�
6Z��[��N�/�-M�{1駟��_��5�������l���4Βw�<˙ f[z���/ɻ�_���.'��ݖuz�s���m,�v���e���0�㐍�J�"�G��,}�2��(�,X�	��K��r�C��%A�F1�2�����$=�i$���7�ˢ���Q�ɗ��)�_Ĳ��Ʀs�}b	�Iw��Z���i]S}��Ԃ�g�I�����E͕t�e��Ԥh�[(�K���tX��(-��!ǀ��6��n����ڱ��$T�ȱ��hU��U��q�XC �Hx���	n�hc�p�� �G}�.� и� P�Xȅ�k���ϽHh�$/ų�� ��)]g��&�X���-=w]c�˲��Pj�ڋ�� ����ͺ޻-����6�9qio��\��o7��1��	 ��#ʕ��l�:-k� `P�A�΄�b���R�y���<��iF��n�����-7Q�E��@h��`���I�Ƒ��V0��`��:(ed��' �H~5 Ԭ��HF��`@�&U�ܣҍ�Q=�RB;g������&}���w_|H[n_���m�|/�Nd�H�_@�~����d4�w���#:e-���X�@f����EHӯ!��0�i�m<F\�EK�`ù�S@)�H�b-�����h�e��m��bs�G���Ч=���O���m�O�ry L���֖*�Y���{4g��̀�����Cv���^����$���T��E��������sV��˃��r]`�����O��V(�u�<9Y��R� �� �M�W,�����5�����L���+=�e�	�z����ޜ�$���䉲2�4��>���
�M��Y\z�y���4:� �-MBo�n�u�6�<���,��Z�VAS�hC��Y�D!�z�ͣ��3�O�L�5����ky��5�uBAh�.@z��uVU��_ɚ�^Xp�� Ed��۳�7]
J�E�<`F�ד����|�v����y�I�/�S,���q�T=����|6��u[�}����$������:�PE��³�6�L���s+xװ唢G�r�%�G7 +26����^4�6*�mV}��Nt��_��FA  h�yXAc��[��hŐLB���|b�]�: ���L�����|�!���w�=vL�5��!�B߈��nb�(p���d����ݨ%1����t%@�,����ڤ�ݜ�w����^H���5G� �2'o� ޤ��6�,���6�DG[2�4����eJtϼ�.t����f���o�{�w����n�ܘ�C7:��`��Kt��� �eRȸlw������=�c��̧/��|�����r�οj���Ţ_0 ��K7.y,���P[\�'B&n����E?TrFh�.Ў[� ��Of'�^�K�����_��oǄ�����r>��\���[�'��qx(�$���4��y�Y��|5"PzLJ�%��� c�M�9��-����5�&hκ�" ~5���#�U�yY���m����4.�"mI��Ys�����08�}b)	 ؘ��GF�ѰvTy.�r�Xȏ�#�T�!��V=~��CV^Xm�
�En���Jǘ�f='�B?*��3`��xfM~����"sD� 6\�gQ8���S��|HH��y5ڥ��)�	ٜQ���8A���(oDI�Zrm��=eYI�����y��c ��0w$�Z��n��u�ɀ)]p`L,�|��?��?	�ZI~x�pn��Iu�q�ևA8��x�(���k��}���t@��^�&W�x���M�� ����{�u�P&d�[�+?���!=z�A[۝𼾤O���E-���OnR��gi�gi��>�N�����Lご5:  �/6a�AM>��F���u �*aw���Ii�I\(E��xp�eY~1���)m������SE���:�����>����4j֍)��2�`5�� x���8�M8��<��] �	��)�����9��I��-��˪�Hx%�Z�/�⒆2C���B[��� ⺅�K!��rZ��RV`x�@�̛�;��B�m��X���+{��q&��cu�� 4��4ͳ���* �d5I�܋X��/�״�ǔ1S��Ei��6Y�u���.
l�ܥ���-�%ʹϷ N$�؛^2A� ��xvz-pb�\�8`|� �c�X~��J��Z��	 # �� 8b	�cC��8��ɵ9��d�����R�\w����N�����N+��:��=�����#4�mJ�&�6 �Η�pHG���=ט�� ���E�Fo  V��L�oDC��̸>�U~gӺ��@�am�b:XBm(���b���[I�?�g�}�5�P; Y��ݻK;�;txtȃ��i0�{���3��pf8�8�/K�I4���=���w��?(h��5p �A�0����X� w �@{7�7�\��c��S�$zp� X@��79�q�$� #��e�}|��	�P7u��c5GXY	�%���L�Q�����Il�r�n{Z�@�������v}m�'�譛�FJJ b�-8�v_e���wsiԥ�1�Q����z��Mq��
�j놊�.�6�D3����v�L��X�ύ.b�M� �����Z#$����G;�cK�'%[y�_g���[c���z�v96��<���Ǩu|K�tK��nb���7���,.c���p���cXJQUg^_5�k+@�t@P���ea��1��+���q��`"�Ǩ��½p��g�I�4��ɻ햲=h��[�M����Hb�A\}���(*���?��������}]2�f�I�5�:�=%���w���Vo� � ����w��oƙ�ѹ���&d6�!�h0x(�.�����
N����5�()�� �<'�QZ.q�����C�L����>�^����MBF:N��d{k�1�mnv9�Ù�K1�d/��l��I����w�iɮ�$[�|�8j�P�k��[[2��3�	�&����"S�~+�y��}��tݿ��_@{�Z�p�硚����Sm��_}�r�h{\;C�Z���$�����uF#�^��Ț�$ad [�[�l��.�?ΫR	��U��́�ujNOh���iɖޝ�=�w�� �L�;��vr���]�� q�m��|��p�zC�.��٠�#�M�0#q/P��c�;�u䙰����L�jj��ļκ�U�@kJ�&+�2�Y�Ev�s��W-��s7nr��q��J�K��E�'P�6�.�T��ςP����V8"�j��l� �v���&�� 1 �<�*I,������W��mk��f�K��s�؋%X�u䦼1}NX���KXڹ�@Yqs ��*/���8��q���T2e��~vxA]����0���E$sN�զpJ�N��uC p�Z�	��8!.w��H�q�9�(2�l&*ڐt4FV䂆��%2�����}�cK�`;����<~�``p�'kV�`a������	[0&Řc�������ѣO�K����ho�=o�A�g���+M��&���qO�����'�)}?xlc�T�`;��{��1����Xp�擸��{@e�{�jb?�2�Rw~.ՙ��7t�U�C���Tߗ�i�/���J�j��׻�Z�1�jSPf��H,����������Q4/ې��n,EYL^�*�l��d�q�W&��n�'��x�G���x�1mnthˁ�ݝ-�{g�ܿ�%�c$l	r�?�u�x�}x֞:�{��A�hh������Ջ���Y��a��7/�-�����ܒPhM5�)pM]����,��@�r �N�~��p���}fyI鶧�5y&��.����M.�m�!eZt�E��6�ʬkL�Qp�t�D2e��``��k��a+e�wV�����'��']j�+@   D[]�9����<�u  ���>}�����*�1^������ip�k����gC�� n\+u��wm�Y@Y�}��5�lø�ݻ@�\
$�e�����넷������d��T!�&���V��e^2�7�w��[<9��= N�w�� �|�\E;�4nwy㚐�4��m���hs�=\���
:<�����1hԍ6�h2V�R��ֶ%�H�;/���D����3��D8r��ի�a�ֶܽ����P��ǔ���3G܃�BX[2���Ӂ߸�5��C�4�m������T=����Hi���ƾ[<���t��g�Rb�E=�1���X��>S�-��ݟ�aT��:�cM[�]���ҫ���?�0-+��a�L����
�,<B���1%-�u=�dMӜ眻�g�1%����A0�Ɨ�4x�o�V���3f�@gA�{��/����񳜶�z�� �]���o�2�b^i�Ll�oWY�7,"�m0��ۣ}:=#�=���M��v�������W���=�Kf�+�����yyjr[�\�9�Y@c�y)�ՠw�w�e�д=�y��終�]�	H/��mC�X5�f!6M������)���z�D%�i���(;��W6�2C��*-x՞p�9ݯ�I�p�H�<yH�Utٵ/�
��/dP\����r]�U��h�uILXd��\K �љ���*����s}�3[ԝl.`�^���:yV����j����������3���Ӧ{h�T���Պ�4��y0µ���֏1��A>Y��v�>��!=��I�H �-�l���m8F�1�}��F�W\�rD�uhR�����5��$"��D�-<�`0.,b��~����_��|��7t68���7o��w�}���}���7��z��ik�.��a�Ha�����0N<���/���^��^��ӳ3��������v�mE	�6��DJ�\�Ui(S��	�y`e&_�Dʑ�ڔ�]D`k�
*�~�[E{�}�e�,�-gP�3��|n��٪�M ؓ��<����1;�oT�8����
���7�Wr��F��zq̳^����mI�\6��6��qp��E{1=F�����&�˯AG�lP�3�xs�����g�W�Q���4�qBK�p�2lc��}����t߶z��Gؖ�����}��/�:��3����BO��r�j�9F�S.�Ib�d��W�E��M����k.e�u�606{~6����Y��w�y$�O�`�Y�!}N
lfY@�S����4%ù(��dmE���L"4�����J����x�0R��3�x/����P���u�b�z� �0�� Q�zR"I NZ#u%�l � ْ��յX+�M�����>Cӽe��v ��0,ψ;�g�g���X��:b�n��_�,@��g�ai?xi�3�{~����MX��巊�h���ȭ�o���fS��s�~i��Ԃ<K��'m�� �@�� ��ͭ�9�w����v��5�N6��|�$::��>G'�y�h����p����bIb1����b.`Fp#�ɂE�"�A��k����7��>{�������x��>���tz�l�r �������)=y�����w��9��Ӂ�c�X+��I�v<y�Y?	C�1k�%��_�hM��g�&W���x�����g[��6@훅e��$=��7�[W���S�����q�2�1V]D���L�|8'�~ө�!�j��49�|�_�,�m�w�����zn��5�PDnn�7hgc�M�3�̙��S7!h��p���.�̸�.�S.��f���C{ p�J����o��69�,���L�q<���HC/_�kMH#��L��rA}ԍ����T(iR�ůI�Y��m׺Lj��utJ-"M}��.���60�"ٖ�)�Qb�k,�kʖd>.2���aI��Ƥ�����V��=`��Ŀ�ݺia�B�,,�����q� ��Bִ.�(�:��8r*�'��V��'T�dV��&��tde�)�,6I��눋r�2L߯i�K[��?��!�����1ں}i6i;^6]G+-�%~��9�Z�徚Z-����;� ���/�ᚧ]ԫ���e+DǠ�؍��ϼU���	��26S���hdIÈ(0]d�ca�}�J\8�Ȥ���wh��	�38{)j�N�\������#ǐN�uâ>fI����'2E?w���?�w�?��/^�`8a��D�&$e1�@���$K��P�3���8â���6���F��L�����L���Z�SI�\=&�U_�F�+ �Ґ�!���p�¾z�vK#�C���E4�U��;HHC�(�4��쵃�g��-��P��h:~n"�@i;T�m<qG�J�Y�k	���&X���Tǧs�h���G����p�k��������}A{���?��];��yR���$��[�.4OX�% i�H����j.����|V�ڋ�Y`T� A�:߽����-� �th��<�1�}���H�������U2�z�9�8��c�I", R�	� C꺨r�,�Xb%TW��}��_�:�R�M�/2��L~�!�ưHchH�5ZJ@�8j����wڢ(�n\}�}�k�<+��M$Z�s�u�&��n)� <E���!��?��v섯��~K!S1K~��ٽ�l���8�_Sr|�e��]�+�E�/E�T���`�H���`��E{��ɘ��NN㑏� 7MJ��ފ[���nY(��H�u�5���
���ck	m< ��l�_#"1h��x�k�|���T�&�<o�5����ԭ��	_i
3*{w�Z�ż�!�3�Ǆ_�4U"!}��3�)\�}SHwy@��\W��V�����m9"[ �����W*�-�9dM���tt\�� <�9QV����zݒ]�;��-�(���dn�W:~X8�;��~ϻD��}����7Np;>AB���O� #����~��iZ�
�(]D�zQ 8ςz�w^��M��zu���DI�Z �E��E��y 8�"�Y�fQ��/���N��t!�%(�����������ldG��a,.zPk���J�!X~a�E�#�Bm�M۶��j���F[�>�Ulx^�R�W\�e�W�n3��a�xf)�$q����{UF�ykk�:��(P�Y ���وQ��2�����Y���[j���J���N��@�1 ��y��yP���[��J4wؠe�bF�M�p�SY��Z����<�dE���Mα(Y'c���Xbd+L|��]7�1�wY�h�a���U�K�^Ʋ_,�MK|���b4��"����:��؊]�c��I~���V)}K�v�\/�7�v|��9���Q2M7�\c�濣\V~�x��9��ŮqK�$\�o��+AG{3dA�#�E!鄎��9�'��!f���6�X:9��'���7t�z�V`�"�;���ӧ�w6o���;]��2\�:�X��v�n�b)��
�,!˪ɷiw{�>x����Cz��	F�.g��r���ܘ��-��y(��&I�$yH�ۀ$�<�3Þ�ݪ�M����I���/�XkԾg'�m���IXfa����-�-���2*n��B.dU B#� ��sa�q�9"�%Xg�!?�x���v�Mh#涶����!�"��m���� �}�+ĕ{U��Y ����ޝ�W��Y��>&��*I/�M�[�u�ŨR  e8n�-��jg81���ך}s�`A���okn6Xh⪂E�0�X�bp�o��
�4 ���f�{�S�,��\�x���Vh2/�f��.������F��$`V��&dc�k�FA��gվ�[�Y�&4����`�'-v��8;���f���U ���WA�,�u�~r�0�d`m��7i8VNv�׿%M���xjVވ��M�Ąa�q٭���w(�&�ǜ�����#���!=��5�90�e ���=:<>��<q�m�(t�6~��l��53��	��=ߤ��.=��;���a��xZx	���4��<����E�ggѢ�tV��&��l�� _���s�i%[�ڼ��V�Y�d]�>�,�weȓR; Q2)/"?�' ������nψ5�u%��M�N�k��&i�l��
YZ����4��w��do�^X�aEǽ�L��lR8��Q�k��Xd\�YS/��k-�U@7�l{H�k��Ҁ����'��M"�	�M�@2��`�{��S��i*ж�y/LFkʰ��
��#1ȕm�5�o8��5]�����x���rx^XT��>����j��}������P�|]�4w����u��(~j�}�8�E)�g��5m`�ģ;P�5����2o#��ƋU���н��@�|��һJmnb����!��k��|��X�T�ˤyC�C��������c:x;��ߕ�<��Ё�3��Ft�N��wwh 8�\��͔��b���~c7W��FC��}�7�q������Yy�bV�[�Y4�,*]d�#6nvL�Rz�Xrۮ%;�Q
�Ēw�}m���� �PW Խ�<��DH)E����B�D����x���1w zq�$g����W\���9-�u�L U<�$�B�qｐ�s][|u\Q�@�����
�_<�$�Ze]쫤U(�4n��l�ŋ�ӆ�z��c7 ���j�ۆ��&��2 6"[`2�e�&8H9�OƂ`�`H��2�󠹪�w��0X�M4Z ���ǋnXh�0���E�N�{&䀰�pF�E���w�ޣ͍M�j9��B���Oa��v������чQ���X8��s�%���ژ�m��0ܩ}��
0���D��^МQ,7R��+�ؾH۵�mW3�k���W�'��o�0�[�h�:h~c�r�n�r񖐖GomU<���5��$	��e:��T�67�� ���\��� ��
5��N��ئT���'[i��v_D�l�!�%��i<�u�9b߾A�h�z��#d�/
X�'49����S�w�K;���,Dy���5�ц�<h˄s9B�id����c��gDU�c薮�V	 V~�؋�m�����B��{��+���L�@�xQ�rQt���"��>i��>;�����&YudMY���;D����7�BCn|��ǳ�j;K��} �Mٞq=�@) �ɭ�2I�
�"�1,�b	���/1�m��m ` a ~��ծ��x��i�ʃt�m:����x�e̕���Yt� 0����2Sq��wYw��,;~���Ā�u� �:����I��y��$�.Z%r
@�#C�1�F�=��,�����փ���/���?�(���p����[��@"����^�x�و�(���G0?p�ߣ� ��чn��P��`��np��������������Ξcno��d@/�?���/��>+�xx��<̽�uN&����@�eLr�c�`mh.�O�dಝ#�X&�u�t���Q�K�������οF�r6��L�j�������>�5�n>B~�QA��6&� dᕐ��8���ׄ� ʭl�[�/h�szi�ןٽVΟp�u��+�k�v�j.��0������k���M5O�Z�������n��쐛_�	���BG~�g>�I��n�OJ �[�k0o}!��7o��ͮ���w��N�)%F�z��=^�4t��	F�>��ߡ�-�҆���@V�b�R{��Z��M��f����e��<�*\������[,w�)�����Y��U�&���M}3��ۨ�n�xm9��2FJ��-�$)է?F[�.=� � {�}�� 0(��:T:^8�S���� � ���w�wJ�!�q^Tyr�5��/�����O���D��\�x[J�<'�/2M�/�Q��i������S鸟�^���i=�6�֪�sQ^�n���0 l����(�-`Y꘎��b�r_�(��ǲ�붜�9y��Y~�(���/Q%Z�n�5827-,NSρ���m�Z����"�����,	���~���������{ߧ�-vy~����glY��ꋘ_d� �Vo0rb�}@�?��S�dz��9�b�-��,1���>pd��=&%(�߭r=�~��+�΄���K���4�Z�7�~y4�>M�,�JhVb�K�V�u�� �|�/��* áepU*ˤKL�
Y�}m���q��y=��%��}�<���_���q>م/j�	\�FW똢�J��TY�+ \x�+��V�2N��,�T�H�j�\f%�[��lˊ�jW|c���.����$�Y��o!��ҥ�:��+�Y�%��V)�6�e��f[�:)-0睷�B���ۂ_g?�_#�c~S�S58�f>�rPS�e:��Sb�O���Sbd�����Y��eQ�1���޹�ےiG:V�� ��"q�h�W�ɖ\w�Ƕ�ٵE��m�� ���i��ӉhA�a��m[ɘ7�:-�|R*K�R��U�MQ����stQ�ps ���+�;A�)�JU �lH������4��t��OY����{t�ތ��
::�sKOث������v���vQ�eV[,F0���cD��"D#s������Baac��B|��]����6=�����NO�iwo��< `L �/P;q��h8rm�>�����@w�G�_p(�*�?SL��;l�-#O����e)p`6�Do�����g��:dcX��EІ��\m�ߘ�r�$����R��础Q�iE�{2�� X�-��2��͏3��pI>������iCx�����kN=g�RM~R؀L����)��C2�ۂ'��C9�@˥Obh���m��ݲ��x�f��$��U�J���.o����|zr�AD��� G�-(���	i��^ZV�Z�jp]�ͭ�泶�4�<o�6�Ϛ���l�E-���~��'���ӧ� ��|�'�/r��7|�Ě���'�O�mV��"��.Kϟ?gk�X�lE6��/�fCFX��̡����&пN�ĺb�%�-Tb�sJ_����2GfY�uK>/�'{�� �b] F�.�҃���t ��7C֏6 �l�� X4np�s�n4&~'n��q<Z	k��ո�	B`��N���$�?cl�}8�6��vrrJ?��=}���л���@����<���`�EvT��lm���=���~�/���.�e��Kr��[d����޽T|�u�m�~� 6ܚ-gk��4�1�Wl/b�1Q��#A�[�})��!{� �Џ��xbKO����6գ]h
p;.��4h��UB��v���!�^�unud��`5󻣡Դ6H�7�	++Jn�W%���>&?��Dt�q[�.b���������F��Qk>x
��3��_ѕ�U�[k�嘝�ݎ^���:4B�b�������t������&�n�Y)�K���oR��
9�.#�wRftxt�
ΣK����A��~����	Z��ⲴN�E�e\�W!l6Y�g��<�iwL�Kn�L�tJ�N���}s޹.dI �ԉUV;$DE(�(3�
 � �����E5Uzh�qU���tL0�
Џ熜�O����7��� �p� ��-��{�Rh�I�f�wBնԳL���B5�SϺ�U)H���`S	� v��.q~�{6���+h�FU`򥒴-�]w ��N�
��48C\�c
[����,w����*A16v�!l4��ֽuw�'>�<k~�6��~�� v�h����b!h48�÷/���� �B�#X�����[�ۮU�4;F��Z;p�܁��ދ��u���>#�.�>S6 s�o�D$ؒ�8 ��r�/���;�O0Ɩ[׿��}�b�
�E�T���EIƓǒ(�g���#3PI�"2�׎h狟� ���;&�^�nHM���d=7$�u��N:)'!�;ɸLt)��M�b,B��2Yv	�aqg�[Z�b�p���3�hsϳ^��CP����
R/��=�!	Tɬ�9퓶��L�5���m��;�q|m�e���t�-{�}z�ߧ�w6ho�� ���5��ڗl+�k���U�u���k���S�Yz{H�ϟ�kD'��Z�W/���-��R+K���c��hQ��E��K�W7��S+�E ���|���(�q�8����a%޻0�G�O Hq�����I����`<,� ���%ɗxH�"I,�xVX��爅�2�{)�t%d�?�����0O��\�pSp�-��lM%���:_{ \뮠y �##	`ѵtx<��Ċ���%�7�[��ə��;�{.�"��O�
�B��]�� j�����LX���gAR���=:9>���*����/pe1�m��������Νm��Ga `���m)�(m�r �t��.m���u:3�/����/o�s�(��c���lq�rm�n���Ϝ傥RQ�:��W"�ݩ���elK�1�հ^"M oT`��P%�<!1�� ��	�u&^C6��4r�W�z(�2ԉ�;���~�P:�{�����S��y(���(6�q�"�&�q��q�罨$��N�����!j�!���z��<2~Y��Ǎ��2zp�f𮭮�{�j?.&��d4��v�j�#y�&=��C�;���q x��}R�R���B��ˇ#r���~;����	�q�X��n�<�� ��ZG�ݬ�Gs]���rpMb� ��݋�h���ː7�{���6�G_�~WfX5��UO��q�s$H�r��@f��R"K��)(�N`����x<���(�o a���� z~a�F_@6_W�g�<`}7�e�&�\c��<6A	�f�m�~Y$<d���� �S�T1~5���VA�II7� �_Ƙ1}��˖1Ԇ�Дqr����|�BL�Ů���❏�� l�8�nt��&fH�py�A��??��Ϟ���!�I^�0��v��o�?���h��C�ۖ;�8����	��d|�:�s�	���m����#���VXt�*��_�>F�����lQ��G���F�ޘ�y3�A�M�`1,6 ��7�7��y�:} �>�F[[9����Ւ�E��@ຓ�`�+����~�Z��\�PǍk�rdޝ�+�(�`����W��Ľ���M�;r�e�(�C�һI�D�)�+�1�:��$�5|R<��,6 ]�X�9�+n�䎿��t��ߤ��۶�����;�:��ۢ���:�����f�-½��t2	1�� �փ��_C�mr6ГgtxX�]�{��-����-�� ���MȜ�� �Zk�M�3�͠�h0w�{,#�_f|��O�4A }��9BXBa~������ɘ�қ�\\S�,w�E�����K3��M��p�~��%�y��z������ů���:�P���-h��b��<��y�ݶg��}����� `�,���(���w��1�{4d�'L��p�r��`޵�gC."Ε07����~j���	��� ]1��wc�G���q��%[����l��?z���~���l0 .���&(c"d�u�sk�cfX���Y8�;a ʱ�l9�p��3TU�EN.6��������l�z2Y�A��1��4�T&���cȮm��	��~~��	�C��pҭ�anX<�s�2-�L�1�~{�sʠ�%�����MCtr2�/N��i8S1>q�kH��Uq{�ٹ�}���`�r��Θ��T����c�&���w徥�"5�mþ��&�5�oe���Ҡ����\��I�b	��s8d�.u��ק���mz��Ր� yPvr�^��l�{�H�fB��F����v���9�9���4紽�!�oc�V�--GM�W�|]_V�&Co]��"}1 JV�E(�+��E���OFC�`�Uu���k���m�I{�	�r�� ��]&qN۾Y��y}�H\u����&��"�^��d%�k���O.u����c=�V`���]��\_�|���lJ�1�W{�Gݮ7*IE�C'W��;�]!N����I���[��ѬqiZQ���O>N�`��dXB�9����IS�y�y p%�3H-� ��8h\��[+ 9���l�$%_��>3n��yΐX�b������X����k ��r��O�Ԡ��68��a����6*<0]XwaI��	_��zNH��͘�7�  x�?A��4etd�Ў8ĻK��r�����3>a*�C`)>88���������sݕK��J����҄�4F���lw9��xH??}�>kL�S�kZ�[
�o�n5�`�[z�e���UB])G�ş����쬠'O߸1E����r�8�Ag��j�/���0,!�� �♼�1��o���q��<���n!��Qͭ��lY����.��Y� ��dw�II����q�Ke�5`�m�kR㖥�q@�S?�}'�l�l҃w���è�0�N^P'+o/���4w%G�Xy��W�����l���S��W�髯�з�=uB�}��$�J�2w���:WM��N�M���a<<�:�E@�"V�e�]���+�k�ߥ�u;�y�B;lN�D.��8�-sD+Q�2�:��ދ �Y
���� �	)e���y�Ӡ���_~�%[|���?2F�Ux#"����?�c��9Uj�����.m�dQ�xU�$��AVh���������ǤW:��,���_���E<&���ʒEp�iR�Քv*��M��� ��
В�At�
Ԇ�=l�@l�FDn��#[=����� �Y1`:� ��M���#��x���`x�b S����{hّ�� �܏B��o@ەqi#?A�,�12���>��` ���ak��q<��."_m��������^��V��F , ]�u�̬����xR�`8���3M
�_��Tڴ�Z��^J��j)�l��ʊ*�������pp��}LG ��pQq;9�Pu�����6��pƊ�(DNܜ;:>����-�>� �%��f%� _RJ$(�J�qv��SK�S��.u;p��1�w�����޾�]��
�r ���0c&���������s4�X�w���?���#}���~{D��A��#_�PӔ���Cb��A5\�I�]��m�)��w�,�<� ���u��E��M ]ߦ��E�)���;�&pK�n�ҵ�
���M�˝�6��_��G��$~B��@ ��(}��5,�+l�J_kpu�T�f�g��VN�{^�I���/J#-�u��]��K�|��vV��"�&��r����2L����7 {�4�5kc�r͓ߧ�����]|�c�-r�d7M<�/aݳּ�@qo�P�������'���O���9m8���g �8������ctܢ7'kI��K�;w����!Mə�J�舳m���m���� �Gq8Z�(%|#}���e���}�e'4�g�6��\�K��ɬ��&�)�\Β=�Է0�s V'�##�� +�^�ުϞ[&���j�Hq� �;��j@���͕��(*�����JI+���xE	�qQR�ɳC:9zK{�=����,�YI�"wshH@��z��1�yhT�J�ș���Ƈ� ��h�:�'O^�w�?��?��zK�'C���t�|o��b�~L���=7������!\���7��CdXE.�o]�����6Y�I5X�~��_r����z�ڢڕ����/���b�5p�20Yh���5O�L�#�J�qU4kL0/~���r�?��l}��1g~������D��n��g��eD�eΈK7<�~�u�����_����_Q�]���F�vL:?����MAfM9Eͯ�u+�v,B� �by+�D�GU�Iӄ���0�|��k���ba�� ~��r4����1�E�"�O�-�c ����7���k<A�+˾��QəT3�a{f
.�ı;�wk	h �;���l�R~�b2�G��Kñ��=O�9٨�o9[�بk�]�\d®�b[����բ�7A�r~����ڂ��8�q��=�=7���*��L�j��x��Y��	๵��MP2U%AZL����N������ų� ��dV�;}�{��)�)�0�y=�WIpR/������''#z��-���}�������������m�{�k���#ņ�l�o��r�P:a�K�d��
kp�}Sh] x�cf���Ƌ��9��W���wzv�ݣM*�P��o�L-HM�%oik������?e�`�5J���F���EܾS���}��쮊�>v1? 
A/^�`E	ܢ��p��Lк��,��IM�	2ޢ@A�/�V��y�7�_d{�k�̷��}�)}�t=/���9�n���em�pSC������= f7� R�V�HE���&Z))Jo�%�HZ�*�f�e#0.������.[`�6��a0��Q
�N�������C��٢?���}BR�L�$Y.��fg���[�:�����'4{g�#���!�Lq�L��2��d�IĞ+�`�Bk0\)!�~�w��DLWC���\�Ҷ���\��
����7�k�};�0�Pj����U2��	������F4�E�*i��j3��:���L"������������!%p���L��C�_�_���0�P,���ȟ#�)���NN�rvvLg��z(���y����-e�|�����K8Y{;�%$������߳5	581F�QU �E��,jǃv��ϋ�k���/Q��񊢜�O���'��g�jX�Y]IoR�j���$�5#]'x��u�Y�z�jj�5nr'mk��:�rzL|N[?O�c$e� r��_3�ꫯ�D6$ʂu�wwv��؉e�d�_��[���x��*)<�Jd�Fۥ&0,� �O��*M�话�bٽ5]�>i����`���$ x��UKj$���H�"�([Y��|k���ZA�2<+Ҧ-��m���nA�b\�������ƨle{��+�<���n�	�#�-'��H�����x��Į�����	�[[=��ܡ>�^��-6��*S9A�� ��6
9a}��n�Z�H��j���*�[L�V-�U,�ȨiEd��O+�l���coo�K_����a���,S��������3?iy�K�Dn���&|%��6��||n]j��wgÂ^�:�~zIcǳ xʑ�~nz�jP����c�:���j�f\���s��/�����.o=���� �c�Ÿ`��}�x��^�R����2+\!tB���� q�\ ^�����T������~_����Ì�%�tpF�����|�����o��}�v0V�R;�eW��g���6C�Nݬ5к.�
+�O�Ch�'<8`hA��� o�78,N�1\�gI��b�E����+�I����Hv�/ܞ�A��Ƞ�S"��?>Q�̲��؅��H<9j�&k����@���`VAߪ�SZ\-�Ձ���4
�@�:I�gQ�CKb-�?um �6Z��o�/?�%H ݗ�^8�z���.d^e �~�x��S�h�E]d���up\�X`y��?�wO�yvT2����Ѓ����G���;���@ʉ�p��z�'�)�fwH/�z�K�!��g/������h���=C��2@���ǭ��+���a�d.r�i�v0������g����~��]����k�n!��[���$e5��qOq,7אkRҫWo�ۿ=}��n�]%�C��=�Ƶb��[�7��EF�g%&���9�>S�Z��R��8cvk(Ɩ�Q������o��y֥��M���\Xx�--K��Z��c��
,0"X꘱��v����e
�u��i�3�ZcV�Y��J66	�M\2�'F7Zi�H���㤭�MB�n_[������9���=_�5�I��%d����xS�g1��.J���	C.�e����>}���X��K4��w�����N���J�(���r|g0dO)
 C�ǟ|��� |��
��ŝX�S�ɕ�����)A��P¬u��c�:��ۼp��P�G7 �_ ��4'��L�43��3�&H~�&��������"�z᫩^l��\?��Y��̂��d��G����*�S�d�F,�	)h'�a���˱�b�wT��sZw��-�m�j�mѯ>{�~��{��ݣn� ��J�L ��GDe�-��N����Y�I/^�!`D��'4Md�vǨw�Q�m�[z��[ӕ$P���9*J�u��jy��o<�K�?7��{���G�����ݻ����&X��zV�>9���f9�A�N�&�����g/����d8�f��kL��@kk��j�Xc�wP���[> �`䄓���MI���U��t˭�-QI����X�'��Tׄb[6l��.��{�ߺ���똺�
�P+�>Ǉ�$5�#(��O�M���cy+��Y(��eߖ���z�e�y���T~��cb?��;�z��|b���^}���:��<g0 n�]����g?׬�pm�I��� `M�6�ߪs�,�r^�`�P����k1жr	��b���{f�%��zż�����.1���b#v�O�,�qM]�Mó5Ygy �c���:F�h;��'�l�����{��=����+n�xQ�iwg�2UɶYt�A]
������7>��1Sה�oS�\�>j���5�Q,�0�^�-f��W1lP&����l[�������ד��ue��4=eFT�!�&Hp���z��bP���:O��Eh�s�2`q(j
�ntL�
hi�%���Y\?��C��/?��{=�w`a<q@jD�Ղ���-� x���e��e�-�غG?<yCo���[���������@���¯.�%H��_AED�����5C\�-͹u<~��w����N���; ����/>����u�>psaH�2C"�X��֭��FI
5�7(�n90c�x�b��s�+��V�̇�?��
{V�w�������Ǩ��eN�.�㺑�V''����TP�X_���C))����%�F�I�`��a���	m�Uo���]��-�\1x4>s@��ˀY;���a
��R�|Y�Zj���)%ܸ��#�Zu](h�e^�x�IF�7%W-(��+���S̺=�J�
b�F>�#s8��"
_2�g�����YR��!Q�~�^Z>�g��s�����Ia��V��YYa��I�zD�.���2�2ښP	������H6�P�/r�~[�z���V�����c�1S �*จ����E�#�4Hj|��Œd�j�"�]H�"bp��O0 #&�`��"6�`˨'P��{S2�6@��US��~b �֒�5�'6�ed�}�������ލ��V�{�k꾐6��7��<�Ux��<G
)�R3�i�o�  ����d6N�J��L�L?�P�ش�$�� ^��z��Q�,��&�Vx��rJ]d�!&�4�fQ�f�[�$�S|��dW����ޝ�����iL�5�����J	���֙��fga8[u�.���Ag�-��٠��DXZӱ��t\Ш��!T�5u%��본R'lu��}��d�:��8�w�����҃�>�w׽���	N7�0�2�
��!N̋�ˇp+͝�y:���es��k�e�-sbV'�L&���V�Dkp �60%o��Q�XS�Xm(G��
��z��9W�ѥ}�(�S*pސ�e��;q�T���@�PwxR�8���A��������%MmZ�4i�y��f�Ž�;��SPb�l�y�'��p(r�!�>^��q��q�o(g���YPfg����U�[@K[<[�j�dʵ�z�+E0�T`(��L�*�+[�?����j�Go�/��M�O�1���k*��36��閾�g�G����Y�I�㢊��v���U�_�ʻȹ��%�O Zl(e���s�t8K4x�Y�&Љ߱u8?������Qkc�n��2j��}��=Xs%�@.�+nܨ�0�I�1m���B�1���B/���0I���q�4P�It� ���y0Ǔ��1�H�Q����6
�c��o�1�D������p>�D+�:��@,�5���7���F�d.w�MU�[j��v��>�_|f����g�slϳ{�-�[�R���{.Lb� @I2��͛W+�2I$�@�b�;4l%IVf8,e�!�tu�����uP�Ҝ8�@Z� kG�`6������a�^����0�|2�0��E]���< ��s/0��YN��[yd�^��䟛'����!e�_���3�\Q�������IZ�(i$Rf!��Sj�;t}5���D�������Ҝf�w���ϖ)�z��f���)S) B�oKtLP�m�L�c�G�r��j�3�Dk�tk7k����s7��q�M,�y��*b�P�%Y_KS+@kb�`�\��a;*�'HK���3h�N,͈W�x��.}h��&�l���3�3����xR$�$�����ʽu�Yk?$X�OѦ�Nb�;L2͡QY�=!9&͢$
����<xU�o��h�wq���*�KŖ����}�"�_���:�k�}���3�UW��9���L���k*b�aF|0�a}���6�0�(6X^���,��5��	�V[�b�w� � ��[��/��q���R�l�D���8W��p�|o��������0��f�;,O[��h���L�g��|�V�~�Pl���^��ϵ�b��2�q��Ρ!����3Sҁ�5��Fpf �x�L���$R�2� l^k.,���G�+�P�2�O�r\p>�d7D��t�gB�@垧�ϵz*�V�u�}��0\:o�w��012'낪�1��1�m��e�[K����'�x$a ̂��fv{ד��@��n�ty��{")��i���͈iU��̋�up)=:�����I�� �s��r�D��ziJ����2C�&y
��q4�]���;���4���ݩ��7�(5�%6�SV#"o�`˳��;T;&B����Dj!�Y�B@�a�0�.��8���0s���S���V���pP���G�<'�s�)1����&yكCV8U�iu{���j�����l��*%F�_� �:��� 8T��Y��s��2*�V_�Y����� ɦ`�@���]�3 �$���	�o������B�|=��b |����P�	V_���-�ϺO��m�E�_z۶�����	R��i��M�u �&� ��WTvѠ|i4I�&��۝�#U?���Ą��� <���I�P�ץn��sĆ�c
z]��$�N[�Y�s�E6�J�	���`�N7ak3�┬f.6�R/�U���H"���ۢM�2���u���0
��Kċ�X(N;�8���b/M>��`�i�l��ځ����M{ Z%�*gA��Y��J(�lV�����`pm�Á:]�ȖOJ��w�LS�@C@
㌑a�������1�슕�|^R$.�Ѫ�`l,�q�_|G��g(e�E�y}�k�(I�5�B�X@LhU+�ܯXCB����Oh�`Ϭ�vU�<�$3 97�0�p�և�ت
�w��FV �l���	/�.�Yb�AA�B����-ʀ�f	ϛpgYg�W��z�/��b��J��+���k
x������_rR)���hl ���x����H�!���&l�%@@_�gc��`X �d�_&��m ��/r^ ��T	��u�MT�Gw�� �K�m��
Y���7�ثu�]#��X~���e�D����t�aF�J�}Q{�N3�,d�z*�xe�p�xedK@�E%e��X�s߲1N������ o�t���}J-�O]3{�KSO5T���d\��f�D��;�ڍ�+�DFҠ�Hy���u��m�<+�n�s�Wl�?77��c'A��C�������x|�B����7�[6.I�:��+/e��Ѫ��[���h�}��?�,����z�V!�e�)�)��HS�� ���*��o����Ҁ�+N%
@-�N���,�;�<S���y�H(H���*����u�޽c�rL��~�C*7sT#%���v�wۖX~s.#Q[����^�zG��fψ�S^j�) �y�_�����z$�����1|ƫPP�G�[�Zn�����Y�7�a��샼)��X\� ��4@�X�%>7,I%�J"�;���;+4�/ 8���ko8���l#-3��\��c����G�x�KJ�;��ſ(���P���HVBi��\���0���W�}�e�[�Z���L&�c9�N/���7\Vi���F�8��3H�8a_��sa"�LX ��:r�@p�\����R�5�j��jĿ�l���-���*N6��8*O�uNi�o�.>��&l6OM�qv��V��=�vt�)�*С�\u�-M�%K�n ����tĖ ��8�����ryq�5�R��ƪ�mı�;�Y߿w�!���5��W�����x��ym=�:�$J9+h�b]R4\�~s$����g������n��CPi�{����a(˺��X���h����<zH�����������/�va�S�SCMX�$�.ْb9u�wkm�q��{��ŋw�?���G�~��Y���*����s���\5[Ū�:�Ⱥ,�M@����Ն*]�+W��w�(@��D ]7��$B�mVD����g�&x.,���`���s��Ŋ��_�b�/ڕ�\�lKj�b���Sa[B�����D[ <��U�g��v� �j *�Ql� �Hx�n���+g�X4�%O���u����5Y�1�]/d>x��(;sE�g�v���������Wt��	p�
���%����>�>  �=��9f���,0� ��`��s�-��&ɚ8F�.���Ӕg>����%T��xs�j�W��>���j��3��q��V�<�����^��i%ֲ��B�Z�����V����Ǻt�T�'��VP;B��4���B�Ds����]���TK3���fؿ�\��ʡ"�k���f�0;�XX~�߻ǂRX��`߀�#.���$Nȷw4/���²�po�G�~�����>��><6�ɡ.�e\�י䮜�W�j�=5,(��׀A�����џ��-uvlg�i����A�p<����unK:x�Ckܯ���f~�чO��	}��N)�1 �������
���3uQ�� ܾ��3;|L�G��o��g?v�66(�Xr��s�������^��6}��۸K�����o�;g�{xn��
�F�=�c�^Zwϡ�w��e)�D�n�`A�� �H�r��x� �}]�E�"%� ��n��xS]�=0�yl�ռҢ�ƪ�� ��� �<.�U���wU�ζ����&� ���TU>��)@�p��0{ZE��^�K��!p�	}��/X{V�LYf�|uyI?��#o�~�l������׿�{�o��7F�ۣϟ�hxA{.W++'�P.�gwV\�֎@¾a*}�w�#�|�^F#���!'�h5k��9"�R�G.됒T��[��Ė��X�&��y�\?M�(��m�I�vs+*Yؗ��L Y	���b��?����O-�p�+�'�p��GC��LHY ����V��6��:S1CHi����X�F?�寠����8^]��h�y�J��i����kU�x��4z�`�����K��-ڂc�����aX%�"��!b�X����0+(��
�$�ɯ�=؛�^+ԕ�^�'��b��[Cs~�Q'AN
g��-�!-�E^`A�s����X!�����|�3�����P���YK/������GfU�*w@ݺ>[p���'��!���Mf8��u�V�����?*@�<(Cݮ�h�����vBt]�XH��QS,cqǜ5�!�X�ڸ�����G��l�N�VgE��fX�y ��C��zS��:��:�0˰8W;�OI	K�ͦ���
=������m�Vϯ{����i����(k(�uP�x*[bm�4k�8b+F�,l���i���{�wyyE/_��^�O�=�OP���c�{�&�K�F]:9�������9/�c [,��=� e�d�\�N�_�5� �&�yG�M|"�.ӈ	��Sg�M�>lh]bܖr�_��*��m��7˄)��Q�UտX���E����������^�����ɵ�@�n�j�KD3οU)�j�����N� ���߹�h��� Z��p���
*��9[y�\{��w���;�����_�lGn��(�K�Ֆ�U1(	���GY<��I�=�n
�1eɥi䚔���uq}]y{�� <�5��rNT�tq�#��%PA���K΅����"q�$�Qg��w���	]�c�:� >c ������/��9�JI�3����Uv�Z�(/�#���K�T��*^�"�ͬw���s��m�cӵ�΍�S��Uu�"�ʊ.�.�@q��4��;e�k���!�|��ZW�8AXS?������'A�ƛ�P��}����|�}��q�s 84�W�Z1	d81��?�B^E�#�ly��_9������9��^b[r���^��S��8+����'=��b4�Zs��)̔z�}����bD��חX_����KVP<[�1A��n�s�r1)V@'q1��W"���hM��b��Ǽ�UP㚩�O�]�t�ڕ��3��EX��h�a�b����V�W/_1D}�O>��>|D���v��M;�adaٯ(�g�/`�pJS�[9��ܤ���A^e�Y �\� �+ G���P݄C|����wC^�Sue�0��_��}LlB�!ʺAۊ�"#�9g!������(�T,��KM�=���/h�9B�Ë�L�i! ܰ�NH��lS;�Ь�'n���Z� �>q�*���*�;o{w�Bp9^IX��Sj媐���>��<}��m$�-�����68[�UM�\�򑁥3���QSbӐ=O�|�|p?����w�M2��bX`����� e% �Et��RF���-:AR����9ʄ$$�<�۔uS��$��X؊b�"��d��Fb5	h�0!���퓬}���w\l�n�&$
�`nh���㋿���BB�� ��HH����g���u!�e/�7r)��=뢗������2���s�P���*iG�"Ɓ9�i.�7rې-���Ԃ_�H\��Z��yi�m�gP&
�I�o9���PWw:tߕհ��iE; �Y�a��Of��; �_�e�ǺL"��M0�Dν�`鎰q�k���Z�� ���y��^��"�tU�kK��nS�U.��{x+�m�Yۦ��@�]"�!�-%�[��$s��y�qU����u��m������)����X�藲�6�r�~[r��/ܪ�w]� r%9 z=���wkp����āPRl�����~������#��f���t@�� x<� x��S�+��*"����rHf�e% xS�nh�Ф��5}9':����ǡD�~��;��;���TM����ڹ&�����u���X�ӎ~6įt��o�.�<q��vJ5Xbb�� ɭ������$Ί�3��
��o�[�W��_���P���[���o8� xr�-#o/+�+�sf�v}��`f��\U �5�V`s�F����h����_)$��(�HZ�s@ּ�m�¿�(��;q���@6q�H��Kr7hv��>�sǂ~���>�[��(��m�Y�w�c�s�h��m�RB[��(��sGw�D����n.J��J���6� �Yn�U}X��f�2 \v��F�h+ V��	�^�np<�2(,T�`]�KνS�GM����&d�}&=�9�@'֍'m��/���pNb6�b�&��B#��n��nT�Ą3E�y��Irŉ�b�r\��r-`�1�6�IS�?(�D»`Ӵ�2��������|Mȩ��� ��uT��J;$;hYl���"�D���Y>&��0�����-�(`�3݇g`��/�����MbR^<�^������c��"Ǜ1�Q�%J ���FO>|�`���7����J��]�>��Ԫ�"8Tשq����9������hB��s�=�A0s!-��9B��J�))ɖ��_ϱ�8�� 0�=5W.Z;Y����
l7h��W�}ӮU'�(�Y#�\���,��}�����۶P,�7	�U׏�ϲ2N+8槦~0�2|�r�VnU"����?��U��]������P�_E"�0Yج�$�c�S:_��2F[�u��㬉�@���/���V��hb� ��{U���!�:�.��,ic��n.3���j�}�}���"����~��]\^Qm-*��|}���<efu�EX0#x�!-���.��� �d�ᗟ��Ɩ;�E�y+��҄k@6����]U�V�e�򾺅k1���Ɛ��p��Iu7��^����W�L^_�=v�*�`��L9WĤ��A��CA����T�.�|���(��_�����~�;�Y�2�B�f�.��U���O>|̙�����`�E[�,�f���HDhɿ?�w����F�ӟ��O?q΃��K�^K�݌_���	�7��U>w%���l,���9��r�%ڮ���it3y
�P��]�8��� ����deEb���'��u[�\~�KPHm�U�s���
 �
�Ѿ8�v����
~ς���ٙ�Nϡ.�c�k�6jc1��b���FX�����/"� ����Ҳ������-b��" �H\iy!�6è���*�2i�)8w#hN=hv�"k�[5�X9�ǔ����<��*��t��5K2�4����q�+X|��(.Ѱ\����KN��χK%��P�(g��.�eK+�ն�`u8��c����+�e��ּ(k�5q�@w˨�=�eX���(a�.��	2��k���K2����˓��[;�PG"��`f t���Ŭ�zjA��oŽ�����GG����{�*5�y?�$�R_�l�+��d�v�Ӕ���<�g��B��F?u�V�Ϧڻ��9goOF����^A?�@h��h����H ��G�t")cyx��y/,��$+<W��`p��og�r|�P�^6պHCaxf��K#D�`AaKp�� 0��=�e䞛�ݻ���v��x�-H>G[���V.�S�xE5�쇎X_��Y�c�'�
Ϊ��$e��������9k�|���S��y�c��<��ߠ�Du�N��Tʹ`�|�=�m�][�ʸ�: ��F�1u ��ϫ�?�������I��MXC�2s��Ǝ��Hjãc���k��|Tx��D�c����u��>?[������Y���%
�=&�z)uS$��AO�h� 7ː�jBÑ�p�S�; ��ɴ+��.hb��i ����l-Aq����#�=��?��A/�6X�ESē��[� �N�K��ʀ\2�pSFf����u;�/G�l�E�ϠX%�/�VS���}W���@[������M��vͫ�f�c��a�(�����X�5Ş[�Q��Ƽ?I+�/OM��~y=�$�d�����0ُ6n�=�T$��AR>�R�٪Č�ɧ;�9D���A*p3�4 0�)h��ͶJ�yh��('��Ż�[^���A�j�_��SכQ�:=[a���"��Q7�Q���% ,�6��[����4�mI�>�`i���ؚ7�����7������CnL����������<�)���oc�E ���h��Q"�*����ocEq�$F)9Ŋ��Zq�[�!��Ex�qB䪯�ՉU�t�^Ѧ�B���K2Ҏ����ˊ�"Jֽ#�{�W�/�g�ܾ+�*^��;�����{3�r�5 e���j'j��}���=��wO	r
)��&�|O,{_d-Ilj���j���S��V~�� �N�]�VѶ�/K�V��޽{�<�իW,�cF)��Eu��.��~�sμ��&B���FM�n�� ��~����oy.��C޹��Zp,��Y��Y^��č1��3��v^(���o ��I&�qm=dD�wԥ����H�������ܮR3���̤��6���J�����f,+��N@�@�^>��S�CP�&�c��oX��>g�Ƌ��b��P�w4�� S��yl=m<A/5�������X�~x���}�%}�fB���ľg�e'q.,6@�`���M�����y�,6++����q�S�����)7�ۀ���/��4�ź	���B��Aܹ`]:�E��Ͱ�rlu���{���*"��HX��f)
μ�1�<���c�������5[����7�S�1����m����JQ�BW>����o���+0��C�'"K	�&����cIb�^�yC�|�+�l��d�$���U����?���)�^�� ���a���$M }�rP�Ūg[����kM�y7�Nn�����x��{��S�Dq��8U�~�k.���
���t���k����)z��ߓW|���j�_��ၾ)QV%d�<����/��:S��b��� �s����Z��\���)��ceS��3}q��ye�����Y�}4�I�a�%V������$<�R���`q�m��V9������9l���~��^1���Af���B��O�7ϖz�m�m�{}�]���t28���YHa� �{��=~xHǇ��0#B��2 � ߣ��#ҫ7�f�)�_�m�(��H\L�\�BX\������Ç��G��_�.�O�>e�`$�AM`� ��s|���_]���9�^�(�tm���:��M��պ#k���|��ńz��<��v�h���-�*�f@�M�"mTܮyD(�$)j��uO	;����
(�<��>;�*-�(E��-Y�%=�;6p�35�L�������
/;���l'��U(�Y������j�M���(�O��L��dځd	H;�(�8�{�@�N�������&�k�I�KVI�������{8�) ��ӟil 샇��V6� 0,�ӟ�m�5�W l��P�\�]�����4�Exyn�Rd�ŎZ���j�k=,w�KB����P2������Ҙ��H;e�۴v�cp]Z��:,�h|�^�35ecy% κz-��x��{�_���* ����{|iHW�B<��2���ʽyQ�Z������B�A��X�:��E�^6uK7�'�Ű����������}c�H�ug����o���Q����:�-���o ����X!� ؀��{���>$�� �1�n�!�.% � E�`m}�>��k�x2���ؽ�X,�?߭9K����"�,���J!jX����<������;!����ޏ4�tt��f�c����(�4�~�]�d��>��̂�3(H�4��i�P_F<0�6�����g$�z*IY��l'=4��-��1B�T*�-�Y �m���kpj6����k��1l��=ɧ��, �<��Ii�M���1H��3?2۞<�c��a��%�cw<���$5ǥ�v���C��4l�� g�6P���S�۬yk���۞?��j
a���(vU�a��b;=;5Z�B�aP��%�.��yϟ?g-w�J�tO���E�
����䫻n�6�C3���@U���T�YX0=��5:/ �&�%ڋ�b�rZ�V�%-��;�W�������;GTV3���Y{�q]�k��[c��Z�+�Z�,,�V�7)���&�m?(m��ش�Tx6� ��y�ɓ'�tx��1��>�e��tagM�s�ɏ�$�u?7Q���<y-����/V#)#�[�n�C�oӓmZ��mѵ�fd�;=��-���8����G�o��h�@��IǀJl���?����n�ˎY�eWuH������Z2�+B�_RE���������#�<�Mr��nH� ����%׭���W��F�7o��g?һ��۳�tr�1�{���#�z�o�mj㙑��WU�W�С�/�3s��K\���w������ͫ���2�����X��N�ꚦ�t���N�?��#E��MW�x��}D�]K[EC�w���������O(��8�����l+�_�j��|�7N�XC��a�{D�̑ξ���q��1+`J�u%j���k @pb@0�o�f7���}����OlYlc)��ӯP(a
�w<eW�x�w�q�Ȣ��?n���gP�/Y�AP���X���6	tw�]����f�R��>
���X+��)�=��X���W,���^�����3b���V�� �G�����ik�R��^�߮��@2>�p�n ��E����~V�w|0 Fb� ���G�����KP#�M^8��7i�_�sO�<��D�_�������q�xF�Q�-�g�{^�6�뛦-����[hN����x۝P����A_9>�\R'���6v,U=�R�v�]J'9ͳh�Ce������*��I�*$�J� �Z?�'Ȁzf qj��D�_�x���.��M'g=�������(�G4'l�V�3Q�i�[���R�Y��^=Fo_��޽}n�+��b%���a��V�"��c4�����!e#�,C2\3�1�<����E�V�F��ۿ�צ�W׈s���Va������bc3�Ɲ�;A2�:k�ף��.2��G�vGfƜ}���s�#[�D����)k�r����:������Ke��T�D	���z{���sx���s��'�ܼg�/�ҡk3�����*�5�����6B -�y۸/��mܐcᩭU_�We�����+�=ZL~w�j���'�t���N�쀤_m���+s��-R`/m�����ehO$��t�qh�RA��)uYS�E�`��a�A��R1��z���W��,���������������+�"U���PB�m?�/�<��ށ��!oe�m���2 �G�h<�q���w�~G����J����b<@ŋjT�IQG<V-5fMܵ�h��?m�hK[�'�d�$뽛�l�Z�8s1������9a�V2�L'|�l�����mY�0���<���RW3!����g/I`�ؐn/_}���|��S:7 �����B����Cn��n�sq>2���&�)d��I�:{�lkݱ����r}N��]�itqM?=e �+���G���@'���l���`�w�{I���� ����s�.(3�[˺�',�M�,�Z[ws$�N�=��{�6�9e��,�u 8�w3̳"�ԭ��O�r������;���|E��=�7����rO�~&�'�a�ν[��~�<���Pӫ�g���_Х����i�1X!�`�0��*.:�t~�Z@���}u.�M�!����j�o���U � ��d���mȵ��Y�V�r	
-�}���c��9���mW�w��q?~���Q�)e��0��}�+��=>���ؐSohQ��1k�L�>l%,IWk=o88V��b�"���a;��=+�"ʪ�W��[,��� N�'���a&��C�
@��b��x�&�W�
�?ȃH����#���JY���i���g#�<ýn�py�wd}F�[[i�^)��g�^Yo�9��ݨTk��ΟuOU�r[��(��ӭ� k"�ޥ8<,��O�������)�.�c��dc��k���������ך�8c7g06�8!��=5����%�ׯ� |Nd�2��6IQ62m\��s8�t�Sw�3���pB����iu͝��gCs-�o���+3�3�#��\�1/��]<4L�������_gHtMP_�ڴk1@�����.e�P�������sB/�4�녋�,^�4�Ƭڶ[%|ܦ�'�G3cdp��%ǡ�����ڌňH��bK�,j���m&�Wiw� �NO����s3���6S8� ~E����;/ n�?s�p�&���ʻ���}Ui�}g�E0��8�M���:\�b�M|���K{���}��6	�M����~.�����EK��i_��Ǹn>���\THVŹ��Jy<M���
~��-�Y�Pk5i�6-;��O$�]��駦�i�#�k��5���5Y\�O�^���[|�e8ʂ�:kp[��E�	�}�����!C4���_��`�y�Y������`Zm�׮��U�Q(1P�T2>�|���/�VƱ��뜛�5B������
���}�Rh���ux'�kC[��"��#Y,��7�b��!&@�1K�������`�n��i��Sn�"e�b��������z���g�9B�UX`����]��x<�{Y�m҇N
@�'�j�9b3{���\;0�I�l+٦.�U�-���і���@-a�!Fv�/^����P{�B�럘�Pn0�D2WJ|W���{F���f��4-�6w��*�����M�t����'t5����S3����O/9�֭;k^�X� +I���kV��]��?��[�o��L!c�6����O2
Iu�z��1�j�-�?�%Ƌ��^�^���y��y��XT�ްO�+�M��^
�Y���2�v�-(���B�jͭ��z�s�Vvs����@�rߕW2'��I�d}�5�ޘ[�u���c-��<�NG��.�>E>T�!�Ķ��D�ν�)��-w#꘼����-��I����	�����{%0L��Ӯ�����}q�jl��xF0��N,@0J�	�$.��λ� W)cD��"��0�=��K{�J�E���n�o+����[�I�d2s����r\��m�:vY�z�b�#V���o f��[X��͂,X�r%x\ZR�Y#�l���յEk6�3ܖ�Q����X�x���t���#>ׂL$�bwU��*z����^π�	����uڹ =[��,�c:tx�O�fKQJV7��'�+�	���p�<8D�`���&ߘ �:���E��]��<ӵ=�o���gc��J�,����q���z<���=�MO�E��iQ�{ �h
+D mh2��|tI��z<�����i ,㛻?R�3�;���\@�!�� E����'�|�-�ɘ�0�Y�����Ґ�϶�ݠ�}�2ob���r~�wݢ�tN۾�m�+�4���yw�6%|jU���YY��>�[�9��K�`	��6�b�('	O��K�����OA� �r�S�sK [S��E����Q6�B���d���W�����j�=Nւ�=`���]�E8�?m�Z�����:R��;�C�#
���� K��]��� �_��F�v���1�5�1|�
<��IX�^Wd��*��0.�)T��P���l���{ ��,Ynm �D�S�Һ��0��`�3 ���0�\����4��Jz�қ30v�S��R�j��4��K�l�=X��m����}��ܣǏ��� ������tv~�n�U"qV�><���G����3^a.d��`�+sC��t������0��p�.�4�$�x� �),~(_���ޣU'��b�h� �!y �H�ζ}���Uц��C��qn!��os���R���L�.�,�n��� ��EY��M� o�תX%���J�NZ�UH���iG;Z/�j(ZY�Bn�=��8F������`�3�v��׹.�N��=v�P��Nok�T�v�b���	�Ӗ�bIO"0����,�n�� �P<~���M���<;қ�4E8��N�
�UQ�u^�*��A�Pu����e�;��Ŝ�l���#HR��� ����_�U�����3��t���&p��GWQ3����gJ��7�]�* ,k!,����+�e�C��}�.�(�,�Z� #�	,�(g���JB�]Fbk��ǺE3��4.TmH^[���7������Q����]�~�K����!�e�{B�?8��~Bg���̹%w�ü2�~j@̐�R�6�g��z�i�S��<���K~�~R��
�c̔����SǼ�H�o�/���"�����O��S �{f u�'ty=���1'�b|;���uS�Q'���G��C���~o���f>u8S����5X,|�� d]��������mƂ���,��6R��g��u�,>����:,$��6�w��Um9��~�: /,$H�0 ��O���=�U����q_)�!��<^,��
֤%���-��B��=��*O�����U��V�9���-1礜�*T|�w^ _��M�y<P��Y<(`KǪ�c��A�@. `��Ѳ�	�g��4p\m�^��n?���0{w]r���T͝U�W! .�-k��d�ߣ�����on�_��S���׺����m 4�
�-������&:;�^�KG=��!���E`�O���湸���|D����;nb�ؔ݃q�����
���~�\�
/���V������DC6@�㘫�+z�������t|��S���O8IVw�؀��i��@2�<{o�ҥ��:��-��	���#����������l���sB���n�(�b�B����ѓtr�o@p�	�2�y 쟋�Wy7�bҲ���i�G���)�{F�gׁv^��x�(���us�W>��=�~�G��Ѓ{G�����Й!żR����".4�_�`!�Ge�2�!�*�_�9������8�E����,׺u�Ԧ>m�����!��%_��v̚�e�5>����J��̜Z���B�]J�_t���ж�R�� 8� �z�������e����*Û���D���C�?�hk�*�(��o3-��^%-,� W<62��d)��Ba���� �ue����p٦���u��Y�y�" ,d�bLd1���:�7��u��k 0�;#��f�+$i+�����و^������%��I�����'��%|�k���s����M�uqy���ɓ���������w�^�� u:��w�2 �
p)���:��t�St��н�}:0���Ib>~.o޾r@���������
@�� �/���>��!죞��و�K�f�!ZAe�s�Y�ɤӧ7�(��G��8���xi��&Hd���m�3��59[~�?��?{B���#��2�#����Z?�.�\B+sM&���d�M�A:=��go8I �]�*�(�]��^�x�hG����go�}�^���|�u��Sx.�.�E���p�&�sUr`�<0k���U��W^�jRżz=��E�b˄�������YG��K��^�xx�[���3#��?�B�)6�"1��Jji��6�y�{��F����-�~XVEun�m�K��b��@�v��� 8fE{(�9�����^G>�1�a)ȸRh���I��:������h;Ƕ
 3sG��j1�*̙��2z���[�,z�vA�w�}��Cp}��\\<O�5�]մUk���ٛ;N����sbX�PZe�޽{��]�9[�x<◬�����=~t�ɪ��s�:�Mǚ]Uq��l�
若�t� gl�>�S��GX�R� e�T�>
�������\Oq��o~����?��Cd��M�H��]�n��e����$��:=J{����)'"���z��W�V����OK�f�x���@�w����\y��}���>����W��c#pe���X�������o5��K������]\����3/��g�^ޠS�����.�P�����Ў�:� �Y~����������#��u|7�C� �&���x�t���ڧn�ʬ�}B�VIxV����eo��߽��y n����ާ����PT_��rb�K�*��zl�5I������䄘��]�9I����n�܄}*t�^���u�iĴ����k]4o�B@&ٷ� �]���v�^�s�m�(2l\i"͚��}Z帇.�x�]�����j�Ē݆bECR�c���I����:BU�c`��5 غh�[���x ���PF�AFgX0�V4�E/��9��8q%� �|f�P��ZE�o3I�2<	2�u���ЀƇf"v8�=ҩÚ�ec��m��(��%,(���'g4�I��A�̹枲�/Jh�]�ǔ�Ylj���sooL@/��B� ���>}���A�0��������>�F��MR��e{�R��{|=$���3��S=Y�� u��~�̺:>.�'�} �
N��Bsj��H��c�"���}�x�>�� `3�!��"a� �{�汛 ����q� ����<W�*U���{[+Ǫ�p�u�6Ӭ�K�!nG��S��Xr-_rq9���/��{�ߌ��aC��M8���w�V��=a�q���iVz����Y7-�,w�	>��?z�����&��b�4�6q�=13�}u=�����~�ѐ=���S�* ҄CS,�%z���/l�*Y�.e?^;>�j��3��T��MV���X���n�w�i�i$�+/�P����uYR묄m��n]񠛢���H&�������R�2��Բ�F/H���2�3s2e��}�ձ�rOM�PF����i�N�|��j�)!m�4�\��W��)��A.Q�(��$gX��r��rjk�r�bWI���7X��l%wT<��h}�	�+�Á���yq�w�O��_~I���_3 �%�/�}��w���c3Qw22 ��3>��)��;�3��A/��#��24����ed��A����:�(3@8��Jܞ����,R�{3@Y��G�S��zi�0��32M�9c/�X������MܜUBcX��NL6�.��p��\��Ugel&\1�
c&����'Ǵ�| ���B���k�PD8变�A?e:�����Ni4xE���ޛ�����_҅�U(�RH.a\�90�j6#��
�����>oY����VP��������E(��"�>7MwE`��,�[�?�\f:\����?1�"w� a���jОo[�i����r�^�xO�~zG���\�-e}r������׈mԑ�-_��7����kz������G����^[��j*TT�o�]X7h�
ӫW����)�/��.��";jq�����R�*���սǡp_��^X�g���y��������"����ȗ���XG\�:i�Ko�)&�9��^cU�	ᗢ(»��p�v	������;�F��kK�:ㄲ~r�wq{ 09�+�`��ؗz�?qI%�IA͑vՃZ�
��bW� �/~%�f�b�t1��|��ă�)����1�Gw�w$�:pu~-��9���c�י�ў�=D����,�HX�h?I	Jн��ioĵx'ڂ�<w�����0��9ԅ�"iR>�2�Ź�̵�Vr��`�B"H능l�erIŸ,�d�l�p����&�/�Hrzw�-��?����.M+��Mb\��Ӽз�Tq*�k-(vL�<v��̀a�ز����)xd�%��N�bhl�<�Z��06,��o�t&�'��TŤ������u��u���q'��!��!������ꊞ>��N��ɢC[y��G��t�I=o�u&a��4����޾���`�������m��g(�=�M�?��	�����)�,G�{�}G��r��E0$�4�����!�_9a0P�;�G�M7��,Kn�����ڂݢ��u
.�H&���#Ń����:�Ўv�s�Py�܁
40��u��];��������p���}��-���W� ������y�k�Y���+ϼ�?v�w�P"��=8�	��G���40�/_����`��$Xo߾��� }g �QbF��O��#�{�<Z(w��k�}Bz?5����M�YBW[�K�SK;+��RN�ȝ�w�VCN44�@s=�B��ʣ@����H p�w���$_�8���6�q@X4�v�m0��pU�-f����Z��#�;<��8(�
Y	�#����LX١H�o�ح�b\���.;��ݤ��N<��/� &��������_���&a%�R(e��p`@  �S����W�������g0�5����xO|guYOJ�t 5�	�,�)�6���Fd{
�[�t[kh�[o��Z0W="��u�~��lL@�X����. �e����Z7�˝<V Ϻ�M�a��_��~HO�<����Z~��.�j�Q�-7��kn+�#�$3m ���M q��g�PJ1�<��y-��H�]�_��4a��R�k�p8�7o^����e�o^����>�{����E<�Y[RB�w`���-\l���]��gwo� S���9@� '�mY0$.Ѕ]����ef�����7E����'E��XE�C�Vjx��Y�9�*g���o����b���9?�[���*?ܸ{+�ݧ:��,�;�%t�~������JnT�]& �u��i��-&���[N����uǬ�I��fTȋ�j��W�8�p�iN y~1�6��=���e��������9X7�"�F��=�X����:7�6<n-�JB�� � ��_p�(�O�'I�ns�Ͷt ����5�
 �.��ߛ��b�xP<~����]E��7q��*�kr��[f~,�\� S�	^�wb"�V�ׯ^���K%�%(J,�F��p4��ْ����i��nJI�7�?b��g �ht���3d�bW�:�����d�C�@4��W�;߉׋���ovG;�юn���(rH��+�]8I9:�8 mLq>�ػ	9rV'�a@0�7/���M�G�� ��y�¯,��xl�Wo����l���z���z�p~޸0�-,�Q 0�j����X�do+��9�[ �7I��Bu1�M1�7Ia� ���]IVl�:v%F��&+k@�{Fu}[�Q.l �=�F� *���}=0@���LPhr�1[M���v��Ui�Rjq���+��^�$˸�����F�!�(���ʝ��{C~;tq51`:1��\ܳ�V	&�p�E������fZ�k���tIXrF��g��0�^`&i}�onGk��y3ˢ�֭U���#�\ ������[�Ni���a-D�Ԛg�}�y%|�T(�aI眚�m؂R��U.��j\��Wr:M���%z}�-���[��渀�8���g[���b�Jt�̍ Qm'Ɖ%-��@�������[ߎ��?�Y���֍�{��\Y�k��HRkbU��e���ۺ@��� �=������.ϼ�%���A��l��̾PV����J ���jxA�~��N߽���uSd=��y��ڻ)��\�I0��=�ܣ�{��	�����t��JӼIp�4KE1��������GE�\�õ�0GeA�-?��n���h~
����_|�M�5�� �-��������*&�_0���H�N��r�
sbum��yVW���Ԗ^����s�pK�G�3Q�+;�ں�$9���b���`�X!@kզe�eig^��-���W�Ǳ��^\U�Kq��p��;@2�
��
�&�>�緝3[�A�"���f틘��Q���ZSm#^���6�D�t�Xdy�6� ��y�h4����N�.(��{L���p'  ��IDATǏ��C��Nґ��y�$Wh	BT�K��u�Вv9˳�O������\���AY�����Q�7]���q�&�[53���Yi����-�&�Uoem�+��y��X��\-j�����_�ƶSs�:jc�X�B�X­���yc�Ib �̒���ַX��u?zK��Y��B�<��~F���R��[K�}qk����$�oTJ�}V_ge���
�����ϱVۨ���S�/�D[�x\�ܡ�Ϭ'��m��Y�x�`�E����H��U�Mx�� ��m�a�v�{h⿷Q^�I�b�+��1���Y x�,T$lO��K9^���;|Sq���͋�[M�.��ו-��O�� E)�P5�*l[��8Q+��6���2���K������>�꫿���������	�<��4\���˖�VF��s;�w��b@Ϟ�2���&/�p2[O/�Aܨ`�Ĺ8Q�\���K����UJ�q(Y�o� �ex�i0)؊�������z��{�W+�G�_"ĕ�y�b��?�/�(���Y�l�y���,�|�"�-���(�k]���>��-s���f(�֕	ߥ�&h�4�Y����~Z*�J�~ ���Ǝ9�Y�mRx.qu�[M�[�['�J�J��L,����E�m��֌�����T
�����!+F���)�g-�R�۳2L��g�׊��Q4�[��mg�k�M_�����SP�zg��F7M�W���{"�����W,�U�a8Dݽ��Iӳ_$i�"���ph��Dcmn4lm��n^�m�D+Bhжv����EH����v[�����������s���h�HO?�ý#�6����Aq΁H@���9�����Wf{�ɸ����F��YS��a�HD�PE&�D�s{5</�S����z��y����Q7���8���r�^�� �����g�j�CʲP(�i7~�T,Uq`H��{K������`~�]e10��ء���k�<ks����Պ�6B������}@Z[���������]��m$s���A8�v�p��g��h1P���5V
��pY�"@z"s��;�$-Td-�Ee%�v���{*:��A<�oۜ������C�+fU<c��"�?���eh�mnr<o�\Z��@]�xS� ��#��� ��WT��� p���siR,T��X�z� ��b� ���k�i��8�d�G�F(,�X��qF��C��W3�M��(p]3/�Ρ8���g?>��������s��O���Ȁ̜}�t�>A��y7\v�N��)6�~��5����a���޼}c'��iY�m���i�ȁߔ3J{!{��n�"]����,���r�P���;��:P`��⚷.jkl��'����=+���c�Em�/_2_A��* ��7u�*:�⁩�]e���ZP%��e����mGm)\���y�n��*q6�q����(	EY�˒f�,`�).�c�?�K��[�ifx��֝�R�����C�C�_�ue��q�s)T ��^�K��0�%��(���uΫe�6�ߛ�C(��*?/ ���<���0T#망i��8�h�����/U�4�^u��� u�u��~��M731C�E���p
�f>�_�[��������hL��\��\�£���f�kr�= ���5��h0�7��3 ���~���b�����ٹ@�j	����h!���� �����VZ;2�͚��c��tcL�1��@`�k?s��������H�q�X��g�
�謁[U�[��Pݩ��n�c�_3Ӿ���:�aa��;=��T���r��}<x��k�I��*�:�Np�@a[j�%�VO�9�ixm�
��M `Vc]��|����5̆B��-��<Z�7j[�݇'U�#�& 0�׺������n�=��wMO~��'#ߜ���& <o��Zy�𖝷��u�G15�����NHm���O(����}�'>|X
�e%Q0���s �RԽ7M�}^�4���)���%�I0�uM�@�pPӵ�s��Е���6�`K�\�: �;�1E��ޞ�� �w���� ��(6-�Wd��XJ�CKzz~����Vz21�S��d��q� X�k���Bn;r���%���b�m�'�^�('��K���O�d��S;U��q@����*)�����8&����C�5+���9������;��B`�������|�_� ~���k�����{[U�H�6vG�������I+���#v��^1��4���W�����X�3(���{���������%����n��VgM�KW��M���p��@v���@�|��|X��X�*u�Zո����}�V�uS�۷�3�pH���,J�=y�~��_�o�[:88(��u�e�K,�uJ;к� ��ĬZ�����\g�w�R�PE��������S,�3m�s��l{J�i2���<��sU�g��q��0� �`l��CDEr+P��Yk�+��;@ �������&�I��H����,�s�����|^�As���T+������:��xp����t�pd��lܜ4���L���2mZU
l������7�kps �
�/ܠ��*^3��5}ެNE�Z���_����zA�*yf��i��mh��ol�-�U5?D�X�[x�,�i��&����Rc�,�����@Q����@V�ťN�����oD�������a ~��-Tf���3/����_�M󰛼~���V�~�Yz?c�o�2�<�Z(ѡ8��W���n�{.�6�.e`ڌ��U�j���s���F1_7�Mc�n������J���k묘�{��!�$a�z����%�
^(����،�i�G	>��5Ā������o��69�pd���;�S嬚�z������*uu�u�ݩg�m]�B;��p�%@��To�2QbR��.���
'� &���J��ط�{��oW2l�7*Z��ơ	c�[����!2n��5�뀁l���Y�f�6�8n��_��Գ���ΰX���O�
�@p��m�\5���B����;n�:o��5=n����Aoӵ7fѬ�����m����x̪�1�(淔�A~�%�<�]d]�y�W� >˒�*�q ���e�R5�U�1�Φגp������C~w&�J�p�F���f��rL՜3S7�GxݦR�~_������iX�P�&U�w��EQ5H�#o�m��Ş��bm��h���.�~����EK�G]��~�k��"8�'�r�]�	w`y��;��������B��)>�������XrV���:��x#�	��9	�]��cE��`�f�_�y ����6w�O��U����Q�f�<���&T��U7�/aM��\�L�E���e��X#v�+�])�8�S7Y��LҙqF;5�ϱ�T��*�em?T�E��Yc�hz�\���v�X��nD`/�7��w��,��h�[ъ�[<�1��V1� V	��VA�{�d�j��Ze�����zm�c^�gS8��� �ȷ��m��(i��%�?��± ���=���- ��7똦k	@�n�m�`X�X%�st�w�c��so˚Y�����[�����=����6Ƈ*t^�$/U᨝���]�5mH�r�P�[�q,M� �'kqe�*E_%(zbL!��c޶Z 	���OB���0���jH2s?}�K���vm��ɤ�����u9�6-�ߖq���c.eA��Yk�l��$+�0�@Q�纶
 ��$��}!�5������뢝�a�� �1nI�>�j1�u�t��><��23�,B����]sl���bP+sBs�,^h�$��I�3s���wb�ʏL&yq!�	:�����.��w^f�����-���z�>7[{�`�j�h�mT)!wT�Z��x��Ti�!�߿���%����P�|Jf-z�*���@�
8�@]-"��=wV"��1 �1��1��$C���}�By��dW�P\5WB@Y���ϯ*iP[�y3��~����d�>�}���y ze�*�	n��dU�W����3�����%4eJ�������RMB���y�^�|�)V�#Y��;	Z�dm���݆l��ӂm
0�<_�/�[٢V��GV��zN6��A0XXlSJd�ݣ�c�q��������0�S,�|��Zٖ��sMin�p��1��.��ɕB�_zn��a��]+�Ǌ� q���Y��f�v��٠)d��Y�K�S���* Tk�os�C͆��Jʹ{�lm���wHj2�D��Ma���r�,ܿm,�,�p�7`Y%�fׁ7ܣv�w��	9���r��y,�8u�eX��|��7�P��-���j���?+��P�����d&_|�ǇC��E.�Z�`5'#l�u x��R��-� ^�|1\���2�B������͢eyH[�t|l�E+n{n"y���x.���c�}�|?�:vS��Z7��-���SB���0�J����)��N��p���U�͢� ���*ECx?��(e���A٦�涓��[��Gg0fq��%�R.�1^�^�G�������I��B��9�_>�\n�e�MFe��i ��l�l}Ӷ����pZ�]n��v~�&+B0c�����Et8�5�	�EL�v �I�܂�ec+pf�@K.�|Y�ۅo}q��.��'+.:=�����wߌ�1e`n��z����צ�#so���V+~Ia|z<f�މy�|vX����P:~�VI;�z3t�o�6]�!�룏>�,�O�>e@Z�I�9R��U��y~����Z�w��E���I$��'��?���ߺc�E.�tw�q!X�w�8W�h�1(�cߤ�	=>@Un�!�C�o8o /�ਲ���P��;��
Ae��MS�Q�4���1U�6�pn�Q�^n����(w���>���'��k�e�ç��h&[׀����D��c�;$E+�B% 3j��W�I ��qF��]_O����J�j;���Q�by�)�X�JpQ�`~!��ú,�x k��J\9�� _��26��-��eb��6kxʥ��+/�-ψ|�8>Týe��.�s:7�76���:	[��Ô�Yb�k���I��\���n�N7�~_��@��Մ�v�n�}��:��&h��ϙf=��f1]�� �=R\&߼yÙq��zs�c�v�9KX�9G�$s	��o�=�s�`<g�Z��C�,�;�D�]kA��F�u[(6�.� `m޿MX��='�?Ck��<F�u���MQx��gP����X�[�Z�1�l�Ҝ�L7���s�h���=-�&t��vhA���:5��K�W9=~J�^��=��wYî��Jܱ�%�C��M�������z��./�jO�$SΝ��F��Y�V�<��bY��XSW�o��pc��t�7� �6�{��i�A��`������i"�րh�N�n��_����,�E�);c�����޼��~|KW�#.L_3�A8ш6c0@;2�0q��3}+�gJ`P�?����Wo��s�H2C�{7;.�zZ��/~m�����fS��,�.�2QR���~������-K; |{H�)ܞ�������!t��U�g���`	���ց�*+c��M[���-��*iY���R��v�i�x����]0o��/w���C ���k�{���x�'(L�ؖ:�wb�m��=g��я�MR��7(���)[ߟ��^���+��X�4��D�Q�$�,f�­��ߧ��=��5��]��0
�}���ko�O���^b�u�Zpϋ�w��tl�S��g��M���X�\0s���� �o�����9߷��;�����XDߟ^�ӧoL�:>��;d���Նa��93L;�~%�b�Ŗ�p��Gc���kz��-]_�=���x�2Դ����P O09?;�/^�4�m\o/�//���vs{>�y�u����]�!�ߴ��j|Wu�M��?�7� �:�$%��̺�.15��Z7I�/J! � Fȅ�x0����*Y�&(V����}�V�����P�*��*�3KIS'ޱ[�: � �!�V�/�`B��;=nT��/����n�#{�})���,���Wtq~i�ĈO�����Ⱥg�ܵ$˵dHՌ��y%��?7�}_�x�>3���Sz��=g���v:|���i'�=KE@�,�T�d^���^���=�hx5�W�^��������Ol�3%��=s�{W�
�bov;G��<ewja�Ht����������h�i�xց�P+/�����$~P~[m^�yH����vJF�Щ�Y
]�b�����L�2g)8�=�H���.���u��*˛p_�B��/��O?��>�����]���ut�<�(�nz�����������z���3Ύ.�-��Ibº��{�����:����yМ�{��oU!HU�)�?P���� ��6G����ͅb��_������� ���zzv�`�V��E�-����K���4�״c��:=�(r�֪�M���yV�l����Z�E�#� O\",�����y��	=6���� �ܞ*m)'l �ggb	μ��]�����X��;7J� �.XR��YS�����Ƒ#�߽���f���
��ǋn�����B�����7ߊ
z3-��w��.�ߛM�;��b�d�oW_3ֶ޺��w�`[��p�d3��z�,��s	5�X� �n�l9�m�:jZ�b��GY6��(q��Z&WI��f����/��EI��u � �����})� �s���:��V�_�ة���Z���Z�C �^7��l ���|��3���8M�"#��_��RNmI;+j��Q�j<g�U��ڲ^/� �eB�U�
E�x�r����Y�����b�]�Wj�����������0��6�$��F�]rμ,�ߩ�Q���=y�1����2% U\��舾��+z��	����5zC�ܰaAz��C�h��rO��^�z��?y�s|q�dX��e�����t��ý��aZAp����]�d�ơ��n����Du��/9�j;H�=_\ ����Qae��P(����vSv�fK�� Pl����&�md�WYX��h������&��,��i�g7 �oq|��"����,A��AƖ�E�����Z�W�F�ժʽs`[��C�9K���������_���` _�֨Rf���3����u���%�l���pS�8"1����yyI���o�o��������y�Y�DYX�����jp���^����y�si�o!��]�5���w���K&����	�W:��U�ɂ� �ժ���7ES/�mcq��"��;�@1 ��{'��ч�2�z��-�{���{X�rj��p@����W�ىV�K0v��eJX`�n�1���B��my`�U�i�lo�U��sPT¨x��+-h){�E�c�~�ZE	5��S3~�Q*ϟE;�U�g�u�νK�~��t�ˮv�i_���B�[��J�ֈM���}oj<�ʚ�/���CI$ ��\Y��&� 8H�J�x�UܓXA��
`���~� @�`�&U}�����mr��kĥC�L�q}��1ˊx������4���ch���o��^�&���I�U��,Y�����uZH���\g�wdI	�5�Ȇ�b(�#ߝ��JQ�0n�:�ؒ���K�,�`�"Zf���$Z�_���V�����Bs|r�e>��S�����5����z�����z�q�\C�҃�9>��'� �������Y��&����BS�{��8�ݵGÌ:���]��8�5 �:�p�q�k�G�=H�q;�_i �|��n��I
�;�CTrꄍy�\�H��x∰㳀Ҏn+U�P[�j)kk\V��&p�J0�(��2�����_X~?��s���'���K������na|�r��̖|X�%~��L��F�ڂE\\�1��@r�@�k�I�W�.�y>8>,��U����!�S��L�ձ.�d��;��3��.�9W��-	�X� 0��<|�Ȁ���B��6��-��ն=cm�t���4�Xp�����|h���'�Ё����w���O쾂$��
�� ���/�+����&+1� 6@3���ѱ��@�R�˲��O��$W6${`�?��]�/����H$����	(=e��V��ZAgZ{wtH�P�za��uߧ��{~�Z�∙׍�AN�L\���*�1���n��K���Nhn�碖�M �y����*�6�^�u1h���An���x����_��^p��,��߿=$�S� #0�`b�Q�r.b���B�Z��t�qjZI;K��ֻ��:m����=�P#���Cl貪,P.9P��Z\�W�M띠eR���S@�ï���&2-������~qR$�0���l�F{ ��Ȟ�����GvW���g�'oY�Eϴ��Ȣ��_�yX� x�����>���o�QH.[�" �����K�K5G0Տ>��ƣ1}sy����KևܝW���&�o�<���3�����m�J�-�?;Z��\awtר��U��0�c�ߦ�6J��+E�_�_K�~\�}JL�����T��;��r
̒z�g)�'¨��aM�*gh��3�7�S|�6�o;��'�~��߲��'P�yD����{슽J࿣Փ�s�cp�Ki+�7���l�2����,����Y��-��~�֤���}�	��J_���;�^�b�������f���ό(�AR���[i^�_ ��"���i��� ���
 �o��{������������꼷ק��� ���c�$6���Iܺ]�H|�^��is�X�a�M8���������+z���(�[z�D% \��ϥ��VW&E��{�|x��Ѳn�;�&
]g,���Oa���vf<AJ���.xn�y�L8�}>�\��γ�NQV���E��q��??)��J��.8�E��܌e'�P�,G6l&��*r�����V�rK�r?���I�{$����#���X�b�K�3ps���_|�{qUex��9�&����7������w�"��e#��l���4P�y���Y[��O��u�_�s��<��; ��'�a���@H�q��r�i)�m�m@�7o�����O���Q
�+��Teͫ���B�C��"
����P��pa�:;;�L~peN;=����s ����?<���}fb6���Hm\����j�YjA��p�-g�I;4��9]�]���5V����r������n����u'��\i��[�G���jG*(s��F.�C��>|@�^��F8C��ꛏ�ْ��j[Z��P$5h
�R_�};Z�T�T��>ծY3�^ ���%��=80�{�OG��v��Y?6㋱5[��mB�̭��Q>��uy�mr��y����C�禸Ū}U�:�/�������0�m��O�ϰ�?��(�VdV$�Bi$l���yu�y#�M�ݿ8�x�1M�{Q��6�e��?�P�����Ք�JŻ� ��Iv�J�*.��o�z������Ir�������gR\D�2%�a������G8a?�[��H�����3�w�^��s��j魪�󐘪FaI �{�=9�
��K.� �p7���D^p{��/>��98��|��Q�E��D&-�h�8�nc��"�����O���.j'�7��9��R��4�B9�A'D�0�e�=�����|�և�d7�w��I�f��c,��F���)�'���-��y��wNF쬓>�bk_���މܡ���o�s"�,lI?���w>�Py���K�"�9E�*J0_T�z�K�u@��>'�kwz�ht�{�A�z��cZM��#��y!,��1=GD�ӝ�0ƄG�o!,�9�<7*��S���-WPg�H�<-��]ZZ�9����m����P�ݥz�M�5%��բ�w:~_�:1�Ћ �#lRd���O[7.	N�F׀��! �H�����.��0��T���Z�/�d|�Ȭ���?d�0���+m��dfNVh�zF�N�����CY�i\��	K��8���hrs�Z(�$�)˜�<�k���b�O(��xK�)���%���~E�8$�YÕ,d�jO�z]�y��k�N��g�P�q��vL�7%��x/�������p�����,W��0�2,?�gV��^	�qH�}\��6���n�.L^�W)$�_��$X�S��xaT�ۉL��,�X���']"�]\������b�Er�V���m��Y���yE�攐V�\�a� �c�
���}ܣ��c���7���.�{�GA�Z� ���%u}}>�-��|2𪼣��܂n%4t�4�V���_!���]5o�KZY����E��v��hcc�����W�07�v��b6kuzt\k��w��ó7������S�ޢ���c!�,���)�`9��1�1�1�B�X�ָI,QI�XP6  � �����Ob����,]��i��4b.rδ�x��,�&�XM��[[[���͛7���Y�>��m�,�<J�c>gI���zw�K���I�ҷ�	�D��;��!5��a/�a� ΋�,C��|��P�7VMJ�.81�]5����o��H�8��gV�.���4�w�8�~�/�%ߟ`n�:-\T(KӠ��g��i��������$4��je�X�ȸ�|9Ő��/�Viks�>ܤ�?�O��2�����#/�s%��j�C!���^������@�W��ue��w����J�0pȉg��޸�W�I@�s�^��������c�����=��p�R�Օ%���=}���Ѫ�ime��%*@�C�t��Mj�v/��z�6�ha�����B�D��#��6���*�����1̀�m�gq�,�n��x�9�H�d�;,,���lz��$�iqK#<繞�6��[$s�D@e�=q#6����;-�<�	��u�s����mރ�x,�3AiH!���\�I}o�K��#L~IWQ��3r��'�}>��E��n� p[��� FH��x)�Dj�-x���F���O�}��/)�S�Z����]~K�sY.t-x���^������z��K��W����>�f�5��.��ϹlǏ�W�(��o�u؎�� _x���t)�$��muZTZ����e���=��_��>x�I�����2���{��{��9=*�Z�*�\Z���5E����֏���^з߾��V�r�yJ6�R�s���Zx>�/�:b�4�ָ�t�;��$@r�발^Ҭ�0T��Q�"Dp� x��in��9o*�b���,f���V~$	v���;���u���/z�d�8��N�o��U?khrO�Y�a�M����K~�&��4�q����H��ۡ��
��Z��~�C?��>}�t���<�^���=Y�eϡ�"�AB�k5\��*%�Ε��X�vxt�Hw��vO�	�M׈=6��Q�4�[;BÉ��:$�S}U*���2O>ݡ�?yğPXx^Gm����n5�|�|!�n뎧��#^�X.��/SY�	/�1R�Q�~�tQ=����Y�;R'���=8���nR򛌙�֯��u��n��#������uD���bI�3�Ns>OS<\���{���s���GK�-0��Gw7�{��kqQӐ[�bD�3$X�FhȤH	Y�������=���J��������<�+]��M�����)���8���1�0�c��Q�����yZ\����e:>����s�p�u��A.�zjg�.��'F	b��;Sя�#V,�?�B��Rɣ��yz�p���?���ޣ��K��	���ڦ�[�z�Ķ}�E�]*�=ʗr�sr�Ej���=z�pQ}ާz�\@�^�)�~s��0�i`�߃iӤ���srSI�I��k�1��0,y��H�� �x����������y�������vܝ��68^x����W�N��F���<�o�ѣ�������5�΁�6��Q����]j4�tR;����$X��r�DKT.u�1[�d#k����裏w�Pթ٬Q�7���9J����
�0�4�E:D��#h\&N�]��e��\U��N�Uo��S�U�n��}��#�3�x7j-��Z�HvV�C��"-,T���0<��|���"磏����P�����j_g`�M#���@�M+�$��h�A���xY$۴j��ٲmĿʒ<g�߲��m�1���5iM�*d%rKU@����4����$�_�}��,%�viq�� [XXXXX�hh��o�Y��9`�lu~�?�O��>mm-Q��)�Z��GtZo���	�����Et��X�x�R1G++����"�%b��n��WD������"I�{'Q��?�L�B� @�g��HB�V�<+&<������T)�у[���&���.��sۊMtYKǛw�o���N�f��kC�TZ]�҃���	<_�$��=�Bޣ�O6�	���:>9�V�A�)�O����$8IFMw^Y/�Fvk]k��I���M�L��1j%�E�<���$��V��f�qO8�D-���:��_�}�Z�۠�ɲ]rl�Ƌ��H��n��Y�u�� �98F,��ЪYXL��4ƶ����L���OP�,� G���HQ����igg��˼���iw�ޣ���y����1���jS��;*<Ev�ҪH�nHk�W�B]�T���2��A������En�`�P�-�B�����;��,��r��˻p/�dX>[�+eW�i��_�rV�"������:�����	�~�ϟ����kw��p�S��awy(D��(_�U�M�|�VW�����H�<Ϳ�*�6�$J�GV��w#�z�[�b\*$N>��	�5I�e�%!�f�"�o���q�d�Ba|��i��,����%�9�HLq�����T��u�O�R��'ˆe��,���&���	����tC����&|�l
\��"�?4@~���VZÏ2r/ժ�������l`��{EEr;��wD/^���GtZ�)��9�3,�ݎO��>���tzܢ��"�ꘊt�l)�>>-/����<�)��}a%��gd���l
��СK�?���a&,,��^*��P���
�wo�-���qg���i��W���~�j(%�J�+�%ɭ���Mj�߰|���
����3��E�qN�^�R�}=�l
�z�nvC^2��_����_&9����U���l6�^�S�V�?OOO9�B,��$�&	��I�\���^P�,d��w����8�A;�<����g�:��(+�U�a��%�?�]��/M~Vl��v�
,�S���gaq�a�'��D�:qU�����8��XB�<-���|�B�\W����"�=:8�Ӯ"GGGmjuHm�S�c�H��Hr�ۡf�ͱ�+�Uud�.k:
>�-���R֚������N���q��{1e��	��]�K?�\�
�s������-/��N�z����$��j���	���I�G�^�<E,\�H>��.�j�[u��]�٩����U]E44�-� ��/-Ϋm	!⎴i�\��!������{3��z�@j�dB�gL��YӲ�Rc
�����7ʰ��e����R��/����){��;0��I����N�lǰ��Z G����tO�'�*��R�I0>��^b۴}�]�$
�ˀ%�w75Ө�Y	��Q�vm	��7_pX@,�
Jx,)�Q	��Ԅ�d-%\���F�bB9���%u�\t\�Ndu�E١�i��&����
-��\��+QU�#��6"d��i�~�A�.��m��J���2;G�b�
��z���hw��T����I�<���g�����%ĺ%��P�[>�R�Z`2\(�T_lF|0H0��ݵ�_8��mW� � r˥��>)r��:�<�AGGGtpp@���꽡�q7e.��H*H,�u+�h�&��dL�Xq���[���O^�c����
�����ښ���*���ɼf�O�d��2]���\F%��'t2�:���ٗ,}�v�i��j�u�)� [XXXXX� D��W���A����x�� Q�Յ%'T$�G�f���Y
"G���t��QA\i�c���~HME��j�^W'X�� ���Z4��(���Z�[9�v�YC������s9���͌>F�+R��������F٣��={a�/R�!ӳ�����܂�Bk���A��[��i:�Cy�c�:dq1��i6���
���$� �X@zy�z!�x��+� FB~e1	�i�L#� �B������v��f��Y��k,��˴���V�d\�){ӈ���*�;��`������2s��4K־�p�
zK�-,,,,,f������~(� ̥��0ȵ9sA
�LёЉ2H(��9�����Vbw�6૯�Y�
�T2E�9*+�X��Q$�BP6bB�N̖�M��O��|��䗉��#��ž���]�� 1İ�C�T�kE�= tl�"���-�-�[�a]�yX��N�Nc����J,�@��NL�	k�۷o���������B	�+,� �fL��k�H�X`�R(ۛ���D���_�[m~W�wE�������A�<x@���lFے� �<�E�U@��]fR3����nn�Ӵ�&�̓m�Β`�%�7ӈ���%T�T�j1�p��������Bl'�]�&ð��t�Z��r1a��͸�v����ι�����5�S�i�Eĉ	sh$�	���}VmG�y�3j;���p %E�K+!���֫~v#!Փ}v��e�s5�f2���m|��LmG�҈E��L�����߰�b9>>f����{^`q�v �pA��Wbp�sOV�ai�I��6��Gbkp���a�LK.X��T�oKKKܾd|p�}�E\%>�6���0�n�*�W��\�u�$� [XX�h��X�:��,�����7l�I��2�Z\��8Q��AwJ&�qvT���Z	������X,!�o�ʥ<Anw{�� ѕ��shGZ%szj=J*�pY���yv��q��S�ݥ��^��-��/Z("���wW�ZxA�dtT�u�=�Ǻ����g��IX���gjpi�R��]�{"���$�+�2ຊde��~V䨮�E��-Td1�H��M�����DSX�����3����EzA(����	�P�<�7�֛�=�l�]���✕J�:�� ���m+B\W�����g��W�^q\�G�h}}=��j�=f�f��K��1,N�&�ù ě �+I��1ɰ��\c|\5��-,�	��d���E"q�MB����5ٞ��ꉊ"��plj�i1Y鸬���s��l�i9g�I�����E��-,]&��'�	(�w9;42�*rsx�V$�C������kA2�R۫}�W	�p7Tx�ʉ�P�q=Ez;t|R�����ދ3<��P#�J�����G��ћ���K��֫�D_	���"*::��>l�>����ܐk���y���r�����Z@�u�"����C�*e�ʴ�T�����2̈́9�Hr��j|�NZ�\Y���xg?�e��>K��,�%�G��ERe	�aڃj|^E"�a�<���j��E �� ��+���"'��4�Œlʴ����q�MM�X�M�%[���XsuH�&��(����C�o�`��|��%��΂Bع�74	֐�Tf�rQ�4S��Ŵ�K�4�K�ĉg=���MWk����˸��;*�[-��SHxZ���7F���t�2?��6��Q���C�l��01�%'���#q$j�)-{T����� �[Hj�RK�j�mj6{�+�就O�J���hKqo�������(�Wi�?�`�]���z�Vת��T�x�[d��(�A��:T� �w
1!h/����"n�]KY`��(ɭ�i���>�}�H{{G��\�b!��"����b^�W�j�������ȋ��1(��nR�������,���
+9�૟�^Im���a��U�v|��[��C
��)L�ڌs�)D7�{r[�x^Ϙ� K���� �F���B��:�x���;������b����$U��Q��Þ�d��%���3F�� ����?��O���kz��!ݿ����y�TJLs��ذv_5��<㌵a$XH�9��xn!��2C!���b|e`\B)/|G�;�k����CFү�`�;��w,.�L��tG�/�f��'=�hғ�ht��m�y�։-����?NQ�G���� /H��p�f�g�wBG�T)�T�)�V"��Y_]����v�
9�ڊ�t@����cda�L[��jY��Hz�r�l�yo���jZ�L\���и�0�Wv���8�Y'��g{���J<>n��a������<m�{T(X)Q*�hcc���m�I�6t���@���X(�=E~ѿK*K���=�8�Qh�}���@�b�H~C�0L�00��d�!��ϴm'9�E=<F�ݞ9��Ź��T �� �>��c&� �o޼ab��AA~�UY�h<��:��5øۤ��,,1�b���R�	�_\#�OH���_�"5���s�U�/d�J�|�Ҿ��R�gE�7s?��^#1���{����@غ��R���J������6),����u0_�����uc\��(��qRk�I��8�}���YL�k�PKM~݈��M�ۊ̞֚���;�XSDvmK�
�zm�MO	)y�\%@��z�����1��r����9ZSDu~�)���W1�v���#z�z�v����l&��DM8fK����,��a�3~���FD��A#)U���i�޽?�{���nm*�R�E������WT�Uiw��HO�]�q�R���j�V�ʴ��@ˋv)����z������{�������hRI��q���B~Lk��e.�?���×/_2��V:���8rL�q��[�uciy��#����"�R��O>�k��Ȫ[;H?]�;iXl�v%�0��q��s������=��g?��O��w�<�ܧ)R �O�=�9��~��_�5�aݿ��g	���ŭ@��}��Q�qc�e�%��8m��U�dv�y��LL[���[�:1�9�<�(��{_�~O+�E��Y�JqQѧ����7����bF+9j���B�J���"ǋ,<w�m%#lN�@�z��;z���N�`!��W���Պ���0��E-~׆��D}��&+��h��՛=Zߨ����*U�G�O��E��E>D�T����[��U����B��KT��T��C�`��%EvCz�z�~��-�W�{|tL�v�~Io����;�d\� ��X�޽{G/���7o�0!Ar+$���N���1q]��F��.���{.�$���^��5�qĵ[H�y<�.}�eX���O�D��F���!�e\~�~(!@~?��s��/~�J���f`�l���㸯�k��?��î�`�� M��`���{�	H�I �yI�!B�(�h�Ԛgq%�1Fݫa�b\Q5��V�a6���9�E��:��r|n�Ӊ�^�~�Hn@�����%%*�"�dש���ZZ�S���c#^�H�9���o���*ѷ߾�����]��5� 7Z���pŧ[�t^�N㡐�I]��Xr�ӭ)����sDk�T(�huyA_�V���iS��P1_���y
�\�;r��̩~���ㅊ0{��%5f�wH�ß���zF����V���9"ļ�b*H*6M���A�`����ݞ_��~{��",q�+��5���gi���}nn�>��C��� Ê����/�`+1`��N�3�z�,�0�<�q�)�� 9bcc������~��_�g�}������Cl/�.i9.�_~�%����-+g׍�`�%x����K��������|I�����Q�޴]�.��,��f�I\�Le�i�9�	Y1Y�
�0I�j7�ȃ��$�ǃ��-6кw�t�<��z�0W������-%�^P��E�C�)�ł���ds�Y*���@�K��Mz��}��z�r�j� hl��$8"�Q���4��XIq��1��'�8/�7��3J!��S�E���~A��<ݢ��2'3sT��.�Y.x9$�&_	���TK�ا ̓�����>}��W�՟�ӳ���ZS�{6^[
��1�[L�xM��P$����l�Z\X���U��W�J��q��B���$���B��1YY򴻻�����Sܽ��Tׅ������ڑ���Ǖ��f�[X?��c�������7��7�0y��$��`gg'V��z|��W<~��0� ����Zlaaq� �A褮�hy��9-\� �#�pI]Ƥ�vd��/Q@a�{��(|��&Y��쑒�s�-�E�f�Kq�G\7j�*�t�D���Qk�o�Ύ"���Y�Xp��)��j?</ X����[����Nӡ��N9zI�������`��k���
�N�����:�͞`}#`�J��0���3\�߽ߧ��N����O�ɣ�X_��{�~���FxG�����ct\u�<�~{@�����o_гW{�x�������!���Т�$�3އ ! �H*��<x@�+�� �bI�$���w鴈�0�wfb�	�p�G&h(wq�H�B��ӧOy>�V,���������˸�,7h1.@&��-������?��?�����-�f=�4��n�e�0N�? �p�	�LXlaaq+ /wLtpÁ�^�X/ZG�X�E�/B~L2�@��F}C�`�z9���q̘/��{�c#	
& ����ݨ�a1BW-X��B����f]��'��M���'��_	�8��i�C��{����.׹��\�㺱�R�K��::�4F�4Ԑ=����~�~|�GR����iw��j�]r�[�-��.y�t��f���Wp�7���}����^|at���=�C�k���zv��!���q�=X�����+Q)��v�]��5r��.'3kԑ�K{�-�����_�H�^����Sjt�'6�3��E/�{�����/\��.A�(�KlQŰX �0�_�"qT�P2��O2|G�2�1\3����m!+H�(˯i.��ܘ���dF�X�8C�����6x��'#��<���qpl�}!���$F]⁓��f,�$������ /F�|�م�/OyiW�a�q�o�`�aB�I����MQM�����+�mI�0'ץM@�[�I� A�%��Mr��u��SQ<&����3�p��jztrL��9�zw@��Uiss�v��hmm�����\괚������j(怾U��ͻ#��J�lR��UdW=_�&�~D~i��������x'y�}���뛦�;køt�u�q�c�l�\�
5�߼9��{O[�Kto{U=�sT�x��"񙣈�����C������o���7tttB�Z���;������	s~ ����C̉ �D�J�e������|1�R�E��q����&n�&����	� ��	���M,�P`[��b�,�d^�e�!�$^7i~f��X��P�`aE�ZyL�͓�&1RȽ�w�MIZ&���[A�O��|5	,�����)^� s[[ۜ�/NsB�&6?�m��d�O����8זԢc2�=�4N�ӈo�y��YWm�Crn��4d�I|O��Ɔ���XӚ"�'�}:<<�����[�ݽ&����|U�n�����o��S�Fo�*���?R�q"�f$���_!�F�/�_�Q$GH�yQ7�O�!E��P�T;��Qd]�}�Nk!�������q�vw봼Z�J5Ϯ����Tߵ�=E�YzsH�~xM�o��?1V|W���z!Y<�w�${z���`y7���BQ��(~Y��T\^�{s��2IF��-e�ǵ�@~q����k�Y��`����#�M�U�D�YSo*�b�ǩ�kBƀ��H��$���yb�-����5H��&1�	&I��0)�u�웶�$n��&�߳�zH;�X�ۈ�K�V� r;��.���5�{JXn) ��p�@��� 1�]j�:Ԭ7���.��7V,�����T\M������uB��ɒQ�N>`Aw������z��R�wpB�b�rW{D]�W�?�B�[=j7:�P��Wbae�����[p{�!� �s	�/b�a�\T$dP����rAR:$X�T�Nk�L�٘�T�B�	�#ܾa������ c�p?�  ��q8�E�D�kk��Lv��ګ<�U� ���\/��k�d3�O�aIhy"=.,����5��N�_F�|^�ud��e���}������c��6�g��<��s�e����h(a�͛���wyW�-���yN��+8�D��}�n���`E���9�b�JhXգ��X`�Ƴ%^-.�iaٝO�mʝ4U��#xJ��LwQQm�T���C����=8R�Y	�Nv���ɚ�	0\|���j�Z����;IZ��a)��X ^#dp�Hr��5]n��-�mXz�d��R�����>��s"ȹ*�/��u!�L^�<в����C	���u��eQ�o�g��s�kz����vK�-,,��]"�.UI���,/[H��d��Fww����l�_&FR�&
5h+[w��aM�B��|A��v;��T�D��ñ�A��Ll�5��4�W�Ĳ��m1mI7��j�IW�V:���qC��s�w�����+B��S�G��Æ�Cm�a�bA��"�~W�at
��^�K�g��@f���7qi;$���O�	�<���Ʈ� ˰�#����M39SR�*�Lf<0ڏ�I ��$�"M�n�g��"�g{{�I?0�Y[[���I7뫞��K�`޳�p�$y�I�q��'>��{(��~��Σ��� ��c�%umYך%wYlaaq'0�iV;L$ݻ&9�uYW�|�y�q�}�ݏ�i����_��hB�."�.� m=t8����ؕ�yvcV�r(���8�0E���T�}j�<;gۓ�N���t=F�F�0J�F]�:������؎��8�U�� ��G�P�{����3���I0�#��@o��\Ga�Dr',��"�!���sIX����u � � ΀$�������uåȗd��'U�]Zr_H	$\7ܦA���Ʉ������q����.�H.��Es�)������VR��Uu�������Na�qL�y�뼎aʃa�ֱ��J0�2G_�	/j�B�@�P�6�C@�":�"ʆ�J����:y&K��!�A��%IE��HM�-��-&Ǩ��j�I��J2vVV}%����!u?��(��E�3�T�6�-ܡ�9�_��u�_���2���	�gXqA�|��S���%X,����c�� 6:i��f�b!��H�/X|A\�n �D�'!��<R! ��@��{��a86��I=y��V����1��6�{=��/~����Oc���`(e=7N�	�1�V2=�ܶ͑����-�����dY~'(�������^Ƶ�Z0��{ϋ� Jp���Zq}��'���2i&N#Ѡ��Q��U��*B��M�	c���0�'��8���U߉L�,��*�]Եn"�b����k~d#�+���8p}� �=���	��5o�D~KC1;���̀�ͭèP�.e�`�р�N_I%��������*f�b��B��|�ii�"E��hZ����䔎�����>�&�tK���,$M�I�Z}��L�vww�ހxIR0��c7�oY���(/%J�A�csNֿ���w�Jx�|��-���a`����_�� [XXX\�B0�Ƅ<��[���Ÿ���4b�.�\��љ��)X|g����u4)������ͽp�#W���Z������L��9L���C�U�?�X����^g�v��w� {z�/ٴ���� p�y��Y��t�vD�H/�ݥH�e��fE��Q�p>[��bR�A_!bƿb���N�����pZܧXDA����H0H,��$Q�!	��B*�賕��2��_�:���o^3q�Z��:�t�d]�8�ǒ��c�a��5A��m�ݻ�Ǔ��Ik�m�0�&�w��{�o��o�|qc���wr��<
d|�"d�7��M���Td��Ӕ2iפ����������
pn�7a�u+�^����D���e��ڬ���ԍ�>S�����^tL���Ǝ!D� �};XU7��ۗ�Y$�@�����a�,�BR�*&����G���X�=GȀ���D� �ޜ�
���$V7�ʨ�D@}7TύK.n�~�C�([��X�����У�#& ��I�[q��Jz$c���H-] �d�was_��^Ƴe���K�����$k5�}%�����7�iK�q���A����^�w������e|b�a~��W���B���/��ĕ'c��6��R�����ٳA�1�6S��o,����S���5�B�$���p}7��.�"�%�眈X�ni�7'�S$l;�۳�-z|j��B�c�A�n	�Y�	���P"�i�-�N�
�a��7pm�ub���w��Xz�-���p��=�=���{�y�Aj!_ /�K.��}��0ݎa)�g@H��c ۍ;��/gC.�L�/١�R*5Y�ڬfl�y`�_��������(�@�^��U�"%�;�:�+	�p� �8&>/;Ǭb���ץmg�T(�_�o ���}ܗ�,��k�gI�&{d���j��v:@��b��k��%�1�w獹���;7���7��nF	biq[�˙!Y�j!!8V��[�����ˬI���(�xׅY�N�/��B��*ǿn����"#��-�y��Hh�+:���%MȈ����?�.IjŅp�Z�� �P��J$-����%\�ay�����$J'�"��������D�*�B��M�}��Z������2[��8�$�y�qϐ}�e�ngg�	�8�/~7;��F)�gF��ߍ�1�AQ�Q������(��/}e`�-}�ɲ��@_`|�_����#�r,�������!�Ҁ�x+|7���^�@��Y����}�a�3rD6	�X>��r������å��!�u�DX@�ś``K���eC,c��;���;0H��+�S9rR���[����
,�B�/�%،%˯i��x	�F��;_����d��ظ^\�k��S��T(H[�,�&1L.i�i�JZ��>A��
T?BQ�E��L��կ�ѣGL�)�ח��[}Ŝ�w$����M����	���Hk�y�%��i�^��}ʹlB`� �����$�����!���sb����a
�l�c��a����1�`ȉmڤ����<���Ӽ��y�HX%����a�3�;0H0�EA��zL��$�3!��>Ǚ��c�T�Kb4�^�ey�$�W%�Vn�Wb���wqq�Jꚛ�f�g˸���P*�����>N,�܋q��7	Y�=cVc� )��?�����K����J�4 �5ݦ�r[���T�Թl�K�-,,,���~]HӼߖ�%��_�&���-���ǏYx���kOb/�R8����,�������p�c������g�#��.���I@�%Ȗ.�Ą�q,	�*���I�4�7K���̍JV%�Հ��7��hkkS��9v��9��`�ɔ$�V� MY)���;�ї_p��{m�(�M�_��W�8�m�'Ex��d�;�7X론@��������>��C�jXqя�C����.�a`L� ����[��C�u��s�,����0'�8Ki��G&�ih9_�JQ�^�)HL�q5��&�qڑ��,���]�P����6`�-���x� ��3h�>9���d���}5���42���qp�k<���,�B���_�����B�eC�B=�
ɯ v�=<d��N�k��Q-�O�U�3�k4�0�����oK9�52.!�Ūb#�~��YD�SP��&9�&ے6I;p�G�s��x����d{���1��p86�.�/�+f�=�,���&d|J21(�>��3V�~��'�w���o��bd���?��O��7ߜI�(��P�`�aLz�k��`�[L�����Dт_f������ �n�{��uRA��$��0�Jbd
9öK;�e@�\O�]�}�Y��Р����)�̙�Ģ#�Ô��m��Y7Y�8�OpV^��˃u��$G����Z� �����jq-֣�øL��xS� ����<�+�,!�x�A@0 3sr�s�M#�b�y�ҊOXB�l�X/
7�6�$]�@G����9�G=b)uR�$�1s\Ɯ.��$
E����R�'k��Tɐu�7�Be�����G��O�c�_��_� ?}��6G�������c; ���7)�4g�:';F�`�[������/N�Y¦E�/��6��d�4'P�8�D�Ap#:�x���9�C`�.����6Y�L���*Z�0� 'a	��0���(��g�b|�Y���y圃�U�7�	B.N�%�X�`���j�Sd]N��Xc��@�q1ρLH&�4ϠqHbRqhBb2AA@��
H�d�B�(Q�J[�D|��'�=>���+�����ƹA�d۬p�� mٕ�*�1>��<���ӐTH΂��E �vpO���_�`�K�C����oNd���K�Z|��A��)n��2۬bp������V /G!�p��D	�"�ъO����,L���ɑE�s�"�&����fq�L9��0M�	T��H2�ۈ�=��q�b������D5����ǽ-�$����>[�o�G��N��H���V��GO��	�љ��T[\6�P�=_�H��ȯ��|�F=���Wb;1���s��B%��9^L�d�UZ��S,���
�UV�[_L�4ڏym1��\��p��/����������������wϞ=���f�g�7C�̸s�%2���B�$�y�����`�[�d� �}��_�Bg!���	ׄ���H��ysH�( t`�ֆQ�w�˞��
����^wyֵ�Ũ֦�)�+��EL�	�X��x���u`��.�F�b�b�	p�O���gϛe��[
��g��
���J����x�$Dq���-�A��/���|�yB2�� 62� �r�m`��wq+N{%�0�k�jR�c�z��=/�7���<0���ޚ%���S0f�y���������k�;����x�8n�S��l��5�w���I�rK�%�wx	b}��9��΃� �@R!�`��	t��X��Z���
��wh����I�!�`��0iǿmVaS����1gDq�#^g�hjaW�̸g��Ҭ�����f�3ޒʈ���atv�887�]MV�;��A4�p�X^����ea{�>K(�OW��M
����a�iۊ�R�v@(�.р�mB�,H"��8��c�"$��d�/���E
�I����B�-�\w��S���9�M퓜"���r;t3极g:���~�Cqg��XI�駟�Ç9Xb�Y���׌���fޖ�;���ya	���ŭ�$�0-��btqJ��D,���0��`&�I&z��d9��cda��<�{p1�@ۣ[ֿ��ǌ�2�����l�X�)	�(&<gy�1,�&-��i��翏�'�.��@�Eq�X\�O�Su��}�Hh���6�E���G�}fƟ��D��w�3�������/e�@���v�ϡ�?e���Q2���	$a��K�+��U2�K�!l���X�����!m�[@�G�21�s�y\�%~r�1�b���1����y*0f������B-F3?�8��Z�-,,�,�/��`q��S��2,���#ߓ	5�`N$f�ͬY���oo"�A�ɪb)�"'�W��iirԷ�Q��0�[���r&���4?�:2�"S���=���,��,���A��� !\Y�� ��Hcb���1�_S��Ǧ�gsD��m���M6"%�x��{�� }�H�[q^9���-Dgww�?Q'X\a���Lђ�_|��8,� NB�d޺��;�_Lu!�漒�cL��w"ݍ�!�}�x_�=�������\)�,P�K�4�W�f�����e1 ��'缷� [XX���0���YOu�^{�B��	����� �Q`�'Y�a��`��6��|[�j�@�!�\X��}�j"��4����H�W!����|Z�_�h���)��'�L�}.s������S��ef�_�y-��#���~�;b�&ۨ7��j*��d��0�~���b,8�b�k� ���8�u���5Xm��$/�6=�YJ��x/���Vd�D�y]�_S�*1���ĻA�!�{�V/��]<�ĕ[��4I�+,8,�R���Š��Zg�n5uL�;��5��A�T,\��>y��<�C ,��?��yZ[_����g��R'}����-�W,�R�B*�*%I���y��`�[��L�Ү}}1�q�p�kېS\��b&�H�q��"�ȧh�e9��פ��U�q�}��g	&a	��&��g+p��������[�xOׅ�%I?�]Pu-��w�o��cY[���B���igg�c�vvvXs/�!@Y�gK�E��8dc�
���=ƵOz�X��{���������[%��+�a(ѷ �.$�rB�������3n�ߡ��b�/��N+P���.����`3����'��e�͊�1,�b�5ߥ����I���|J�d]@02�Ģ�bѕv�� CX0f�.�g���]����K�=�XS,��!;�=M#i�����O����7���?�o�K������/����?�����JEMQA�,��S�!�
Y��������� ¦�'M�8p?�A��	K�-,,n�K"1�U�	��q���b�Il�ۥ��N���_�P��
���'���He)z�Ȳ�-l ���<G	��x1����Q��J���1�sen��|���W�W�����HS��Źf�~�	�i�8�h:�9�~�3a�y�QrD��,�� �]�]iLd��U�Ǚc�0/�Ͱ��57���ﮐ�0ryNy��1���Ϧ��1w�e���ǅ~�w�$�plXyQ� ��$H2;�w)g˞$E�E�@�d��dh\��e�� �x�{�Z���~�j+pֺqϛ��I2q�$��`�G~�嗴y@"���sX�Ņ��kl#�І�s}��v�K(�7K�-,,,��j|�a
$7��k"�mp4À��w1Xu�	}[$��K�D=��)�Y~}�L�AD�u&�p @;F8F��Y��'O�����s�Њ��P��K�u�ǵ�
	�
��,Y�&���b2�<���K��؆B���{��;o�:��>��r	�T`��j���̷ ���x��0to�;�b�XDc���� ��V#6X�7#�q"��L�e*r�A~e|��]�ö���x�ɺ��}�	F�����Ax�[ʷbQǈK�e����a�+%�����8������c!!-n���a`b�_d��I�4�k���cE�AFx3%���z�1��EI9�.�@vss�8{��κnuR�$�M����L7h!�p)��DD2�j!���R�K$��(F���x!���Hc���x����b�q$|F
�~������Ըum���'��9���t	��kȌ�n�%Z,����@~A|�
�M�x�"�B����!5�+E�t[0����]�"^���������k�dX�%���-����!d9�I����H◄%��
���0������zlY�u}���AVzj=,~�H莄6! ¨��Uۄc;p|N���9T(إl��;�-����ѷ�~K7E�0m��ybzǅX�`�EX����&nd7]����e,��Tq����d�W'Z�<	���(�sH:��� �j`�jL���� ;�[tp-�g��RW�YC��BaK0�x�> ~���ĂA92�#V�$��U�gLr+$L,�W�a{V�vߓ�?+�뤞3`Zq�]_��kHB�L���mzo�x��́"���!�7� [XXXXX�0�,8��	0�o.��T.�9�#��1�p�Ip�)�{jQ�8P�H�*���L�(�ol ��u���	L���"�����d�g���4Am��j�w���g�S��a6Rv�PHR�H,Y��F�_X}5�\�W�>{�8C��"6p{��~O�N�Eݎcݐ��]�x�Zq\y��3����zv�$�RfO�|Bd����$㻉iY~�m�J�5�1F�~����dn�~[XX�Օ��(��>ˊ��-� ���Xɱq�1b	��������B2�J""�cE~*��(bR*Run��T)����F�Z��kM:>:a���I�Z�@����Q-'4l����E�[#�� Jr��\�X�<��6��1�]4;m���i�_����B���/B�%�D�Y�]�bG��N-�d}��/���-.�q��iw��l���)�*rszܠV��׊���:���&¤V�i�,ERֳ%�<��	�����X�:���,�¦�q�u�:�Ѽ&I�'�Mi˰<iǺ-�~�X��W��ol��/�Kz���8�[�7�{���1��?�@���o8��_���̨Xlaaaaa1#/��I�e��H�+�V��󴲲LK�UZP�dii�V���
��6m:>����<�����ϖ"ŧ�T�Xɡ�4���*,V�(Rd�6l�jyFnh�&�\ZF��8��q�Өui�ӴFO�l�c
����oa���}����ha��{9�3��;_=*�ha	
��OyZ^�н{+��2O%NZC�V�Vk��uJj�6�����:��m���Q$�]�%^�;>���s1n<�Y��\?$�syH�_X|At��Q�X�w�.��b}�#)im�+�$HZ*�}׌97ݝ=��MZte�[;�0>��g�������3ʃ����wI4�7����C���ի8�e�`���D�!�A ���#�"���]�O?z@�o��ڒ"(sT�+*��J�	l��Rm&�''���0q@�~��޾�%:�S����8L���4S$��y�đR���FBb��w��(��4c��,�Ib�w��,QRҵP,��1"!��兂ER�-<W�1ENrn��_���}��z�p�6���*�|�@e_o�j�t贆L�uz�{J��������C:�?UD��c�%�p�<+ҧ��)�"y�s������,Y��^��w�����ﳕX6r]�IZj.�|'�m&���s�}J5���<�e���ӂ�,Ͽ�կ�Tj�B�k.\�2n��n��"6�ѣG��g�Q�T�~����ʊ(U.�
l	�������a�u.��D�o�챛���"&k�ӟ>��W�`Yf�[,zTȻ�Ϲl��G	�yE�+�l�J(i}uQ	9�}�^�+�rH��Om?�$�8
]�lYb�K�?"$J�'���W8<��8�}�:��>h~?Ld+ͼ)��3b�c�T�)�[���9z�p��ⳇ�����U�Zɑ��� ���c#s�����Q�����%�ؘ�ťU(���;u�CE���K-��$x�x,KHD�"�B��ViZ���j���"�:#9ǌ+"��X � �(����)y���y�&����)j�k2]yC���3���d���(����~��ܗ(c���_s]r���K��`T �����<�A�	�f��4��n	������Ō@��;\U}�T�.-/U�ɣ-���?��O�hm�L�,qM�;��o���hWi�Eb7G9E���Z������5�����L��S�%)�>:.T'�
�[g��.��шz�Wc�׮�H�+p�(aա�j���_�/>}B?�pK}qɓ�v(�k��a��:��dWuA
j\�Z]�յ���TD�u$�v��R��r�qr,;���-!�6&��O�+�2&�i!�9RR�c�7����Wc�|X	Q�`�R��7��b�,��Kq욫�d.�v~H�$�"�X�� ���"	����?r�������	0�� ���={F��ɖ�O�2�Fp>o�4K�-,,,�0�i�{�܉�5�ۯI�ol�c~������G;��'�������"ݠz�M~�M���,�(�.UO=�Q3b���$Y��\���lw�=j6��kK;7���0�F���F"����Ud��dW ���"<w~���M���{����уe���������pVq���xj�p|_��H4jw٩��C򵞯�r��#&lA�x�n�'�[V�=~=Y��16�H�E��R*�AP@f��V_$�+�j��/��4��j$I��KkZ���f��uɾK�b��� H�w�}G?��#�A����Ĳ`��W����a�y(P@��r.�ò��o,�����c6aX\5�{�|��35I{-�9���D?��1}��{�����S���͠M�Ma��%���(�t���C�n�|ERzy_�.y��L]��Ӈla>>�Q���BvUu��jl�i���
��w�F���:�;Ɨ�L�m�-�Ͼ�����=�i��٣v���ScF�z�)��Km1�v��"Ep;�tZ��r���UZ])җ?��J���o��	��7[�\�b�3��m&j��f��� �pw���X�k ,��e�i�>�>A�Ar@�p��W�_��X,�I�y]�I�qN(u`�L�˺��p���&�L\�1&Ч��w�WQ|ȵ�]��2K�4�(F@��\��IR�:��,�������zJ�&�0����˄Q�m�IBYp)�b9���yE����u���D�R��o�ߛ��v؊w堇}N9�V>��C�]�S7a���T̗9~������K����k@��Ť*g�OcHM;��"������z9Nu�:��|��hkc�~��}�x�*e�:רԨ������ԉ��+�xp����/��(���<�˥*=|��^�|��Q����Z�"�6�R��Q��(�{��䙸�(�d�$:B,/�X�Lʂ���4��O��8p����_'�5	�X5�df�v����;���s�$s���%cQ����މ�Y�J0Ʊl+ߓ�%��41V��ߖ [XXXXX\)�(��3��cnI��	f�e^��h�R�յ��Bɣ�
pCUD�o*�X�@{*�!�[J�h�8O'8�o>�qX�CEP�^�:]��|HKU���J<ݡ�z��s��IT)�L4�;3��Œ�ل$LB����8�)����H[[+���Dˋ괏��Q���J<{�,���u�z5�:QyW�\H����c.T��&g�.�K��Z��>�+�T����n�!��13&�$3�8OR�,�VJ�p�;��q@z�	���>��g&�@pa)�$S���Hc|�8������;��Kb��ܲ�ka�Ji^k�f��t�1ۢ� DA�CI����a�kQ8���Va�i?r���M46S8ͯ�� ��q�m������M��o�ڹo����0	�&����$�S.�����%X�N�(���F����|��9���p�n�񕊸ֺ���P�JX����5���	�W��")y�7��P�~W$(�������
�yB/^(�{��;�l-�z���9BLA$�4�3޳x�s���a�*���"$�o��X*���"�߅9��n�:���\ۜ�9\��j5�T;nQ�4�v����95+syZ^��r�@�_�}¶:6\��4Wqhks�66����{k�o��v�ܕ�X�w(&B�b&ֵ��y��<�	����)�=�o����_����_,� �b��X\`�t�",.���u^��1�c\���x�}4�u���m!�IHb4����B��mƷcA�"�1Π1���C�f� �C��Y�)������$��V�maqa3�Cr��Vdq1���{�?���c�h�P*�@g�E�!E��઼En)��I������� ��F�޾�ӟ�ݥ�ݚ<97�&Z_����tO�iX�9% � +��n��iE����vy���~�8亱ڂ���� 1��I�@��1I�u���;N���%��j�D�n)7��mm�����A�:�,��+�5O-5NN���m�^<;��ݦ"�=�K������&m���Pʫ1D\��B$f��q��|5O�乜�\�P��9���X�+luW��$q� ��N-B6���%�����:ȭi�aY__�Oq�6�}�1�:���G,� <�!E6i\��ں�޹�P�!�,ԓ\g��8�X���Z@Г.�YƵ,���a�Kg��|������_b�eQ�`<w�}Fl����cK6�Ur���]�!�Nc�I��u���"�P��8�%laq�`����Z��B��4�����+8�;*5�/�hii��@�� E�ɘ�\�a���I�����ջSE�O�	�r�[��2U��+穘G�_�%$�Z��啶���{��P�ة:4���wg{K	3���W�X�2�X����ƿMi�������3ﯸnr]ΕU��ڊ		�[�"b
L�wV���{�����F����\F�U�	�O��!��C�۫S���,�jw}�J�*�Jd�(��Ϋ�WrL�+���6G�FȊ��XĢiqҿ�G � �_X_A$@�8��0���i��\ # ���������Rn�o�f`lb_������9p��Z��H�������@ܕq=�>�O�m*�%Y�8��q�ež�/ܻ��=Vf �J����hIo ��������/���������M��=l��94��14f� �Y'L���\o.�^�	��cI�����m�lo$"b�w$���Tԟ��Ď���,�X���L�^���;U�B	�A��1`�a��.��ר:����"��.�c���`��T��Ǐ��W�t��#�0��bHH��mphm}�>��#P d��%�/b-��>��1�%�w������K� �3Ǎs��6�*��[������1�j� 9�B�����<���-j��������iБ"�o�*���J���"�G��K3�R*V9������=�n��Գ�w�a&��U��u�3I0B"
�a.�,��48�<�_����\R�i)Ss�p޻w��``|�ju��ފ��I���;s
��7�1�=�!yύ�Z{�w�"�����7�p�=x��676iggG�QB��(.X�c��>`K0��:�_}��z���pQ%�`�00�X�c<�2	�����Oj��<�F������
�����`sa��P�'{&��r��A����n��fG�_]��^N���w�p�i�%ڜ�(��%�r='JDS�C�.��j��Y��Q�e�6�׸�g����CM��t!ϴ�Bx��T���`Y*�TA�A+���^mn-�bU�f�AAg �OT�U��V��p-t\���l�uCj)RPk����.��ؽI�0�rJF+���`[`Wh(t&u#��H�@`UA���T�>�Y��y7�Y$�ܖA
Ar@D����\�7rǾ(�@bA�9.���:_+�/%��Z�Z�N��&�^�����BRq�v�j������k'Cᶦ�`(��~2]�M�$��I������^�|��� ��`��s���2L����Ƀ�Zk7	�1��0������h�D�$D:y~��ow]p�:�Xsɰ�
�����(v���mơaQ�w_()g��{�j���#E�����o�u(_�S���s���K��R$����l1�0	d��q��&�cd��<��G9��y�=��8q /���y�!;y�ᅰ����I�(��Dq�� C�-'*��z"�r>�������Ȼ⪛̧c���{?+�����25H�X~A~777����t5���r-���Qg�	��qr%cߋ�T	o`�n��&d�*p��a����w������=zD���g��H������^�xA����I��=���4N��!�$1S0@��~��K�w��%��vۈQ�6B4H n�d���d7Y�baaaqܦ�w��r_ͺ��xԱB'"N?)�Ry�tTJ��-p|o��{:�Xm[ȫ��t� .y�
�SD���(��G�߼WBnKq̱�y��/�ԩXB}NE��3q\�Y�C��9΅i��jϸ�K8�$0=Q�+�ׯU���!�����7���95~�2Q�iY�	0\���Z[V�1�b7�"�*���j}�Z�J��5���l�����o��Xծ�Q�����=4I?�� i/�E�5%���f�5�=A��X\��ŻD,�8�X�/�$Yk �s�oi��|�.	�.:~�H%�׸��Sk��;����p���]�q��&NZ���������G�8���9l�N\�mB��$˜dyX�)��2,�0@;!����"܂����,,,,,,F#�;��ƾʘ0�y�	��J�@V�Օ*�O�tz�$n�=��cK����Y���e�S$��!ы�r9(q�S�qJ�?ۣ_�������&?�r��;�����Gmnm�Ww�b8q�.@R��ߌ�'凫�W�����۷oY�����%�"ŀQ�W�~�woU��O���:�-T�[��<��7��V�55���j"Cn��J��Ksml,("��Hr�ݝ��-q��*j|����Pܤ�ú��N	�'-�ȫ����@J�H6hȽ X��$4�t��:n��j��[|�b�Y�)1�BXL��eXb���z �K�*��ݻwl���ގ�b�{ܬ6�m�/H�%�bt��s�����+���?�!�@�7oZ���q �%�=��6�����[V�]N{�g���p�;����f�/�G&��@`�M��m��K�q��Ջ������$�c���oh�u;M����2��v�����
������w�	ޥ��zƢ��4�^kRo>ON��V��a+\����b�����n�h��q�^�X�������"�sT(���
f@�����o9�؜қ������o���4��F{����!5�y�851gax�����"�����*!��?}��=ףb����*!�I��񱜣��Oy5��B�-^p�^^�Pk��ĵ\*R�𵔋m�q��V��j��5*e��������F�N�m�	CDW���ȁV����$i��dr,dhȹI�`"�kG�5c4�lJ]^��Y�8�eX~�ז�Y'��b	�uR'8��%ϑ$��D�%��G�9I����Y��,w%�	�
�q!���ًq������S�?iD�l�8�fN6ά%�h��]B�4��������7>�R
7G4Q�y �8�b!���*mln�f�������z��v�v���8��Ȱ�q̌vL7�b��6?�׉�Wi�]���A�h'�%Z�}���i���"2�\^#��S�U���%�̻�G}_%�V�Z;�2���� W�eZ^*���Ժ.�x��{*_�b�Ljs:>m��Q��h�~.
B�<´�U�8��x.�\��V	+b	�K�Th�N#-�.1��:��,��9���NP�#El%W����Rcc��\ZQ�H�<n��'��,���
5��xv��A.�"�r�܊PwC�c�I��^PPcʥZJ�� �Z����N��b4D�Ƴ�K(�!dc��0�@�q ��f����"�˼$��ߐ��)	���Z���fV��I�#�o�Z��A�Ԕ=U��q@Z�p�R'X�M~�*�q=�,��u6mO�Z�s5��9Ic��Vf�_�̱4��w��E#.������'��wx����1˚��7j&� - �VT<\|fAmh$���S�$���^\��.� ��_�ܨ�;\.�#�C⏲�}���8��F{���j�8��y_ҳ2���a'��B��.��ىNɿxWs��]�X)ғ{�2?��+0yI��HHp��P��s^&=^���J9���:˴A�+(R���޼=���t��Ȓ���9`�.s�V�	⦅dV��&��!-Lj��z��"l�A��
\�?�і�0j��������3��I�/�����R1���B�����c���ڑ����1�ƕ�����h*b��X���\Ǔ[B�q�V�!aI��\X�`�Y8��ɌN�[s<��@Ɩ:����ʌO3�3͚z��k¬�"�����VX��$��z&���{��"S�)oS��X9C��gD��$-�I�հ���ыj:����@����K�n_�5�l��<�� '�/2qQ �O�<�Se���'��� ��j~LԒ�J�:K��E��EK�1 �bZ� ��޾��}��!��9^�~Iϟ?�g�~P/��h�֢�K���[XXXXX�')�D��N�d7�%���yɡ��}|�6�(��K��kr�+$��r� T.�dHO�.gwF�_.���|����:D{u���oԼ�ڞ'$�Z��q�q����!Iܳ�t/]q�b�Jh_@]D�*�����z�
��E����J����P�Q��%O�ٜ��E�C�����!�m=?T7��Y^�D�7������w~E���R�XgX�1��y���i�Y��� �
Y���+�$��2�)��2�n�� � � "���*cܥ��&!��.�Qg�A��&��X��^�#%9��g�Ϳ�8������}�H�%۲-[�,Ŏ����f�!p��I�c'�ĉ�ؒ-k#)����}f����q��=0 f���p���U��U��+B�/�c�&t����>*Te%�+����[�������m��?�����jרt  �j���B��e�=������DfB~�h��\�ef<�&�7���0�����FN�<i�^4s�P��p!N����g�1�9f:'O�
�Ã�e�we�6�L@���a���
��PCGYhЃ�����Z�#�ǖ��}���p��;��;.^8�ϟ"�F����Y��V���h�H��*R#Ͷ̌�����l�}o1|�����wí[w⽺�5]�%�`x�^N��� m�ג�R_U=C\|`�����<h�:����f�s��ͯ���N�����u2��0��oul^��|F��JC��D����d��E�5:�o͇{�V��qn���V��	�q.'9��<����4��nġ�8� �Uuy���H��~� @E{��a����ߐ$)X�"B�R�_]�%~��׀CG���Jp��oj0�oU��؎C�͜�t�=�	sܧ��}��O<�A����|�IK�~�@��� �ҧ�P�l�`%�>���Uh{[��t��%���]��������R�v��K�.��/^�/_OǶ}�����hI�777�f�	�L�������PCqʴ�4���Q���*f�춳<�Q���"S�	7o/�?�wݴ�?�����K�Ck.2�հ�Y�=���ʍKMc7c�� ���E@ȅ��։�tg9�����,|��RX|@T�Pj�s#Y����	�A��*S�*�B���t�|��00C���\괻a)ί�̇�o�����{�é�($�E`�/_��(��bs,Gǹ���:��?�T��;�^W�|�اᛯ���[���7���T��̠e�0 �=��3�� L�[ZOo1��7|6�7��F,<>K�S��\|� ��*�b�I{� w�0}Sz��'ԛ�>��o4�(��gY�j��9�t6P�9�wѳ�P&ؤ��=� 2P����_̞ya����љoۑ>�_u��,l3n9�Բ,_��l@�H$��g�?u�����{p�7m0!��/c��ݽ�������_�F�PC��*��aiz������aֶb� �M��i�K���,.ŉ��-Uͅs����)�E��@�ެ��{�X��Ό��v�N��YX�Lo�w��"\�䛰x%ln��}�S��vK�N8� ��0�e��v(���p�ݲ�Gh�-�tw�Kq~}z�f��sfnv!l�_
��]'����x.d3��8wL�lP�&�d.γ����Z
�?�>��p��7��"��sKD����a�K
�����>�������	�oi~��{��"����J[�>��?[��ﬀ,8@��c�[�S%x> ���/VC�<ȾKQ����W��h��1arp�N��7ߴ��	H�~�3������U�#	nn�{�ws��"H��"f:����{cc+<�,���f\��[{^~����'�k��jR����6ܿww��٫|�-b��A-v���dn�rC�R�.�a�B&�>�p��v���X� �]$���"����_O=y6���3�m�~5~Z�_�E4ޭ��G�0~6vb��GW>]�:|tW#��,bt�������kއ!W�I�x��c���)��,�7���֦=K%�g�g#�R_~y'��l���/=~�ʷ��^�@(ί��7g��C��n�_�I���`=�q��'���D0��8�n/���u�?�	��-ea�ߣ���	6k�`Q"��l�7�MeE�<`Ds
���|iG���0��c�/��>�% �WF�+0�GFP%>
����w�*�� Y�.S���ԛ�ˇ]�����
,��ms,^�B;k�"�kѝ�h&�HY���7�'l��歛q!����۬@:H[f�l�<��iJf Ya�D�[���|�B(�&qׄ�����o��Շ��͛� ��<��ַ���S�^�w½�wM��94m�&fѓ�9z�qƛ��� ���H�Xc�`��$*[5�� m�u@U���ԙ��;?Ȝ�����:��oc��A�nh��e�AP?����2�T����<]v�΃�a�>�]�uݭkJV�>c��i�r�E^�$ ��f���%��q�̄��#�w
M�l8v|����LCf�fum+,?\7����_�
W�~>��V���aq)2�E���e��~���v�/�\����_s�g�z��G��V \���=��s���(�jNvh��@W�&���sp�K��Z�6��φ��ZZވ@�L8s�X�[���\0~.3��mJ����~W"�>��v��ӯ�ܺ�-��c=lls+�7=�l[�t����d�}�-�)�s~L|�O��k!|6�� ����oV�#���k?����T>�u�>��R�Nc h���] ���. .�v1}�����]����S�;����v��x�q�����*W��|?�|���˥�r�Mc���Z��\�@d�̣z=�x�RJ�����g���,���f����^E�87˄nY�^�:�i�0sn�Oa������Ʀ�E[gnbV�L��SL���ݻ�B�z-���xy.Y8��-�;o���ջ����N���L��A�h�W�<�[�슠�r��M��B�f)!���������U/D��J�|��T2�ϧ�"m�����SO�=À��6#zT��7R4��`kG��Uh�fa/>N�lp�AUfj����(�9R}\�T�5�`)*-�����6`����㏝O\:�p&��p:�<q<�n�E������_
�n�_}}'ܻA��e[��ڙ��.fCVX[Y,A�\���
��U�1l�΋�����l�2�d��y���1ﴏ�@1�s���L������ u)Ι_|D@������8�;.<N@�q~aR�5kue-�[��+���oE�`р��j��o�5�-ow%\�	$��f��7�/|�3����o���\�l���sJ	
o��K/��?��Oe:#i�8�`Ww�Љ�f� @��z�	T�t8(�Z�zO�t�	�E)ȼ1c���1����mJ.��x���zg[����P� ��q�]ū���W����5����0/ Ί��OX�N�ꙧ��/��~�i�p��y���O�~��7f�\2_
 ��M�%�Y8�����s̃c�ܽ��s�`�ba��i�����}�7�G�xkc}���nw��̄��s�ҩ�֖�/����p��-����Vv]��CT��M~"
 |������^t��h��ۃC���2,$W�^5�^���'��9�OО[�;��Ӥ��Jy%	gzO�K��B/)��~rήۓ`�����S}���KDU�d�I���?�~/uC�!/��������ԯͣ����Ԟ��0���h�9꧁�v��雛��Q����m���k��nG��T�������3��Ӗ�`.�H���m5(��=���x� "Y��`D����JOW��,��}9T�u;�6��n>U	,��~�� �����$ �/J��U^\<�PFa.�Ұ�-�!�X]��եp�n	wN�on/����s�φ�'O���WW#�X6��͛q~�[ҝ����B��w����j�F�'��9*n@��B0,̠����W�Ay�Ѡ��B�P�g�G�>�E���p ��8���}�׃���71�P���+�_U���W�6��q���@c��0����;�D��Jp9��� �&����$,R)�`�A>'�K1��������/��",.=�/f�r��K�s߆�]�@Ul�D� ˼�o�yf 8�H݈�w-� ERp���(N��7-�9���9�|_��6��ǟ|b/��(�x\�|�ڋt����6!,�^)�C�$��o��f��믛F^9�<��d��c��
Hخ\�R�<k^�
��	<'f���9�T�EJ��=%��T�6�}�`�8�~2�Z�;ux���S!��cn��瓦^6�J��FBy�=IS�_m�� A`^�h@������b:�Z_Ou*���8�U5�x9�T�<�֏y�24B�&bs���n��a`���{�m���,��ҶeJ�oD��~�US�;�Z�h
�g��.2b�/�L	�\j/�E`/��������:�� ��<�T�0�����U��\�ϫG�GϏԪ����j���N�i��[(���V؊{"s̔��[ox����X v���������z�g�r�i�����[��=7)��Q�C?�v�_J�TP�h~q�d��(z{�σ`�*��T�`�3��$�:</>j��X�@c� g��7�(s�s�ԉ����6� `W>�(|���᫯��<��b�,;��63��df�l+!���N� x�������|�(i[��M��[�6�WVV-���&".-/��+k�<(VfZk�w �7��2��z�����K�L��g7L����oF��[�J����Dl��/�X���{@�"�7c����&�ȞM�L\ӐGpKY���'s@����S6iQ-�Wl��Q �X
Pοt�C�0܁9��,����:$~��?�>�D�Ky�ܴ�z�xp��|����Q���F�c�h \��ohHsD �g'�>C�ڮ���?�h�<�@�wH��Q��e]2M���3TMQ��ud�c��-�Y���xd�vx��N�i���]��-�+d.�5��3oqQG�}��ѮWQ?06l�άq@w���Az�0�|���w�M�4�)����N���v[����ʅÞ)���^ssEBC�Gz��sȲ���5�7�v,�>������QH���p��N��������0F��ڝv8
��n��b*��U블��#W�qh�@j܏g�F^Ѹu_/��pGy~c� ���R����h`�d�����k�ڵ�|.[ٙ"�\ml��R�f^��1����bN��o�`�r��*��T�)�(effrS��t�J'\�x��un߾nߺ���M|!r��.0��Ͳ��V4�Hӟy����<�ͅp6����C�0[p�ܮlb_ ��" x��J��c��� RQ�5�50��Nc!�����ήa����o�9~kRS�/�0p�DNZ^�5���P?��a�0E,Z�����ߜ7K�X?�����O-���}S���k�Y{x!�˃���n������:8���1�fE7bY����|�S>�W�����M�v�G"R��CU�4���I_��w=�)���on��Ih������&�N��c�������O�oC�k���h�)�M�spa��ҵB����:͞��[l��J���m��xغ�O�� ����q;�$�Pp/�7\�؟>��S�?[��H3o���9�����0>���%Y��;$X-�l��
a'{�x�����cG�~}�v��c� ��������˗V���=�3��;L�����p�	4{��.���s��Ħ�}��Q�����ݤ|�kP�>�����������icn3r3NB�c6l����'�� 4�"�w���8��"sv2;]2������ڝNaz]��z&�Y���ge�`@-u�O̢ݎ�����F�6	�댜vk��ob;NG��N�EM���<�8��3v����D�K�v��Ab��9TN��*?�9ƳZ��^~	���}�w�z`0$E�D�x����_�gO=r�)�,  �s��x��a�x���B\�K�<���7�e ; �K]������m@E�}�~�����N�
6!����gl�S��?-��i'Ϝ�x�<'��-��@��9,/Id����7/���.p-���G����O�d́�iT�a���֝ӷ���꯺J��`�c-C�"�&sQ�	���z�

�ۭ;�t��� a=�ӬW 1��c�����K�J �2�ψ6j� %H���d�W��＄��2�,��Uħ(:tZ�4RU@ZxW�Ci~�?���^�p�|��W���a�jG��s𬠹�Y���4�T?+<`�a�~9O�l\�!䀪���1�.H/@��x��'��[�M�he
�L��y���4\�� � /�^����lnfS �`�Yf�x��/g��f8n���*3��fz~nޮ9�p,������Ր�5�L�e��
�ߛ$׾>�q=����3Ϛ���E�-�H��?�J��� X���䅏JȒf��2i���0H�p�a���{�g���m �/��X��C��\a�N,ܴU��f�^��p )/=�x�(K{�����o�mL��˗�-��Ch;/RC�Q�+��ғ\]>3��Ht��zE��X��#�sH��h�F�y7���F}���a�pz�xGٸdꤼ��0A��1<����(h_�;�z
tE�W*��9��:>�s�+���k�����Z�Z[��y�$�����HמR����s��`����:%�@��>����}i/�o���:.y(i� �Q'��� �V�+�37X���+5��l��q���\�ۮ�κ_��V����n~g��P��~����C��&�[��7��t�P�� �Ax�ŧk�z��q��X��N�?�`f�>�d8~�x�����0�
?�e��%��S��sy�'���[�h��!ڧ�4���4<GFmn��ooT��yV+���jmkO�]�Ў��W��IE �N0� ^^~A��f�~-�td)�Gr�=}ټ�(��ؓ/Q*��z�#�N&�&�E�^��@P�Lm4�"�q��k6T$vj38/ĺi��\+8�|=������Jgڤd�2����d�@}��|�r�M"uh<d����i���
���?����475���y6X L�85_����,xEZe��0-�s�u�û�toiZ�i�a��M��ܕu��n4U_iO6Xk۝�jj|�~&ƻ���5���~!	�������xv�?����?4t T�i��}6YBqL��	�I|���f�Ӗ�Y�T��k�����#�`�g���J*����Q���Wh.��A�r)]$cN�/s�D1�Y�y�!M0�:���>0^�í��F�1k��Ν���`Kh~���,�_E ��%y�A�f�E |.~Κf@�'�[�G�6��"B�̭fH�4Wh�
 I����8��Q��S��c��>�ԁ����R| [��-��_g3saye5\�q��	3��\����b���>A@&���ib���:n���z;5� ���;Tņ��?�X1��G��~`��,F�C(�K#Se$��##�c\�	6�aQ�)�fZ��^=m�JU�L��1i���* L�d.$�k懂gq^J�@�L(�6�����O]����Ґ���M1�֏����:R��(`zRH5Y���^�})5���Y��s��K�AY�@�H��9����� �~�n�W+�{�ظ��k?��|N�����w�j�y���%K5bx4��B��QPQ����*?pOi[��DJ���<�q���7��>B��e����GG}	�J�4�7U��	A�z��+!�^*�=��@��\/J)��(��}{3 �o  s��%^�{q22![ɀ��p�ef�H�,�LЭ"�U�[�Vj��ϔ�V9(s�ϳ����������\s��B{����0��l���a�c����-�<��gN���Ç�a��xlib'ny-�_���Nw�ie)e+�=L���u[T1�(���6N�ۖ��(�H#�� G 0�RGnMp���>��t����r�OQ�4�-��J[+4�� *%u(0��G��	�4���@m�]��H�b���nۆF��)�M�(�^�j5� XmN%��"`��3*���q�6�uRLB�����1���9_`GCCC�Ǫ"�/$P"�gx |C���~�W?Sw�ai�{���[�g§�o����*�*��n�\G�(����#V�XL��q�W���H�YQ���s+}��<�*hX+��G�����!<��c�����r��$���<~�I�*c��v8ؠ)�sKf�YV���f��G�*�eE���ϵ�Pk&7�6�!>������{�y5�ݭ��<�fƴ�D9\]yA�M��⥋��o�'�Ҥ���zmI��\_n��u��K�B���?ڷ4��/_�2H�X���b��v�k�Xl��ř�Ma��y�-i�� \H���	@S�R�r�ׅZnA�r�u���y��H�8/9�Ѵ���u�.�����8l(��vG{5��F�k_���y7�5�o�Y��Y��4�Б�AJ��C|�Dk�xT�G	�4C�+�n�Yo���5=o�q|}0�-��O���OYG�O�B�J@;jF�à�{(�\��/�SY��� m:o� �W��6��K��Ҷ�y!�˄��w��g�@6�j,�Q|�H[��(�&<������0.A�>�K������c��V��L{W���Uڛ�je�uu-�_K��K �	/a�q���Mo�&��� Шh˘C���[)��HR^Q���k�<a�Sc�(0�����q_ +�����Hϖ�M˱���`+77k����	#�PdA>��V��A�4��ӴHP'���j���U����<�+Ja��o$>J)i|����zh/�H)U"�TQ�/����R�(�
� ���cT��]�!�8�:����4�S�@p�z#�g��B���j��'��_ק׌Jc�2C���d���ɋ$ `��Ec&���L��DD���Uٶ�A	�J�OܪUh|�- �(���bȊz<�e���i�	��py� �R �� �`[���A���E�����Y{��7 xsC��&�<0էg����	�����M'�'�P��?W�j��V����d���M���`9�v���_�vb�B]��gnm��Nԭh� X}+b��!h~+�5�����p����b&��g���iX� �n��r�WG�
�_#-�H��eP�PC�4��7�PC�K�T�"�;��Z((��- I>�����U`j?j��4Z���?		�*�$��w4xFx7�鳟4�{���8��tW�i�Z���o� 8D���ʏ2��$|u~�H������@�TG�+�B�V� �=����'������!$���i0�Bl�\l����"�}nݾ���l��HS���F,�;eS�I�
��e5M�K&	����N������^
���G,8�O> T�1�8E��"%Z>),��q���N����=�_��*����jC��s��"�T���k)��5A�8����0:e�i/�)6��4��Mk���	��l&�GK㬍�Y�j��G����5�wjƷ�aH<��^�T|�u����G�[��Ah�:S�T3�R��%K�K� ��%��(Ç�����~��6OyC�i��K�T��돋v�v��hFN�r�N<d��YK�±�'�����S���<�0]o9�c9il�@�*�I�k�	�}Z�
�U>����0��'��~,��I��.���t� O8z+�]�)|���n:�`*u�<�T��5�&�(�4�Kbi�T�!'���)��,L���/�8 �ܟ ,� K�/=~s?]|T� �]:/3cF�D=,~�=�̇{��{qO�}���,s�k1�� ����x��fB�`��eQ�e�����&$��E4<�N����鴑��PCG��i�i��g�>�HR�����@�Fs��^�^���k�P�z����;5e�Fni��盹{<��i+W��L�!�9�Bڍ�M�z��v�lx���*�����Ώ���`|i��H�m�]7,�.�1�	�;��=}�ES6�S(�S2�����u�W�i~�<�Qi���F�n�g�	7��ӧb�N��zcm%��l(r�����X )5ͅ�/G oѣ��Yy�Ю~��e�+�\���L�Yx �\�oI�D2mFbH@-XҌr/́aPu��݌u�B�����4��R酤�[D�ib���y}��"*~�KE�&�V��BȦ��l��,�Ь��j�I��$�W@6��c�K~4͂�PC�C�����R�2�xzf���M�����O��\τV�e�z� t�l�����ǰם����ޔ�Oۗ���.mKU`��R ����m�&��1'�O	'������hh��9�3�(=�,��G�^�/J	�# ��?� ����wXaf�>���(�-���g�4"/�0�P�,^0k?\���6�7x�:�̑}�:+��YSzi� � m�+@Z �^�\�R���{��9{�ڀ̍���կ�*����7�,�W���"t7/g�f���i��l�<�����؇m l1�⢁��M�,�����ؗ�&��.���~�@��XRFA~�LdXL � ?@'��_��	�HG��
T� o4�\C}���Ĕ���E ,��_}���S^9z�.��q�
��*J�A��Q������k̂/_�6Y�ʴp.M8e8���W�W�#Ə1����j=���1��3�nJ���I{eR0��{�*Tl$��H�Ӳ�VE�AJ-"_��"���SR���Ҽ�>莮���:o��BR���:�yҴ��lç� ��ڢ�h\��M���(�ڧE>��_��U5�{׎����X� �)4������pi�0fa����Z%P������l��������AJ9.bRzJ��y�:��o�G�3��][7����r�\�N�e��s��y�'J ._ߪ�&O�z���$Q���� _�ߞsP���5��<�?V�nmmf�.BZȣ+(�$9�&�E�e�h,�T�-�mwܒ�� �_$˳�Za�.�1@���fy�-8Ҽ�)����h�0}���E~�*��Z7���dA �]�r�6��%�8��h#�ٯ�xu��O)X���M@� 0�Q�dKmԔU�d�C���K:���[H}���9(?a��.�����k)�sֵ�����
`3?�H��
8��LY�jkl�85t�T�-Ɠ*��ꤱ��7M�O�
� �4Rպ�:��UH�`¼�J (��)�JϧD\)�����*_�ܪ��u���U�_��ٗ�u��Օ��[�ח��������vO{!{�S�<e>�ۑY�ź�eª��T�G�ƹVd�wˁ��=yT%p�|�}N�e�GYE ���(�3x+}Lc[d�tAU��ҏ3�̃t�[��������h{�V�b�����.�i����n��Q��� ϴf4*ɶ��;�C�0� _)ŦRh�������v�-v���\���C���U��<Zu�\n�1��zq����O��I����!=h櫊I�X�8&mA�Ű
@o�h����6Y12��$_Y�=W��o<�&�flSNRHI��z�e����P2�ԧr��͢ꙙ�ĐO������i�t��Bu �(P�0&��_,���{K	a^���??����L���+��^S����M�B�O����T���ԁfπ���%a�0����k`����0U�[_��H��1�#ͻ����&	;�����ߞ;{�7��7n\������{����E��a ���߶qW��Qm��#�7�sbޙb������{�����)�%se)����܎�!�X
�8oeR����"5�]��tN։�����7t�4I��x�@��X_�@H���P)�m��Y��mS��7K̘��^�����7)T��Q�����t�e����5���Fn~;g���lR�O6-|U�㞪$�P� ��*��@�4����$�b��&��PB��O��9�ۓJ,�-&̛2�
�ƺ��AUڟ�JuڴA4M ���Sh����o}�[�K�赱��0���|��'��Q�W�
Oc��g��W�G/,p��Q�R!`���2�D�Ʒ����R�;�)�^�����u�W]���
�륽E����؀,���>� ��=K �F�> ���c�DXH���7�(s�*fGC�.��殄S��b�0���V%�6�fJ]!$���<�	5�4`X Xy|�R�P�A2yN߷�*)��� �$���IeZ��K��^�g�V��A�x����}h��� ;���e_,$V7��o�&h�(]�����*-�(���OSڦ:� � ��}�yi������e�(�����&M��P=2�J��Q�D�	��Ѵ�A����G�L�#�z���w��E���s�~�� ��s !R������]��m�zMo���m�g"lY 
�t�y�_	-}�*�&�L��<m�/��=��_T���u�u��W�ӷ] 7=��y���?���K/�d�����`��h������ݕy<< ��W^�߸1d�УM�H¬T0�L�-�N������ʲ��p��B�
Tڣ���I�]��wI��GeW+ &��F1�MKr��3) �ےN3�f����vU6����[�Wk��{��# �������v� Z, s�3�@��M1q�1a���R	���15�*�{�0�UR��>��0}�w΃c�SkAUTg�H�$Ȑ	u?��^��<��d�'�9*TB��4H�c�i����P̿�G�xN�@A��Z���� .k?�� M�'� � �d�3F�e�SNPiu�U���W��(U�4�bj����[��(�
d�^c9�O˺G����s�:唗����)��>�O*P�[A�I��<ɥ�������EP�V��#m�4fҎ)�<�L���o���@j���/�k\��s��R(���9�u��[�J�{T)�;K���z:g�{���,��A�5O��[U�b������^u�L'����Ѵ��i�OG+�����"�D{EPl	 f���`�Zy���fP#����v.e��6V��d�������az���~�Z��7�|s��xX�Y���c'i]J��G�BҌ��(}��g<�ߘ|��B׫�t��me�Q>��R��&�v��z-����H�߆�(��N
i��{<�ͻ�B�al�"v�4��|���G��ʻVe��R�8�����µk�l�� �h���o���&�h�^/�
PBS8R�%�C�~�iva|�O ݔe?d�k��=�kI�'�c�l���k�g��!��J#D��?� �! m������&�����?`O����ąF�����9D]�����}���P?�S�稏���16�ør/��O�ύ6q�~��V�k�~���N{%R�>(�^�$~���λ��K=����<�<��'U�^Teu�Z��ǫL�Ӳ����[�L�Տ_����X0�j�0S8�����
@Z��Z��v���:/�-|X��<�P7h��⭏Rk�ˊsEE&Yk���K�[L7��D�-r�f���[�5`�3���l�jm�� �݃���%]X �dax`Ҁ#���N��������()z*ٓD�c���/o��Ny�1oIs��Ϩ�ޔF��o0��6𷀷�.�~!R��S����M���:?��ق|P�t��ϯ�ݑK�3E�].֥~���x�1)e��̴�������M���*PѴ�vUL��� ��~h�V�����/�˗/ ������φ�^{;�+] ���L�������[��=X߸/� t\��:@9 Xk6Srx��?��e�K=�<?�]��Z��r&߀Ni2!�X���. ;��k��R��^��w<�KY�i7�E��Ƴ�HX �/2��G_W�[�u�!�`������f�ٓ9O��E�s$`���Q�O/#�q���������12a��\y���h� -˦S{T���Pux�x~�������ޣ���`��^ŉ�� O���js��lU]����c[є�_���P������u��QU~��v�4vh66��935:7�cq� 7�]��-�]���Ι�±�PP=r�$R�V\����Zc]��vB�L#��_���/���"Uӎv{��mfV̢�n�s�,_�o&�u��o|S�r���6��b|������eP�1����"�����񀑠<~c�^��h�Ny��(���_�U��0���E|�aW�a>�d+�7�F���Q����
��q�)���c�p�\K91�O�yj�_�_��ʉ9�@xR�i�t���W��, �Gq�G�L�e�2SF��+틟�{�VPk�\�9 �A&��X� [h^�������{c���'� �%�-��W�*��� ?������G[� ��5h��D��׿����> 8~���k�*�,�c�|>^φ��~sb=�5�V�O L9�?�o���Ԙ��M�(�,7ډ��O���!�/~��ꫯ�P/s�y�:P�ޅ�Yi�h3�po�g�!�ô�g?��=o�/�����8ךA�{)�������2���~�(�Cs\Yt^�uHkL{����J�}~���>hN���~�㣙�Ϫ��'�e������Ve�������*o���a��7U�n���My�\�s���(_�xp��kN�H�� �S�"�X.�͵հ��δ�X���l�˞�$i��3c���C]:ۖz�\��h����)&bȵ����l٧��ogÒp���ڷ�� \0�mr{�1\KK�;�y�4�����C���x� ^2�jYP�c�1��_O�'>00 ����ƍƁ����Iyy�a�؄�^6x��V��<6���J��Ǻ�7������C�}` b�o�6sF�v+��B��p�&�P�W�y�J���K�0�S?6��?
�ARj1�Whmdnx� Ш4�x�2�BZ�.��B 㨽gU߶%�v�?��� [��/���qY� �)�xr���J���i88K@m,��`�����D��k�ӝ������ �h�\�� ��}h�b]��h�8�i�`y@5�2.;Ʋ�S7mdWNz冧4��K&��Ͻ� Ŝ��6��?2sfݑ�T�B�1�8'�e���̶�0>�5���3��Y*͌�	`嫭5�P�V�c�OcT�4�=I�����z@�-��2~����{P�a�My%RU�������~<�~Zߴ\���(k��l�60[�(��-���h��V�y��>��q�}��y�R�-�%�f���t;}I��ߘ?g�-5���&Z�M���B+ݱf�Y
 �>��>�  >c�"�,��[ے�����/6�l �l�J P��ϛ�
 C<K�K�=c��0�A�5H����?����l�0
�B6}�E�� ,J�C��_����H��C�x�Y�?������uQ7�z��@�i/{�q����p���p����&�Q��3f�{�Ǝka��#�&~�w��(�	�t�0����u�#��A^��o�O��m��נx ����-����>0.`Dy�OhhD�W�(��)Q�Y��+��*  ���5�2���x�R@){�)ZQ̧y7)�f��r@&�&���z+��o�c|�������'?)ͼ9�� (�Ⱥ��[o��8�Z��:�)2�Ѿ�������}���k �� Z���_� ��~���,���oƓ�$lFH��Ii��SEו���%�����0�Q�̟��jP���>�Ni��Q�T�W5�0����C�X�0��8�iKL��sk�_�w].<s�I�꜄������N���,������POz�[��fcج���	l�JtM�j&OD�����͇�����5_��x?��� "R��*�zZ�ͺ�=\y��V��7�M��1nD3-3^[ˣ-�ϛ�m�����h��;n"��*|Bs���FM%��K����U�Λ@{0�M�|�L$ۀD�C6b��Ɓ{0������(���
���a���g�\Q �������0�<������/��	������}/^�T��1)��Xri('_3EѤ�*�~����'��*s���C~,e��;�R�QhT�a�L"�u�	����(�ӘxR+A�Y�X�|yEǇ�~��Ǭ� Y@1k��yZ����u�}�zX� 6e���=�?���oXåe����������`�����`�� �5 _��j3}���q�^?�D��q��z��T����ԬH(��$k"��a�j����2Ș�D�.��w�dɪJ��< I^�d�9j���]���J{ף�Kx0Y#�\Se£�/�{��wR��=��+���_�K�<8X�5��<�I�wNY6<�uڹFu{"����*E�a3����,�	��_�#�le�Z���57�vHV�E+�>3��Ԁ6��j��e W�~;*b�\T���y�Rn&���bo��l�(��6�>u�4� �Z�ٰ��Ih0NJ�ܪ^&���Gy��ݛ9�eS&R� B���1L�U�t�-�3���Q@Z�������s�р��9�&�50JbrDԭ�bP�G�9�6�4�WL|�d1���|2�F
CDY�,��DY1p��>�5�ϙ��5{��H�"����!����P����SAe�fT�u�����J�O;�>d�Aĺ�&���� q�۬o�N� ��c����6��>e͕_�w�Q;��P������~+���oh#�0Zk̪Y{�����G���������f `ˇ5������RNѕ�"��@k|�4��~��P������|Iq����5�_8ƽ� �b���ʋ�tO�-W#	�鏴�Ǌ,^���t�B�f?���/<�����4M��%�'z�Y�����R�A�g���u�T�@��@�`R��b^����@�r،�������� w��0�婓��Pَf��\�)Z�)�l�;gA�R��rm�]ȶ}�)\F|."@Az���r�%4�->��F��֔�*���Xd
l�E�pŴǶyLU�Q����K�،e>��ތ��"�1.a28��ʩ���4 21��,Q�L~�����2���n,>b�ĸ�� ̢D;�ʟ�r0)lZ��qF	�φƵ�_i���L��s&6L���<R%�h�ѩ
�YB44<M�\|�,+��ѳ>f�.���>�6�^!,D8���Eެ/��H��K��U{�אx��L�u�4�])�um�c���+����̶ۛe0(�v��g�6ˮ̗@�ۛfQmP0*�'Վ{�k���̲w�E�yH�˷�i_� ��Of̲�JcO(@��&����@P��R����ν�@u~�����F�יs�8<We�@q#޸��#	\S-�U���Jϱ�$��V{,�n���[8�k�0�F�z���P(b]ķnX���onZ8�sg�[�,@�i���L�縧X��,�hu;�	�p�e��L!�4�]����nn�lm��F	�9�|g��_�mZ+�2���ie4�'N��<�IƗ��|l66�m�'�v�d%��eB�Y!�Rj�Hfl΀D6nv�i)�&�H���{��U;Ɔ .�a��4�{�a.�T�S�F��ސ�[ѣeJ�q>Y�� (lF��2������V�M�wiP$���)'&cB���D^e��?Xc�1OS(5 xw�k���Q��h��i��I�Q}�<	�ؓ_|�%[�X��b�AC (�Y�\Y������G������;��o=\�4W�4��6���i�d��u��Y$`G�)����˿�0Rf��	0��-2k�O����W(�L��a��̨%��}�c������|lK`�F�{��"x*
5��ߗ}Bu�|s4��/�y�E�.��y~�|��J�K�.�q��Y�A/9Oy�joU��q̻i���6��_'- �AB(	9�_pC�Gz�f֎�����ٲ����y_eA�Ӑ��� �~/�0�C'�K��_؂�؅� �9@+M�U���ӰP��?��R8;;��&q]Y]����ƅ�1�L�V�*)q!o!���M�# nfI,W�r�����kŴ�wm� ���r�eI��av�S�!_�x)�8~2|��Ǧ����v��ת�Ir�J�Δ�Yux�~I�e>��.�\�}���͘�^�EB���R�(Ӓ�f���F�p�-s"��0)�����X�\�ƴ��Rɼ��0=ژc����U�c�ʷC�m�n�%7����e&�0(�4����oL�mNz���;h���}a�>�����"pS͚źL0�'�:IY�#V0�K�a~a��.�@��N*-��+�Ts�����z`���4����0�Ei��˗�{,�����b����k��0�+R4�`]V�ż�Z����0m�M����$P���;/Ǆ�ᩴ�2���^%W������� ��8�RH�U�X�@Y|4��R�G.H���\�S9}*�Sdiŷ�k�Fi���u�WyA��S��}��N�Z1����t{m$��߲r`��@�a�� �f�J+�:s�A��I�O�������[�|�c]@�B
8��,%�*���G���a^�Af0��2[��^�j���~�3�`>7�;q��_vȺ��Aj���3i���09s:|����R	f���|n���M�M�?s3L�-3�6s�rc^0�qn��@�&B��K�A�����?(c�l幊-�w���Bd .<.>~1�?��u~�ŗ���?+��N2���K��#��ԬJ���|m���m[БXr��bL�V���4`Z�qi�����4K
�1� ꆁ�m�	s�h����M]0������Ac���)m��vlV0�֋h��F�h2��^�PKC�B9���,���{>�b�7J%��?�g�9)4̻��+e�X�X��s�z����Ȼy ��(-?\��Εn#I��\�ND|�e����R���',@��� ���b=pk11#X�z�u��@)�=9����eγ� ����Us��#���U����B�a �4�/^~�4▎��gm_@;N����E������ DP1����\�ܽS樗���?��]#`χ�|��f/3k�8��5�'���V��=FY.�����S���S��cau!������*�;I�~t�p�{0����L,�B�>k��\�̄3Y�g|w�i)B>�%oߟ�aM�>�W'X��z��Z(�kW�ZT|�ZY z+�G��w��3��Qǳ����w��́�(}��� ����P]悋O�FXZ0}]J�O���T��B��ܟ-�fU�3�<�!��R��v�9�2�[n��&X]�H�ka�LR�[7o�M�E�F+<�����53�N���ؖ'�z*<q�	���b�ρ��6�I�����-��PN�^�&�� 3�<_Na#���!��``�e���WR}6j�|dc�QN�t�#�aÀa����#�I�|Θ�<���CiҜ��S�>��=��m;��C>n�S�,ƃ���	�+r?&w�i��w��G�&�Y��ﷷpN�8�E����~�-,y`����������!�?��(�:��Li�$@�N3ý{/�<s3~�-Mm���(/�\�u�  �V�-� c��#� ��CQ���������ʏ�gi�]\h��J�Wy����iZ��~�=�
�W�Xj>�/�\��~�>(!�YYY5�k�$n�*ӲɧZAi�R�)�3m����h� T��G1����J�j�O����6�I�U\s�v��Q6�e�i�E���أf0�,�7��OyjՒ��&}�'�?���@=-/�Py�YKY'��Z�z���I�i�]i��KC{���Q��R�7��� Ky�PD|tB�� �0�@t�0y~��g���&�v��!�A�6�V�x��b��D�k��ہ�: �bR��.� YT��_�;qS�O�GL�67l���L�b�y��<�,}������凥��4�ZZ�d����&Н�H��5�#r$���\DS���)=c�tD0l�,�00;�%L	��b��P����vq�e�VQ�i�L��8�����,t*]�4�>ȉ���f�6�h���~�G�OM�ZE�fq�~iI��@�� ��/�Y� ��j���z!
��^��@��V@T��2� �< K`�}Wn"��h<YW)˚'/eٟ�;��<�(��(����o<iR�0K����J����k�����/�3�-�6u3�0��Y�j�Gv��|vi���ǣ= ����7�'��~������Qz%���wߵ�������ܲ63ތ)u+���_���������3܏{+�#�@ ���3R�#Ɛ�@{i�2HÏ���xM$ϝ>�|:�DU{�>���]��[b�������E ��#<QP�T�^�{�m8,�v� WYC�Ǚ�K!Ļ����C4�Z�<jh2hV�78���db
s��^*i�x�Y�y�ʫǆ�$����⾵��7#��td��t����ͦ��
0��_m���̙h�w-�b����:>��M��2.��؎�·�"`c�e�1������I%���MM节=9"[3��-��Ȥ����~�L��{%GA�X(ߢ7�CB9������;��l���a� �Y H��$�J@��7�TA)�"6����H����,t��Ń�GߨK�M`Z�&c�3j���J�J@�o�,֣��\1F�uʯ�\�:) ��9�KZ�FM��ҷQ/�:up^y�������f�D�!�*�Y��*O:m����5� ���JK'Ɵ�Is�`����[��O�$�fo�^w������C�KyrEj�6ߔa����3��~(0"���3\�~�v�?2�����t�̳��ɺ|%>W����>����n���gθ+�bvp��p��c.����Ҙ
�x�"wԅ����n,����y��p��ⷆ5��q�t�g��Kϥ���/Zcy����Q�X�~���k��w�����vS��Ѭ+���(�m���!�
��e#b� � I�%Wp!^|�VfV�b��}'ߤ����=N�E���3a+\��%nw�h� �V�lY+�Z�@ �f����a\��/>�o��h�Z{i�6O�V�1�����mx�L�i�a6A���ݗI�t�b<XTl��4�NøC�V�L	/�N�Śg��+������*�}/6Yk�+<��䌺���%����4�0
�<�b������X�Xx���!��:����t8&�+iH���?��K�?S0 bA��9��F�~Kk�e�m���F�:L�sb�ߏ��q���NHk<��r��7V�PB_�F�y-�͊�̇kY[Y�)Ϛ�y�`~��-����Y���e���`�F��q4��;��/[	Z?��s��^�Zf��Z������ʾ���~l)����Ң*p�L�\���TH҄s-�И
��7�%��m��2���XC�E_�s�����
��ߊXMJ)��2�V{���o�</I��7��o�����0�[Ϥ?�nw2���������ϖ��5�o�-�)H�L
�{�Q�Yi|�	�������v����TH�d�$@��o 	&�����#�V�wd��@TJ� ��	�s����8#�@�n�__�膞�t�	��my�_6��++��TL�ܜ������ܬ�z�ȍ���OY�b�ĢE�}0�ߔw�����ӗا�cĦ@�����K6�8�[`O9'�93V��ubب��n~[��8�����hf`�%�%I6�B<�a�0��ˌO�DD��RF��y�lD2�c���R1����	LCb68F��L�4>�[C5�Ш���)C�\�&{M��!L-���Z�8�(�s/�
��6��+�1�HK��S��,����k�k(�p�#��)o��/u�J�R+���?i�|�x_&�h,56��=����3��2a��!�E�#���v9m#�y��<����q` O�W5�Y�����4�5U媞�AP��l�`���b��C)��sx���4�$���@��T*o��Z%|�;*--'��4�G�vɥ��S�_`{N0�f0L�z  pA�K�A �[o�eF� ���n�vmm�̛��s`s�OF r�4�P���Ǘy5[l��*ۆ�Sa��3�����X�e���6 y���qc�S3������]�>���rrk#W&�X`���x K2�}a�m� �庻w��z1J jRG+�ĨG�gb~�L`��!̀7�V^^�����)�__;Ȧ�*僤�fWD��u�A�L�r+r}cACL�E��lP�M�\D��H���	���wC5�P?�NT�P��C҆z��M*����T��[�=�N3P�f��M�R7�>>��'X!���~V��5�u��������>i�o��}�[�H�����0�-�Y��b?�$�D�*��Ǒ�z~@{�w� �[����j�^2�U0.H�e�Pu�zŬ���z�;ݧj������ΫA{hjb{�J	/��Ǽ�D�rBi�|�Q}F'�LT5~�}H�*��ID�B������Q�aR��Q�Y . �p+�5l.�8��fE���F'��;���(�+ ���@���Q� %�����35^��a���M䕕�eT�|s��~Ñ�p(�_����7��k�ac-nF[�,�P�W"�l�,NX�ċf���ϗ�<ׯ�(�;�MdRI/ς� ���@uk-�e��K����R�.&F�k��|�lG~���)2�EO�dic�>1"�u��J)���z��N=uc.m骾��6�Pd��14����0;�����4��'?5mP��+6W�pT1>5�PC)�i��u�}w�aJAsi����Q�ֵ'B���^C��������7�Q�)��!Sb ��uu_	m���{��*�I���{�<[�%�{Vm� %�L�<��}�NÜ��@���/�]�|9_��V��!���[�Ҡjn���jF�gŽ{��L��P������[K���-x�tcZ@p?�k��uV ep�n�g^�V'5H&��>���'}�UQ��f�03�
'��`O0�WV�&�:]�xq˿{�V4A~���>?�яL������4#��3��flM7���CKQd����b3�r�R���Gs���[�z���V��Ri!
e��� K���b;� ���?7����ؚ�2S���w�匟2���"-���ԋz��Ď�$!׸���4����B+ļ$�^{���M)*�%��e�� "���[���K�u�k"�q��M���PCU����cR���o�<�O*����N��y���]�&�K��UZO}�eуŰu=w�!��I��Q@�y�l���xm�tA��f?�תm~d*�#j+E�@���|�aN5��=���U�J������u��g�_<�����߻���a�;�}8}���������݂߆��	pD�P�JU^_�a��fy����y^���U���5�b�~e&��Y���a6���N���Ϙ%0`sk5��t���m l%�7?lhz!�m%�&O�/_��e&��Re�41���jbk>��0/|ɺ\���[������؜�=��F�{��	kק�+��ϤS�Le{�Tǀy�g�zFyY�~ԁN�H������G5�yJ{^E��i�j�����~��3�0��
�4X���%�}@,���j��yҫ4l��ۻ�C�u����I8��g�����7�C3�-�d��5��~�
Ifݲ��g���3���.�^K����ǫ��0Ӫ�� �������q�~Tw���>�R���^�e��x���k�~S%�	E��
��^��R ����*�j�U	��sn�`����Xc����6��i��jๅ�~O�sΘI1��Yk��z��	�F�����F��Q ��㸴o�Ҳ�uBwo/v�[d9��m�����8ϖ�'�-��.��ȿ����=����w�t6G��f5�Ҟ�j��i�*�T��Δ�`9졀4�P��쵊�,����9�v"� 
��z��p�[��ha˥֣>�N���Ǳ���[�A���q?VN^��(��S�-�zʕ��r��-c�ƃ5	���\|�e�!�ԔaN�*AB?^g��~h��iЪ@pJ� �a���u���AP�g5��oXm]��O^�!ˋ:E4čw̏��Ke$�k�f���c�����Õ��p-�έ�NVD�9�E�fp3���,���I�A1�в�������L����7��N��y4���z�n!��;����?Ν=�z�Ik��4���js~��Y\j�����ꄌ��AA�H����/��0��=V9d�;33kq�׎� I9�㎄kBi�i|o�N�G��9�Z�x�C�9�9��J!TE�]�߇��H<��|�;��@,�P��I>f�;�X#��W�^��*����}��e&�����q�d@�@� mx��O��ǃ�	z:v�Ώâ:mo���7�"4�a@��4�G��0�������3�-�X^>�{��UD����	������n�c��f+�a׊�u��;��my�PT����)���D�����o����za�ė �Ŧ���#3�����͇��|8}�T���
�=�\ܰ_�@Zlp�<T�{6�ILw��o�Pm���:z�}`��1������3�Y���%i��������o���<��q-q9^{�5���W�*���	��CÚ��ӟh$�
���^w����)��W -�D�L0G�Ɣ�N �nK�����/��/L(@=���+�p�ޜ�Ԋ�E}�B��S.���������o�<B�m�/�c��;�SY������iz)�CM����A�]�P�̇�c��*F@����Y���(���?b���l�ǎ���M`e3�[����\H�-��2i�4ؔd&�q AE���Ħ�Fw'n�l��X:#">wG�s�`\�	���?s洙3!?7�'�x2<v�m�Hu�D{V�` &V�LY��6�PCY�ZE>�cXR}�{�3a-VT쟞(�^Gl�o�� 0@S&�*烼h߃i@�;��/�8��3 �}\�{�ա��~�S'�n��y�/�IJ}a.���>�r4�[���N�	d�~J��S�1� \�����L��ƕ��O�0����kL��ďU�9�nLw�+�w�TJu�דBch���_}�	�xɿ�~��y���%�~Q�ߠ��}��s��][��s��\<�b>g�6����|�\i�[�q���6�ƞ?xlJ�Æ!,̏�|#�����D?��Y�u�VX]Y���@(�[�ۥK��g�y6<��������.��Hn�*R�( ���PC5�PC�E)h`���J R��ĸ�o�3��b�HCC��/���"�X`p���VR��.���4G6so�c>��'"� �p��e��� �(�@�����)��Zc�>2N [��=��n���)��R�G���t��'?1�����4�N��ԡ4{����4������~�y�*�;%m�-�������ws ?h���6�7U�����^%�Ư<ӣ4'��u{����)��<[�3����;f",���t7��Q��	.��:Q��Y����:?���mv�&���ֈΝ�4GP+k��ٙRBN.��}�Qϝ;k��#>�9������f��WR�F��PC5��AҠ`+u����0Ȭ�kzr�0�_���ow(,� 8i��OK�Ҙގ{�R�K}4h�T"ܦ^@�r�s_�R?|�cV@.~����`x�%��/.)�(CL�,��꒩4}1˯��teJM9�CS͸�l�����%�̼�(1�G�N}����V��80V܏2�9<���h�j#�Y��_��\�8�KY����~
�ŵ���naQ��N�/t�| ���Vi���0y�A���h���
���ݯL�mnl�|��M�X�B���HcY�;�X#yS�˪����x�\{�]u3�[�
`�-�y���m`+��b\��7��Ι�8i�Pm**ʤ�V�Zm�����w�|����y�g���FX]_�_����o���[J�07g��'����a~n�z���\��7o����Ek����N���PC5��tRU0�~����\��(�w� <
������t҄(e�\��{,`�am���?6p%�,&��d����>�{�4�"�f�/��/���	���
+0E�Ve����sf '�_�J�u��o�-��s,p����,c2��4u0n�ï��$�=��s�4�|3f�b����h���s�������+��b��/����ߴ팁�͸�����7�4�/�5�o��o >.[Ќ}�y�O�%�ꭷ�2�� �����a���l� [)�;W�Ʃ�
�� 0��kT�1�A?����:�!4�Y{?aG�{&�U��Ӂ>�!�w�eŵ;���U}����5 �Չ�w%<�� ����`q)���d(�q������2A$�eAGb��HH�ؘ-����irٰ�GP�&��"�eAǿ'�.`w~a�6o>s�o|���g���WL��80�b��ַj`wӷA�4�PC�#֬?�KU ��T���}.?4�2���J#�-�8h�@����7 񇯾~��kv��tnv��`|^l�:@#����k��W�VS>�2����U����d�/ ��B�ds~��(χ������X��JY���`���vb��Pw[�.��G@R�D͸1.���\܏c��1�[�z�+�� �.��@��sN��9�\�r��N�ѯ����q�E�n��Y8c�]��i��_k\8F|k�X��n��e�ќ��i�Q���h���=h�?;�|U)5G�G��Uȳ�粭�fHn��K��{��.���W�7lw���~����CȢ�7�6���;n�hu��B|?�����<�&�X��尶�f��h��ef�P?>l
��U'}o���j��âA����${ �F��� F�\���� 	�$S^�F�޲/�m�������R�&� �x܋_}�U3�U�f�`����\n� =�-��1����8/�'k�% `O��m C�	 r-��>pϿ��_[��ޟ힌}&�3u�S��8}҄E�%}�	7��>L�I?_}�U���o�m�w��駞�gE�e���| �h�	"��t�J�RT1&�Wi�Ȩ����w�!���_�����_��ԺS� � |��N��(�4��0��Jô;�pp��k����N:VW���=�=r�ir͗�B��D��0.�];G��� �7��
�S)-%�ީ\C�q�}�F��pl!��H�ɸɠ�&��I��" n� �G>>�>ʓ���j���K�j����?��:pe�c��r� p .��0Ƭ�]����}�g�	sjZ������ 0c��)#J�c�m�4�����f����]21�CY��8���~ �+]	�>�fm���U>�+81�9������-MSdkƛv�'�z� o�F�|>׮]�z�<{&�O�8  4�p���o,�H!E���q�|����pP��1�(C��;�bͽ��<	)����-���w핆�!�t�j���̓|��5��xՙ2��n�.�z(*~2���N�k��Y'�~��Y��@
�7�4�8@v���0w.lEʙ?Ӭ�8�I�1 �noٷ����ߝ����>�Y�n���jhڈ=Kf��>��fej,����B(�G���*���~����π(��`�쟀5��:hYeq�v
i� o/G�����M�:Z/�mx@0�L���=� �?2��{�n��4�n��_4�~�ͤ������_�e2n��rK3 0�R�0�)��ז~r��b�eƬh�f2�0ocɽq��<��o����'����c,��g~�ԝqT�kᙸ?��#�����_Ǻ���O�OC=�Tg�~����B����&����[���'�n^�ɽ˧����骝�Qu�S� Ե��'�̩�7=s���pl�;m���Bu��PC5��R?? ���� J�,e���!  �IDAT̢����h��>�ZN��J)D�@��8�J��	6��̝"�� �"SWQ���Ahv���? �k� M�/m3����|p }��u��� ���G���A�c�HP�0��H�XM����M�Y�^-�I̴�2h����3e����YPFf�E��|䋌% ���,ῂ�i.�`����AP��
�q��PC��2��L��`�uu�4�l_� c�KI9�66Ͽ��U������<����w��Q~��u�E�0��b��v�����.zaC5�PC&��"��	���2�D`�{�O�SVl�]�RT���囿�V����P�d6��� �>~�Ō�z�nL�
?�a5��|�-�L> `�Ž��	`���ꏲ?p�	M��.;�p	@����=>�	�2h \E�&�5m��<�&��*�p�sn�==8LǊz�h�9Ǹ��g?��*�q��HW+=wX)��mx��:��A�5@�zJ�=�����N렴G���4H���7E�4�e��t��%�nQ��O�̳m��B�k��}
�v����͂�PC5��$Qʘx�|��)���tH�Ж�(��H���O�4_D�F�HY��4��)� 20g	�3��@- �(�� �� �O�������$��G3��[��d�y?�YM5��Ø�F��8�6�'`������]j�1]��7�ch���Lkl}��p󼩋��4��dk.��N�4s]�F�nn���UB ��@�z��àa�+k�Љ�*�pؖ��Ώ:�t��Y���Tp�v����s�i��2f��s�)�}�\��H�ӹ��ӡW��k�ݾݤ����au�9w�ē�'���j��G��1�J%��4�R�N^J�k��I[�r�.�k�]J�B��A�/L�僋9/>�
��v�����>+3`i:˲��7>�\@-ZL����6��`O�����-hG�R(16�c"~��eӔRV�9L����Ɵ߀V�#%>��m�����M5��_x���:����!��:��k��`����<c�&���<4� ����q`�0��+�6�O�+���p�����c?��P�����m�9�|�BԴ�橡��IB�J�Ls=�kn����L�}�<�.�y*�L׿A{֤?�Y!����ܡ�d�K}.�:�:��dq���П�'gTC5�PC��۟<�j����9~Ugi~\׵i��<L  %__�� W�0��כ�iH����a�f��A�0���G4�hYi3 �>��Їo0�]���h��~b��1�G�����~���-�@V� Üۑm�d�s�h��+W��~�h��� |���0?��t�f��m�����y
OQ�eV-M1D�D�~.��v��_��,-�Va��o~��7�W��{�lO1��	&ҶslҨj,����/ì�CVTk=Rw�׽�����*K
���N��N}w�S�֟�F�����O��O��5�PC54I$�h��_ԃ+o����:M��6�o�Z@$������mK�� a����*PV�D%��A�����`)Z���U��!So4��NLv� 8� T� �T�7��	L����
>EYR��������_}��qf6�<���_c!�����&$ྀi�,�����63�hv����,5��w�)�4h�|�M+�13��vB���5�A��ԓ�pOߨ�����>��{"�`\���d`���S��=��U��a�,�iW�L�z��&��������+9�4�|u�	t�3�|���z�׍��$��Oz�Q� ��Z~�ԟ������F�=�Ƣ��{>VY� ߆j���&��O���� Wh�  K�V����QcEEV�ZL�e���l7ڔ��Ἦ�oʥ�
���ި_fЊ�|��+{����v)]"m �c�˵���E�`����h�ѐʗ�_�/��#��|����r`я ���[�~��Vn�L�}��	h&��s��ZJ���8��<`٢bL�rSo����})C��y�eY-�G�O�
����3Zf�9~��)r5�P*'�t�����Rsh1�iJ�~��Ͼ�B�T3>
�9 M��:�0��6�4ցD��L?���GS)LcA�.��{+���ö}T��s?��Np�¼8��awט�A��n���j��#H�z����+|t�JX� ��8��Y�~��߆?������(e�v�� L�դ.�����(��믿n Kit<0���o�m���y��q\ZW4��zV��#mZ�w�}�4�|3�m��2�b�8�5 \چf��'�2�`L,�x2��X ,�/��}�@���� ���[6>�\�� � �RZg/l��Ҫ<�i�m�X���p�{P��?��i�y~�Ѧ]��o�� az>����@0�)������J�?0Ɯ�~��_�!}��Ai����Lz�Ao�S{��Ak������O���9L�bb?��b��L��XJ($A��m�R���]l�4 �Q�m l�K�Z4*��Q�� R9e�w7���9ݗ���`s*5�PC5��"�� V d'o�0��T>p �Y/ @p�,�	�& H���O+���߷k�K4�R�S�| � [@���GхhP@�Vy��bt\{�����{x���9Ni+}���;��q,
�e[N��S=���d3��Y�	�ݝ��U�3�$>������rl���T���?� ���GX߮�%��7iؠ0w�xژ�iW�")�篾^o�a������)m�7�}�O:�[����Z,�9妞:2���Ro&.����+�-2O��s,�u\�/_���Tq-��V;~/��V���<F�q�r?J����K'|�N{�����T���\��J�s�^&Ș(#6�֋���D�h0`Ho�I����7=��:kp�8s���e�n	v8�c>4��꤭��*���|j��a�|'!
:�I���@�'�b�]�$c���-d�Q
.+.�d����<y�������ԁoɣ�`e�"���� �i)���`Ȣ��(+����������$ے��?�48W�l��4�Z�8+Е�9R;���c?$WQ���R�֜����q.��i�r��_�H{<��qhI$��$��ڂsR��H� KK@Yi���Z|o��b�̱�m�v��쓿�K� O��cI̥���z8u/��t5CR�cε��<O<?���5ZC�%�t�%_�R�y���>�C��tC0��]���vU�B/YG7�����f�BՐv�H��b�]�u_4��}H-�����}���p8%T��ioO��%_B��$�v{��%�g� 	D	�e-����es��`�$K$�	���\γ��L���0K�U`([o�g�vP���t�v�ѵ�H��U��`2�|+E�V4mg�>u|l�9��%/�Lن5�v���3���;�rJ*i�)b��� �j�>@Y&/��ݛ����<]3[�����}M�|��1�5��NC����:~L��C�S&@���XX��I<�&� �l��&�T��Z�9��)���R:��O�NF�Ha��Wב��p�H~���"�D��,��dtE���kB�W��~׫ؑ�o���:�n�SF_����[�Y�I�YwR���4���/�����;/���t�� ���ׁS���_�e '&������Ur%��U9��H~�#���}��9Ɂ	<��ZX���gh�)h;x��9�n��ה"i[2hIo�d���1�@N�B���>}J^�y"��)\Ȯ�9s�RU�h�:�^�ۺ��BxT;�|.?W�]���ہ� i��k o��ƶi�Ө�3���T�ڍ_�ݣ�)U�#�0��'1�,�s���{�l��f��|r��L�ɍDd9������'�p��W9�(�!�)�UEcԑ����D���H�o�n݄�冭����I�ߪ�>]�]׫p��J|I��o���:�b�V�lo�<�!EQ�Db�i��	�Tz�_|�'���������9��PZ�����"`׎�|(4�R�.V6�AC��
?S,��+Js�1��T}NŔ�lL�8�]�ӡt�)bovȹ��Ү�]ژ��Xݙ`��b������
CёK��c�}*l�����\�c����"�.��9^�k����&�����@���M���[��z�R��\!bg����A}J�����zS}�U����&����6������6���DH��&6s �R���os���#�I�b�p����]��͆�-[_��ꞯ������p8�"J3�֒)	����_W��Z"����pƶ���	���BL*Ц�g�<����^�A�������7��vM(�d�ԇ6�I�K�+��֢��0;OA�9������1L���?t��E� �8��ÒI�8�<�ۜ�(��@�-%�c��������,�2ܮo���N�7�wm�\/jZ1l�!HA�	=�3�d�mg��)n�HiBb�K���;�lw�L�c��wש!�f��Y9���ܰ�LX�U �H),�|����7F��|�J���wH�({�X��y��I,s��ka�n�Xq/RW&]P���k~b>��n+�t8��)��CǔT��ؔ�wC}�`��RH��D���8�l�I?�aCF�)�ũ���u�ό[�"�ŕ��ݱ�]�txM8����,�}�	,�_,�$�#|�6���i0�7�.�Y���nKb�u�����.VӒ��/Xd�ZZ�m��%�>��yc/`���p�m��Xn)��k@d%s�yC����0f��%����R�}�[9��^��7��~Π:���Ѱڀ8�{�����A� ����@�B�K�J��SQ*�M7'��,��������+�S����>�s���YPV�XWAM�� �U�&ØY
�߿�u�w&^��R��+dy���w�`�p�AS��O�h�;�ײpy��D8�c:���nZ���U�}?o���|Y���x-(���9��R8�(c���_�vJ��!���%�<��Ti\vq��b_f�H��S�fV���,��)���O	������:[s�D����|����Oѡ?|�P��L��=� k�>����Y��Y*@j���o�?ï��v��$(�e���)���i�7N�ɉ��SE8G��S�ޤ�ݩvݗ�ty���;���x~Ysm@I�D�E:?g*ݷ�)�?����FjM�����{ж�UU?�«�&M����d�S��v+'�����o?^���Λ��Y���ʦ����@Ǘ,�Ia���I ˩��q�f���0L(T����>>�U���~�zD�<��&2|�|��.ܮ߅��*�x��Xh��[�����K�~�!33�jD���'~�$�tK���{�%	Y}��r8��%�F Mӿ�w�o6����8�r���}ɐ`V̐%G�`��eY�A���k>�<���e�	��DTǩ��gѵ����(��ͯ�;cX����0�"�mL�mQhK3e�/�V�6���
o��?�=�VK+    IEND�B`�PK
     mdZ��<�`T  `T  /   images/69c28b0d-a0ad-46f0-a190-03e6ecfe42fd.png�PNG

   IHDR   d   5   �0N  0�iCCPICC Profile  x��||eE���6�G��y�]�$�{�R�f�IvC�]�%�l�l#[`�H�"Mw�J�"�T�"H�&E@`��3w�N�]������@��79�Μ�=��{I���挪&��y����L��ǞՕ^IF�u����X�����#�Ox���{�%��H3������;sp�@�4,¯X0��Q����- �~��{?G?K�0��g9z�xǓӛ8���V�)�V]20}�n�$���^�0IV�O���Ṡ=a`ͻʅ��;s�̙I�*$�̚�x��ci̹���A��$c�Z�?<+I����{�\�FЭ�m����%�����<���L�Ze)cͩlf���:��լ�y��C[7MV2M��4�9�5�kʴ\����Ӕغxx��6���Y��"��t%,I��]�*��,iƫĿ,1h�HZ��x�*��&��;�%��I�8S�ׄQ�u ���M��{���K�<@u�ǵ�1c�%m��&���_��^[�/X:<4k��j4m��>o��Dғ�,�6�~{��ǆ/<�����{Hl;�$i����6�Q�\�`��}yl���d���䶶H<os
�R�^�e���vLrjr^�<�6�-y y2y5��a���D�.{7�pfõ5�6j�Q٨�u٨'FWF�0z���F?3f�1�c����M��{�������J�4o�ߎ�x����<q���X�UN�����U��j�w�ֲ�-��կZc�5�Ys�5���'k��k�θu�Xw�uo^�{�W�?�~��6��l��F�o��&c6�vә�m�ك�[m�b����R��~?�-��f�׶�f����ŗ_�撦��;�֫������fױ���`9G�g�.;mۮ�������p���|�̖�&������4~�;��~��]�w���ִ�Zw]�}i���'̘��5���s�7.��ߞ�w�^o����3�ۇ�:b���6�7<�w�6�Ȃ��wZx��K�?p�����!�~w�CO9|�#N;j���=f±W�k�?z�~'�;��S[O{��#Ϝx�o���ܕ�[~A������{~���/�����g-WO��랺�7���C���֭o_�w~���w�u�=�w��>���G����d��G<��s�<?��/��ʌ�����oLzkǷŻ_������p�G>�+V�~����>��kWrQ�aCo�u�6u��7F����5敱�[w܍+�3�:��o����q�������k^���k߾΃��y����x�57�������MO����_}�1��&4Ml�b����Z��q_>{�˚nn����W^H��>�b�\S��76���m��j�ݶ��C��{}mA��Nk�x�umw��ؔ�v~��cw٤Cv�:u��.����Wz�O�r�λ����=~��/���7_�֊�u�ڪ����͜3�p�f}g��C?������s�܇�=;�����p�EM��[��{8�t�A�|�!˿s�w�;����;b�#�G���|o�cf���#����x�'.��U']{�/N��ԫN���K���r�yg�u�i���Gǝ{�y���\���2|���ɂ��]����.�t�V��uE�\��U�|�Օkֹv������冎w����C7/��!�}�I��s�%w\��_���>|�ӿ{��7�~�����}����O���~辇��í�\��������'���'>����������n���]��U_���F�<�o+��ګ������׶}�o.}�^����<��'����m?��Ã����n���c��_���a��Fm2��Q���Yc�{ĸM�ݱ҂�ی���wU��rƪ'�v�ꧭq��W�u�������/���Fo�ކ[m��ƻm���'n�|�;�O~�/����Ħ-v�r�V{m��ˇmsJӏ�^��+���gϱW���ߪA�dV�kl��W7�n���-;N�ڷ[�O:����?n�f��Nyt����٥���ίN흶���]/뾻��cfL�m��{�q���o��[��{���x�l�m���}�f-�}���^���s��Լ�$��1��B��m�nKfpЁ�/=�퐇���w�=l��7;��v�nG����}�ǝ��K����[N�������ϝ���/���鯟���>�ݳ�;��s>�ч�~p��x�G~��A��$�|�����m�.���/?񊣮<���v��O���k.����n����w�#7>yӳ�|�����[>�������z��l������~W��߾gֽs�s�������>t��G��GN|��?���鏟�������>���9�f�_vyv�粿6>��c_x�����ˏ���Wn{����������eo,󊷮���8�����{o�k�k}8���Ώg~BH�#�Q�Z���>�ר�G�ї�i�_{Ӹ]ǽ����g���ʯV~�ʕ�^��٫��ƅk^�ֵk߶���>����_��FS7^���޴�3��_ܲq�/�3ሉ�mq�m���o�n�6͓j�}e����v6�D\-oU��G�3�o۾�ݘ���a��k-3'�z����~�ӟ���>���b:v�\:�G�n�z�{t�����f��Ż�f���\�͍�%�=�o�^�������|p��}�����7�>�o�9��m��������?|���-[��%���_?(9x�C&|G������X~��G=~�k�4��q�/�o9����0p�ܓ�r𩇜���;��}�1g{�������=�S�?��.�鏯���~�=���O,���G.��e?���+N��ȫ��Q??���9��s���/.���n��������7��WO��̭�����o���?�͊;G�n�]��W�g�{W�o�}�����������w<rˣ7���]���O\����<��ӟ>���<s�_�x���������^<�3^��o��r��w������X��-�����o���a��޲���]���g���Go}��O>\�p�����$��W�x�+v|;i��v�A���b��$+���O��ϕM�i_J	{�?�d�3�9V�qi��=8�?b��}oJ�2<88�?pm�|�A+6i����4�����c߲$�UW����Q��5���3�%����e��@����o����	���u}��_�{������ہٓ��z�7^�34<�W��M��(��y�Q4~���	�Q�x��׳�
�Q�uo�w4�)_������������=�� ����3�	���1��ch[��������1�����;%}�y��H{)��P�8|�/G�C�9����c~B*���~-~9������8�$^6f��(SX���t�{opPk=�#?�w�J�u,M[��I2�,�;�ڒ�I;�lż��[�{.r#���F�m0!�OݚZ�O��c!zP�1��1�g�i`7m��A����Ջ3��įyJ-#w��	�x���a�i1ֱ�>˝8�A �!���2l�¦�]IS���Gq��k��m�')ᘉ144�d�2#ѹj�g\������I�$�d������I�3�)������V��Io18�ªF�.����S}H�K�y��o�9 �fH�#���a�_�-=z���;u�e��O?f��>��/�����ygo;�V���䶞�����i��Ɩ�YK�̩����{����y����Y������U���3xn��X���>�}j�Ȯ3�.��Xi�nk�m�\m��_T��_Ze���m��V2Wh��3�[��Z;Zzz����{�:Z�h���O����7��������nZgWߔ�=�6�9������cZw_w[W��{ʤ>���JoK���޾��=���;ۦ�Vwo�Z4Xʪ���9�K���7U[�ϙ?ܹx�~C�����׻GW�ݩ��g�j��i��ˤ����v�7k�ĉ��t���v�t��:�wBjS�s,��ur'�6ZQSYfLZ��&�f,�f��eJYf+S�uw�t���6��wZ�}Y�V�h�i��h��6��czo_+&u���O���5���}RG�g�Lj�I�A{tt�AD]��v��=��%���gW��{�ͭX���@(IԪ�8�E�3�-�$�i��fj�ƫ��fV�o�쩲ZVc���N���Xi�:�t�ʴI=m�3ڠ?��Y�t:�8���ul��so���v�7��?wwC��i-m��܎���Z<s�ҫ66�xz:�M��ySWKo��}=m�NoñT�u��w��/�0��6KþHE+S�wNj���Fvjo��S�^ē[z[�v�����tvu8� M�v�Nq���d����=ܿ{:!��=b���ޞj��9*�;�O	ae-�ˑ�5m���v-�kZ5��A�xժ���U�j\�TU��p>�?�'�y�ʈ�3�,�"���&��*����jF()����(�?�)�+�*��헱�`����if������Wߏ��폣#,R���Tl�s}?�j"���^���6j�BK%KK:[���3!,�X�#��Tq]�FhL�;t�<�2ص�0�B�1�T�*SȨ訲��;�U��4g�E� WX*/Q��Q�,�R�V���W�&��Q��]���L���t�����Q��>2Yr�E�@ڌ����h�N�c��d����SS�IH+��"}͠yZU2]r#w��dF�1C�R�V2�C�;5nG�%��P��:�D�l4��b#�e���؄�n!ӌ����Y��~�a"-#���N��L��RCH���L��t�	bK�;2iXfhaIYa�jk&�L�� �*s���-Պ˨�e8$zTPB��dF�\2Nrˬ��W�p��=Q�ϐ\a3Hڱ�
Ù�֌c�'0�`��X-�7X-�<����i5�S=�jLm.�GB	�rH˰5�u��J�*\�N�8b�0�e5�H��'OE���8t�tC+�b�P`�2�_G�@��K��h�(��@�Lׄ��'�a,ܶ��H�Y�K����O|tZB(,�Y����Y��5t)K��p,�|4��`�2�DX�ܱ�����9����`�$�J��s'��fp'4rYc�l��@P����AjI�X'��TX��1�f�`Ka�i�q�Daͬ�U�ۚ��:"#���+2xr���`2�G���VO��+�|�G�N���q�
�Bp�N��zlL���R(-�Xr�U����=Z��z�R+;��C��x(�+lj��� 6KDHN���RؐU�����#�o��?B\�� 6��`�h]i	3ѩ��ㇲ< 8T��p*]G�L��
����3tU�FZY	A��*�����*@*!)����3�5�!�#�8y���P���#���4��G�Q��a��m���@��4�O�b�Va��La4�j	�%�����sKR��"2���I3�	�	djA@a�z8bBZ����R5l#-#0��� ��=[M�� �O�������:� �}!��'U����H��	�K#SY��&AJ��BG8.V�r�����3@�)�E��n�H�g���#H������r)&N
mD��M��:B�#f�VaVP=�� 8�
,� X��zB���S�,I�Le�uոF�u��E�J�82,Ug�Ȋ4U#�~c3 +��%� ���R-�#С4-!�aN��W��lM"��w�u�~�	!g	�}!: ؊ʪ	�%ͬ'4�6|��3򪁓����΁�HR�z#�;9�0&D�j 2,��0#�'��0n�V
@2�ei�:
Gk�_Gg�wZ�0�0�=��
�����H����`�kI88x�;����TI��:x_B.�����U�.�"T^Aza�X�)�1r��ʔdqFV�+Ek袁����%�Ṋ`�@��$�P��dP"�iI�St$?�p�Q��a��`�8���"kD2��?	���SV���=�w�_��Ffjd:d���*�����:B1�&�H��]«�E�ˎ�H��ړ�E�p5h~1Q}G�S$q������!���ܪ�����B�p
���	/	к$�ǁ@	��q@�̳Ba���e,�qF>�.��!�Np.�X����9�T���I��������8���!� $mG@��b��8���j`�@�
pP�=��)+�ē��QPG%a	J@&,��(L��F�C`^[�R!#Ќ��Đ����`�1��3��-t�Ȓ�����.P��I��&CA>�pTI�u `:Npy���RE�-f�n����3$��"��rW$A�&-�jJ�gGNF��� P�N!Q�[�b�{kT.%E�y�������|�: "r�EsJua�*�����\�h�C��22Eq���\|E�d��*r8GFi�zd�by����T 02��4P <��a,� {՟?#�,.��Ud1CE*XŎМ���*!j�����LUt��XU�1.��~� �
(oɬ��K ]�K��H�R��=�T1J�B�)q�Q �F�{4�k�Qj +ǖ�Ǣ� -l��9������diY�)�F���3�`=�*ziV�3.�TQ%OQ~&U^�L���#+q��ڦ%o�H.�z�H��%�5*\*rzF�Ukx�	 �z��U8�`�Zr�H�r[���^ZVE.V6�����P�.=$���eu�'BO@.�:�		]GO�8�9�*�q犒?�����r�)*��e��'��APM�<��*|���֖G�ZJ8d���K9׬	�W��rr�
�X��^�x
NZ✰s�YVO�=	;�dp�]�ӦH_ѓ��B c
�M���x����D����ʰ��PM�Rg�%���Lu
	!.#�4��l�49�R@�#k��=���Gғk���G�7z��Q��8O�8eje^����}������i1�xA+�Pe�)X6��� lܧ�Q6�ٙBl��Cќ��g�L)U>� �*���@���2	�!�ecJ$YZ���SaY�T1B�
�rA��Q�R�F��+�Ѳ0���9�L��)��t�ʞJ�U��K�&���\�0�.0Q�3T����*~�*2T�}�����zO�oJ5*�P�`9�T%^3j2K	�T�2N�mI��.�Q%�8H6lH��@v�D�dkJ�eѓ������Ch��AO[�5�*�'$�(y�礷�4�)�6�Y�$��-�	E7h$�?Nn����5�|W�'���d%ޤhAb��@��p�F���	�l���'M�w�0����<��HL�x�(!���t(��t
cq	���SD��s�OHN������9hp��FGM�T����ܺ!�AHka %=�j���z�Y.[�|�{6�~f��ڗj�
�H/a̤�$\��en��IپѮ�! ��
As�2�OX�QퟜeJ�#���Sde���*����<�*דe��dd{�$-!0|�����ؚ�j�Y��d��WKuGX��tr���F�y��>��EX�9���K�U�r�h+d�q�j������x��e�:�!�zF\,���V�P��9u	֌��!mQAO)X6�>�'�iJz�}R�����@�	���@o�-�#�	�j�m��(�i���2㊚��@J���G �8�Jz�-�Ee)��'U�8�s"�K�$+�Y�jP;�R���H����%�6�*l���)k��<|YA�)E��-zRI�%�B0Տ�t*�S�X?bvʌ{�.�ӤU�C�T%=��a`��ӣ�|NI��,�Cq�4g���m������)�'�-%������yM�Z����$W ��gĜ�QO�!!U�:�	��=��s�|�XV��0uT&U��_R\�G���)�г�F�	�A���aD�L0唝C�/�秽	��<x��E$���D����j�� PL�,�E$�&J�D��0 My֌�"��E�h��,�*d����X.�;Iݜ��J��k�i�a70��\�T�6��>MY��	 <�D���!�/���e!�Є����=���{f�t���'l�c�.
��I��,$�G�P}O���hr+&�~Nn��n`����i��פP�f�b����jt}O*	�L�,^���ԓЛ%��I�� N ��P������ ����e�� �p�L�*t�����N\240����=�����z�����^�$6,7\�d����V���0�{�=V�g�YW��Ɉ��-���Y�y �K�U���dPt1D4�;`����DO�讑�HXmޝ��5{�������?wh��>&��x|��������G^���*K.I��K�t��������4�:dP����H���H�#T ��{�JIǫ�S~%y������ h�/��\+]��ܓ\�Z�R��x)���"���D��c�����U�hϵ*:u�I���"x#^�������i(�ʽ���v{c:��C�-F��Z�I�����YF����7C�ܓP>'(�6�KK��V���rNbk������(�V	hH�ؙ�� xG���'vҩ'3����>�@J�xuJ��]�ͰObe~9�N<W�M�|6hDrR�r#����f�5�(=i��$N �t�HQ�o���M^�j�#�*_��õc/�A��)����O.(���� H3?��t�x���4�<	8�G���+�$\���f�̌_�R���r�p�9�?BA�7�F�T9^�2g�)��'�Hs��HL���8A�� ��ۚ零,גe䋤��61��taF伂�3g�������ʜ��o�z��V�F�7+�n��.3s���K��]�|�J��Ѝ�8�;��q�/RYDG�QE/�u*�Z5L�g��t�Ϗ ���,7͜���'��Z�x����r�.+`�ĩ�n��Q� !�UH&o<��7'�4�U�+��kԊ���@�T��eF�����^+h5�!�;^���{�X�C��C��� 9�ίݑ���@�4��u��Y�9��+H/�&�nq�2�	�ȯu�d1��+9�M�l=7�)xh�T8��M���>a
E*���b����
�IhWn�E��j$S���o�.�K�+��X�R��
 ��"e4���ר���?�"��I8O��+DՉ�Aa��'�:�zI%d����ݞ�ys��[--���^ؓ�Y�\�D/H�DR������b?~0I�ϓ����C�k%���Q��y)�z^���!E�Γ�%�$t�xYD+oR�@f�P{�y�!?�%��t{*'c��%g�[�t ��n e�������O�I�dA�G�xe~A�Z�~0Lt�H�����ێpL���T��*��y��`B~9V�`�y|b���<�E�k/��כ�je.�y�Yo���qs��j��
I3�I���y������g��z}`)=%�y�������R��/a�[-��� )� S���]�k�>�_/�f�	@f��Y�0T�5�T��@�ԯA���,�K�t�5�<���;o��̸�6��Ht��r��Z�]�Ԇn�3^s(�Z�(Ȭhu�s^�_���w� Y���cO��10	�)�[�)�7r~0�% D ������A-��)��L=��0��n\x���@�5�)>µ$bk �6d��Y0�	r�y8R�\�<bFK�ޜ�U�[`F�@:�8�!����pR{�����GÌ���	�H�<o�a�h8X�d�4>��aA��y���*����!�����F6�*�y�0ٗ�cH���Z���a�n�$O�g1�����P�D�j����Ѓ��7���"��{$a����6b��-0���2�;fȨr����cz��@fao@�1M+��9�[�V+�z#��6��b����O���0ئ��	2�L�4�g���0�KY��GHNI��[�0o/�p��yxeP6La�#$���pł#��@	£�z1��}��ȴ��ĆxН�a8%�~�Ȕñ 'h?n�0nһ�i�:Sx�2��@r;�!R#�a8��c */I�a=o�a����Mʤ�k�ƹ����0�),�f���խ�Kg޽�.����<��X�v�#� o&<o�a�~�
��o=)�q#���r  ����E�"<�'2����rވa�kK�Dz?)�=��@Hʻ
J�6-��T�⁴<�J�x,"�p�Ap
>fa�J�q#�4Ͳ�aCʺ=�ټ|#�����D��*#�F{���2�w
 U87Z�_o�0�|����7S�,�mHD5U<�Z�CNJ���a���y^)����SE�04���
�~�>:�y��a�=�,�l�y��H�b�<����d�tg�������^��0��>���a��� ��ԍ+-�����މ	XH�T ��ވa�+B7��@B�r9Ȉa�o� �ӤB�����g�ܬ�,t���(1t@z�����Ւ
��>Ȉa��ZRp�*S���1�D����o��/��LF��5`p�������`��JŞ�м"��T;��rO���@d�0�����
#�u�[`	�*�*�I+�<VFC�-�@��W�,�Sd{��^s�C9o�a0�I�$G�y��?��a(���i�f� ��a$!.H�2�|<>��H�_A�*0�1�:���'Dw��"�A���R��{�,#���)yH+�a>���H�.���9I�L��"b��0.`uX}�Ï1ZC�����=�����:tCLR��T~àU��
�WF��v1�A5`�q%|R�HJ��,��4-�v�y3r
8���W�o�a��PI�,ر�F��e�I�:S)���Ak���2:�"��-0Z�<�D�g��sSà�����������yC�}_cR��>���|MAE��>H(`�i�k*b���_Ae�O�gY�&�"��O��@���1���BE��)x�R��ރS�������x��OY�:ӾN�"�Q���p�W�l<o�aEw/>D@�;�U��8*bEy��K�t1�x#�Q��^ri�~�=o�a,(���8��vz=�F�~�!�T��G��y��Tg����0
��?'��Ǩ�6#��v��/����/߈aa]0�B���X1�,0hHj�*b���^��@�P�R�`��0h܊���a�~�O��\�n��>1��9��t9�y��(k���7S*6{���е��`�' ���#��pm~o`��`0�sH1�Ί���{Aj�uRGC��Ҥޤ1��8UGC����T�����a4}7U`p1'��up1r���K�ky����g:b�|*��^$�uC~� /1Lx�����g:b�qo�#�q)�;�h�>^5�i�b�3���a�^�Oa)�
$�g�7bL!y �GP�i��-bL�|��y� H���1�PޭhE�<I�sވah
xU��Q��c1C�FS�ɏ��w�1�~R�TC�1KG�)����ݐ�r���a�<��C87#��/t�0T����i±y��#��!�j��?��M�wL�0�>���[�U�L�0hUAa(��Wf�^J��0huO�2Q��U��(B𴆊$���+ӷ�x]7�P�wx����t'�-0�zC7��0��y1�f��>��I+<^7�P��;�$�{�D��"��V$���SP�e1�c�Fp�H��&b�
�4�
�M�P���-b�J_7d��|�Dcx�쀀����j=~�à5�����p ��^'M�0��K����㐉*lP�d��&b�߇�TW�����>U�ݕ�a��W.�u���;��F�1 ���&b0J�@NH��xC���� �I��}��Dc�{����k�����DCu�`8�Ӡ}�a�
*�=�F�c|��D���zhv:�q�0����w����R�ve#�!��^+��QXl�-0dX:�V�[�AFxc�1e�!y T�9[��)|�l҄q��ue1��/��l�O����xa#�J�>�b���EK�Ҭ�-0�ʐgY��#?�Kp���06sϸs�4�4��h#���4l��C�|l������\�#97�y��A$�BH�y��t���җ���s�P?e>^f���}/,�y?��S��>Y��
Q����-0��Jc�P��;��[l�0�A�0�^�2��8��X�ҍ��B��7�I1��YAH#U�Fj#���c���.Hӕ�-0�h��?�q���ECu��7v�����ك�MgA|���6b��p���0N*�-bk�2=�N8Һ�Q�[`K���y+?�Y6��.Z���k��պ�3^�N��� V�Q(&�[   	pHYs  %  %IR$�   �eXIfII*     (           >       F   i�    N       %     %      �    �  �       ��    x       ASCII   Screenshot�M_  �iTXtXML:com.adobe.xmp     <x:xmpmeta xmlns:x="adobe:ns:meta/" x:xmptk="XMP Core 6.0.0">
   <rdf:RDF xmlns:rdf="http://www.w3.org/1999/02/22-rdf-syntax-ns#">
      <rdf:Description rdf:about=""
            xmlns:exif="http://ns.adobe.com/exif/1.0/">
         <exif:PixelYDimension>512</exif:PixelYDimension>
         <exif:PixelXDimension>960</exif:PixelXDimension>
         <exif:UserComment>Screenshot</exif:UserComment>
      </rdf:Description>
   </rdf:RDF>
</x:xmpmeta>
ǃۥ   �IDATx��\	��U�������N'ݝ����$��%�T�PAk(PK�-���*GgpFf�aTD0��R�Ț�HBBHgOw:I��}{���~����~M`�)o��{�/��{��{�����t�jAAAzǆ�?4�@��?s�O�q�L&������gn�5m��sz^?��\O$�=��'��s�����'�d>�,[(��q�`08��T*�u]���7�5�\�iӦy���~������v�y��H��o��cǎy�幻��۶���aT����:�7���32����B,Zt�0<<�M.�����B�4�a||\��|QQ������&�_p�8u�֮]�s�Ρ���V���ӧ166���y�B*((�&ǃ����b�ܹ�7'����̙3q��Y���L��=uuuH$(/+GWW�ܯ
�O���Ba�K�,�/~�����X�����8�u�%��<_|�E���t�r�-&�������X�j�b�;~����:000`�J����h�՘={zzz�x2g� %�%�D"����A�2������
��ىy�������R\\,DUWWcŊX�f-��(JJJ�
���F�I�����w�Ʒ��-���/��1x��سg�����BۓO>�O�Ә:u*����V棖��de�
�t�9sFh��-ƶ��bW�&���ϗy���k��1�u����bp�����A$�%Z�~z{�L�~<x�xVD�Rs��t������.�;v������o߾]����::�+��If����d������,J�O�8���n
��¢B$I��7�o�^^^.�w��Q��_�r%v���Y�g\�O�ʃ��5u��]�VN���������t�2�y�
Lݪx���h�$?֮�(g!���'6b���¤X,!D�#j	�U�PɳQ0����B��5�~��{��7�0 f��0_شɋ#�4�v1T�_���b]�,��@ȇ�Hf���f>�hѢ��E+����ɜC���3�I�x�7���o��}ٱL,��~�i<��S2�
���=���1}L�>M0c�����w?-�9��۷�6�#���a%�&N�
���@o�!�5kֈ[���a���v��!<���^?�
�鋷.ǚ�����#�UH�"�6P�]���˖���_�y5��)�<�G[F�hQFΚ5K�e�T@��D��~i����^l��|&wnڟ}�rh �gWw�0�q���C�'MP��9Gc�L�c�1��|�����$�82�~�҉�����8z�o,�Au���}�1�ܼ/n����l�^g���sB>�Q�WlX��Wcxh.������\���<H�@���ac|���%�M���O��Mz���?�;���:�o�Az����^v��98AL�x�`�21_2�Ea{M >d܅������%̇�����Ţ���9?0��m��ju6>�㩩(4�DM��ѓ��`��-�1�z>g�����|�U����V�k<"p8p� ֭[' C��O�{f�9���L��z��p+
�!	����� ��j�+�� v����iB�=p�]�Hl]��Ʉi�Rg#57��=ބ������Y[/y�e>4e7B�~�A?��CQqQM�'�'��ߌKD�!l����e�����'�4��1Do��tu���0r1I�Dk�$ɴu"�,��D�	w[�3��8�������g3�9^\Җ��+)�$7^���j�#O��X4�W^yE܊���DP�Y�h�J��W0��?Մ���G��GQ?�$��>.��Ȑ�pl2��n�(��/��b�m{Q���I������g��>p��xv�sު �߶�!�D7v�u71u�E�	��� �}f1z;�����+;�m�^�$U�S�Px^�~s��6���8��_��|doV��x��ۆ̴
�ߧL�2!�رǞ��6�5Q8Y9K3���.K&Ƨ,��@f�W^yeTd#�$𪫮��ի=A�.����w�ox(���a��x�h�)�j�qT��y�nm�֝X�0uxk�Q?'f���p�Hu��b6�}�jj��~饗T7W�`��{߇@\8:�}@����MO�>]a��Y�Ї��,��j���^"����D�H�d�?���Ϳ��[(()����j\{�����;���M����@�$�ј�$�!�.o��$�	���gz����r���}�>��	�ߧ@��[a����aU�֥��+�����	��=�h�|���Io۶M�}�Oki�n�L��n�,�ZQ��61LǾ}���+�r�q=<�`��9�t���g���Ͽtܸ��Qie������f�l�N��xOn~e��{o��������"��djM���a�9S+\M�!n��������:}&ۧ��2Cx�͹-;�0����$�����K3�XZU)�z�j�#��`�5xm7��
J#0q-�I�;����������E��V?���*[ vF��$��lү55>K7<{��,����v���7�|���^{�*�4!p�<���b��u8��chinFc�l�r�mR�y�Gp��1���0~��lz�}����y�����ؔx���s;�9���m7>y*��ق���Rn�ð�x@���JG����g����΄�j���L$CI�&�.�<�Q�y]-��U����ddkk�7�,���aDg���2�g|�'>T�Ջ��68��Mg\&�(**1�A��N(O���_�a:�����i-��)���4ݢ���u�E���U��ш���7���������K�d�bè�$�Z8t�gH �[5���<����YT����0BE4U�5m޼Y\�M�*���>�g���?x��	�5
�Z�9�4��
�8��X���S���R��B��y ��Bg�����m)�2�DabZ�@�����B=�Z��r�W���tP�k!�ģ\e��Ć���a���鐱���L�wcZ(@0��?M2�:��Q�d2��!�Ak1چ�E�[��Cx�u�|i��&~D�lncc�T��W����:?4�f�$)�9L�>f�*�xѪ��:{����A'02r���
��+82�%��船WQ�O|�1��]�V���ۢ�Q(�'7��W3�)���D��p7ݰ���w8�w���9�d�����֋p�g�=h�Ap�
���qY���s!_Y%_ˮ�ϒ��?��e�ҥh6�^�ڕ�����D]��x����)Y(�Z��������O������ѣC8��i�D�9iz&�=���MN���	�Qa��hYKK~����t��	|��_�*)�w�}76n�(��I"Wm���U�n����\47\Y�����P�3$`bJe!n�v
���[�;bY�$�{衇�*�]�,�'j>��(���W��9?��3f���s3
�Ѯx����]1|�.,,BIq�x'�+*�|6,���Ѥ%S����-T��HG��8ۑt+K����p�����t)�U�뮻��C�7���m�M�������w�2ֈ�����%2�䔸=�&g��3�
�y8N6x��i�̪�瞬dӶ^�z��/�Kɛ�)�!,f�&�E��kL��}n�#�.g|'O�0�tA[)��vva_S�1�"�E����G�벺����sg0v\��U��
r��/�aI�Uq�^6��B$}��qajV�i�!t0��CO��_?_���1����[-4��'���{�0ٸ9èT,%
���EN��FX�_~���ҩ���^�ü�LVz���+,Z�w�!K�t���Pҭ>�K���v�'Lf]��݌�?3k��၍�����8��_"a3����z���a����x�s�Kq̣���>��0��|y��jkV֠w����b�fWP�ۿ`�&�ch$h�(7HPs��#���#�0^N�4#L&���$Q"ذsZ�����ȑ#�b[��\�T��4�ֵ��I��	�@�gE���q��A.���z�_� ��J�V 2A�h�P���w)I��C�?�k�p8��hJ��0����_�F��S�LpO���'��3#�_�'�܀Ϧ�{�ĚL�D��Йֺ��9FV��n��׿�)z2a%3S�uq&�� �n*7��A�����yo�C�0C\�<��pg���d��
J=`�?5�<�����ȏ�Zc����1��V�U� ��jԚ�b��Z��Ԏ�~�d�ɀ�����Xh�./jb��~sc�=F�����������z�~^}yJ���>+��ɡ��s��t����A�;��.� &|DQ��h�册�~�S�c�/���EA�~�\����L�k�|� ��g;��A��tF]f|H����Sb�)�L�O���n���T����Mt���w�Y��;ObŲ
������qB)##O�%h6�Zh uv�I/K�ۆZ��6d�.����)�Ux-F�����m�7�p����g����>	�H�ןk?'~�qf�aNãC��KJ��4::&��
�`c�%h�њ��Rc=�dB�0�/�pK�0\!����^�JJ)e��#+��s��.�ӏk �ul�_׿m�1�p�A2��y�X*$��d>!���&�~�j-I�9��<\zx���y�5*:�

!ܪ3ݸ����ը�*���[\�4�(śMq=�!(�{�FFG$δwv���u�g`Պy��*t�'���w�=�&�PW����ńŅ��CG����:䷪�'M��8��\."S��u*b��r��r�eV)��ta����(K�ٛ�E��йE���s\O���1�SW0j��ͻ��
���
}�~�C��q���X��m�a8�.JN�.�*����k����p�T������q?k]TCI��_X�w�b���9�����:��ɂ�z]ݚ����)縟nq5 ���,*�y;��B�����˲�|��Mt)x�@���4� ��8�p7��
� _�C�a��``8᭮�;���D�f��İ�`m�,􅔇�leW?�	��0Q=�$��(��BH������7mͬRj��u��.�~�[˱Q�pc�l.P �y5]�bX���a��6��/����|��	!�q�&�������P\Tl�Q㦆�?`���O�+@W��(�C�q��7�����{������v�Y�b�����.:�Z���>�J���7��R�͠�8&�W?>;'��5z<�bF���T&�Ln4�;J�/����{Yjb�A!��dǱ\T�����gcf~W;S�}c���X�`�� ?�O�������c�O��٘p���a/�Vg՗�럛�ç�x�E���p��ϙC,a�i���쐉S�:k�pA��Q��Z����s���5�h�4<��0v�9!A�Bi�U����B�����@���m%l��t��R��;x�Q�Z�ޟ�a�1[8y�.]�B�$q���A*0�a�L[���r3�^t����BrkYNV��o�1}�22��J�2���xg�0�U �W�������gP^��I����o���:��颕�0�%�ĺ ^�c�����8K`Jy��G�ĤD��x���Z}�L�����Ʀt���J?F���ߟ�8��A���-��W[m���<�C7UZRlbKe=�����F?5�p{J�ƽ��dI����}Q<��۸���*Jw����\w�u^ �&Zf�ݶm+�y��n�N 2�d��C��	�c�Ḟs�'�n��w�G����4�.���,�s�8�N.���z����Qok+���~�Nى��L\�˦=�=h:zw�25U�8�Vn��
/�������[)����-6�2��߸��Z}x�u���K�)N����g>3�w(r�阬�{�}F���?�?bd8&�e� H�r����K`�aI��1��pu�����}k���t1��ϵ�|�� m��\�;����}�̕5�-[���L�a��1�;f�׃�=dLޏ��s�2D�����0��EgV�R�,7���1]��p�1�z�-Y�L��i�,�	���^P�d�7+_H[
�C�Ns�.������`6c��>����ڴ�7p��QL�H�/����EU'Gv�!�֮�h1ty��{�m�F�r;�%Z�����@��\����Ĝ��8r����S**+0��5�S�t���m+�I�����	3Q�a�=�0FW�l�L�L��D5�@�홥]�Vyy&�I�	\dY�P'U	2���
����'v�wz��\�Z	�����༘�0��*�D��.��2Cv�[;�;��2/�c]]�x|�⻙��zo_�r���i�S��|)�!�&>Y˝����\����]d���'w��$�N�\��jD�lX���ß�nŉS��{iu�b����$�Ӛ��d2����5�=���&���݌�P����\�k��]�r�2X��Xt�$2̜���D�=��u�o+��N��F�BR�]�,<��|�te<A��M���%8�ҎO^���2�TvE�M_lUz�5�բi�\	d�P��V�/�B�8�<H���B ��|V������G�[��o�N}���x���N�v�\V8�v��v̩�!o8�%.K_�ɥ�F��ݹ�$>�f.��q��˘ݝ��M'_a ���5v2�������3W��n��c�f����4��O~2��%Sw�A-�9�ϵw�S���r�iQ =�����v���P��m��$aB��/ǖm-�ދ�&�9��Ս�.Y!cI��Ὄ����9s�d=k�>;w�\�2�	�2'�.@F�g&Lk�K��E�k�S���a�Aw�eř<)h�`bd����\�9
��4r��M+�Zۢ�[Jm:����N�6�f�'�i�s�҉.ۚ	|�ߔzЦM�$;�ݘ���ԭS���Bg� �_���#j�b�e�=���mݺC�@UV�^������0������"x�J��qE-?��#¤P�wJ&l%�A�n��ß�t���O��/6���^sw��׾x	�^X�M/��L9v��#�J�IZn���p�J̚Q��ol���r<���ز��DJ-�ګ��n-$�����I���R*@����o6O Z��E�L��ƹ����$�o�w��f-��V[��rsn	-*`������uwP*���`;��Z�0p|���"���uxu�)d튱�����b�DI��m�c�Q�T��3��(.'O�����6/��Aj��Vgr��	܂����|B^+�	�p�wr�������Rs�,��F�c��+�ڧ�8�]�
R�౧�����W�P]��ġ�G
��X�*S\ar'b^~m'b�3�|�4<�����s{|��eI�Ua��w
��,_�<�*�Α	1��]�*O �;���7|��-D_?^~�%	�'�����ӟ��<��vQ�Q jv4a4n {/+!3�;'��z�|��E�s�M7�������jr�L&?p��׏��;�z��O�8��豱QÜ~<�\7�eHIUY�i�Ej���M��_6RQi��B�+�޸)���̟ہ���̑������)(,.ü��y{7�G��\����~W$K���}�{T�i~:�����Oh7M���.q��VBەil��W\!Ȍ飢�.���y�slT�uk�I6� �iz�INS˥�(J�N�#MJ/w6�T*�,��B�;�m}G1��$�{����1���Ƞ���~1�ܷ~��^���08aN�hAw�s�C�y�k$����~�-7�V��G�{}�Z�	ҷ�)��;��Z�����uj{�&Ҭp��7�K�;睫L��%��ubt��O��\�56:&u����6��B�S��`~�d9I��uх�Tb���n���2��i��{?�V�m�v��ǅ�wj+ĭ6Q�����y*�
VH���R6���0w��+Ԗ�T����d����`͌rY:}���seͯ��[�� O�z��c�&������K���K-��ӟӨ,��[�V�@�A��c�֭���JB�`�b�M�ƠOxLKџmR���*�'1ߞ� ���\a;�LpxpTV�r�0E=�{�D�v>5�s�_�AWIw�_m���jt���񂮖`�ej:��+����m�W����O	�� &�|ހ��H�tj"�D����E��v��������v>�z��e�7���ͽN(J�P+�
i^x���J��gP���&?}����8����,��/�ʽv�9�j��!�4O�t��X*u��T    IEND�B`�PK
     mdZ?�>�oH  oH  /   images/a038ca8d-f9eb-4e93-ad0b-b831193aa106.png�PNG

   IHDR   �  c   ��T   	pHYs  �  ��+   tEXtSoftware Adobe ImageReadyq�e<  G�IDATx��{�W}篌�-͐�_�K<aF�	�!���2��,�v��?vON<J��s��X!�c�l��q�g7ɑΆ�eA4�+a$LV^�0Y4��H`$�&X�H[�����.UU���n�����>��3�]Su?������BCi
C�
C�
C�
C��Da^���|y�!�3���̙�D_L�0�h�\�}�)!
(!
(!
(!
��,_�<|R����G�4%���wB��Ȉq+!��!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!DAi�Y����s���fj�H�U����?�[�I"���ĉfd�n�u�CH��R0::j-H��V�q�&���!YQJa֬2;w�2���aj�UnHV�R�͛7�� �f�����*�rH�A�ƍ͞={!�RJa�=j�l�b����W<�	@H+�R����wlxx8hÌ��mڴ1xmY�c3��QJa4�w��t4|pl��J��۷oG�t ���B�����n2�c3��BH3�^�c�vs�u�����B�t�0�f�،t �-344� ��#�v ��7m��o��1� � ���:�>��]��F�(a����%1��u�������k���Q�[��aZ��ߐ����pWؽ��{fH�t�0 ]�2���h�Ha ��H �!�:V���AL�gi��T�fvQ�0-F����{��F(�0(�)4��1Eƾ}�3�I�����ne�(���<�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�((�0X�k,W�����`���^n�����tQ٧�F��w�����4<e3��Hye��A
�ym�U�STJ��H�&�^�ϲm�h�wM��a�>\d���Y̝����-C4��`����300h6l.|�TXap�$�t�fɒ�ٯKj^?|���׉��ƾ�X���ā ���U@rn��ǎ�cǏ��V�j������{�k$����WD
'
����cEY�x�Y�r�Y��>Od�G�O��2�'&̾}����7���`����6.�b��P��K���ua�}����̓�
��Zs�e����|�>�!H��#x@lzU��z#�<�DB-e��s�����n[{!��j��A��c����G��`���_ֽep^e�i�װ�D�8P��<�,`������W�B�4�f����3\!�A���\u^���ݾH� ���3\\��S���}�RfwI1G%�jխ�E��s�h$2�Z�H�;|��L�~�����T>U�*#$���'N��wܑ�v� �=�]��c�\ǲh����e������Nmq>Q��(6"F\[�R�����Ê�DqTFG�N������ka�dA-�SSS�,aڶh�yx��c�1Y��󊨂��L��N��hHm���5\��=掠2�h��lz�f�#����]ԏ��������@�{�/����mՂdK���
����Ƶ_ B���$�o��!���c�S��p^}�Ka$��M�o�H�v���ip�����J�mHIҰ�)�4��u�/��v� K��Eژ	���8��V�/������эtD�A��}�N4 �Z*�o?d��A:pq1��{ר���~9�_nQ�?��9eօo)�W��X��4�ѮJW ��,�!M\\���Eͽ|�oS3���WT��^�z�w�=���
�<I}���+a��H~����P���g�\�z� �G׮�^\H_�\��z�m�4���Z �!*�����Ho�MvqjY "Ktl'N��SB R'�<�I헃&N��Ge
�{lڴ���aO�@Z�G��YY�5��]m�`ִoQ�>�(�Y�׸�KҨ�H- ���}� �B�b/DC�Z�E����pa}�Վ.��^���g�~�Ad�y�{�(�����=yD��d8�mAZ&m�jC���Θ�LT�m�$��i���0h� ��!��B�))dyQ��R�+5qq}Ǝ.�o�8�$�_*�aZm'-���@>e�4ۍ'�̥c���
� �'"�T������~Y�Q\$A�A{n�-�\�[�� �@~
cL��r��f #e��c��,@jTI�PP�=1���X�����~�o-���e�޶c��EeAdA�1�,e�~��0�yͪ I�D���~ �=��k��|�J�ŋg��"ұ��SY��+$¤�3�v����&E������JԾ�ㅱW�5a^��+���RX�2�Ğ��}:v~���t�f��2&s��I�n�.�+�d]([�6rg��ƶ_&�m�vE499a�Mۅ�/lVS6�]�w�4_��d9�(����Ʈ�a�9�^�ViT|��:@��I�%��0�Iۅ��x��W+�M=Y0QRd�ws�'����t���va��*=:ǎ�&�,�'n��"ei���K�=d�^��.LV ��Ŭ,>w�,��v�,�]X;r��"�Mj��2��G�����`������e� n�k#��x�!�/�r���#wV2ǵ_��Ο���=W}���m��������c��Ap�ȑ�s�=�n����č�n�0�D��,B�j�i�"��ݗ#�2�B���l��}���Oaj
ױ�{,ɷ}�EF��l&�n��*#� ��mYM��>nDL�3.���}��0>�R��}��v�l'��L���r�Q\�%���QЙ ,�d�/��""̾���u��-Q|�ȝ� ���
��t�&���[�va��kn������|�ap�"n���j���w��s�tl`��NpÕ�u�s���pR�%���6�����1^�����>�{�y��b��pK�������\T�>�hZ�cmf�\R���t~�>�>�i)x!���"j3H �iB�S|�ܫ!��o����$@t�l�$ĥ^����yEe���;ʠ���|��e��"~ ������Hw�6�D3V���~q4�����0 ��ls�s�P��&�g�9668��-[��ۇ T@v�n�����t~�ϫW &A�*�5�*&q�c�7��U�%
�Vx��<��-Z�PaOJ�\L��u���z%�IB�t3c�%�d��RD��I`����a� ��w_C�/.�r1FvO�%��y�N�g�C�櫸�(�󃋊�ݲD/*z����jj�Wl�d��z�1���Q��^�}�>�08a�D�b�'����7AVYV�qϞ=��T,
j�;�W{��&n�%���r�y�yD/�C����t�2��,0����pe��!ݕ�Hصkׇ��D�4q�,��K�`����y�V���b�-�Dp�R�1M(�,�Ȯ��pO�I����Ep�~�t8�v_�0_�%�0@�A��=���V�8눃����]s��)M�e�-��Kz���E�[�֮�]<n�Xk����-(R%�0 '�СC�^��5��h�ɚ�-��8I� �f�.P��H�Еo�Z������A���Ks��ej�=�QY�r^!�F6��� Bf,�8����k�gw�=Ԭq���'��~��,(����G��h@΅�̬v:?�+"���DJ�C�蒷)�0
.v,F��l�k��,:�#���f�E���k�����W�Ư(�������]���?�h8��^�Y�xͶǎUV�YT�I m�miw�b�F��x^'���nwق8����ֆ�۞Q 
ҕ�f����|8�����Һ�'챴�o�K�S7��PHa��(0.9��R\l�^"((x���+A��U�|`�<��%�k��X�^����*���ސk�&Ƀ���.�wc���'��k��G�:��w�[����Oi��""����X��XB\@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ@aQ�fdd$|҉0�����@-�[o6o�m����y�^`.��#����W<^y�<s�ET�y�K��x\p�)��y��k����r�gf�9=sּ4sμt�\�\g����_<sּ8y|��f��>��a0����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������8��_=h=?P�����I#���xײ�߿��K���/�2׿�/|� x�淾͐l�0J���o�S�N�'�9i��ߟ<i���Q�T�Ț�@ڟ����1W��'���@��]����u��g�q(L(�O�����
��ȃ��c��ϝ�sH���;�fKC����sr>/Dx�[�"�?�o�_�QX1�Q<����
� ��P7�{�y�[ V��d:N�/���"H�H<�����=�kQ�:-�Z�5 EU�ٚ�4O�D�����2G��	��/|���R:<��?������i�Dᅩ�V����%�#*R�_[��P����]Ha$�<����@/"�L���u�}
!�"���_�<�"h��kY��mo��%�; �ߞO��� ������x'ҭ�|��(I�k.�}�o}�*�Ox!�����t� �<����w��E�Aۄ�;�-�;I�N��a��?F���4.wa�r�fAź��	�:��䝲�"�������O���>FBZE�;�4��C1�y��W_y���u*��?<j�T(!.@Թ���>�կ�ܶ�w�/����>ω0��O��?���{�����/~>|,��uf��������4�rA����0?{���g����/�ϞgOiǟ����;~�\:���ο7�>�!��5Wg��-s�GO��O~�<��݆�xṓ����>�[���C��4-�S�|�L}�3��2��΁�*|�aɻ���l4���w6�>ja~:�������O|�R4�s�����}�4���?P��Z��=b):ߛ�Z�x���N/���.~��)��SBPBPBP�6���g�������qC��i��˗�_������o�>�&2��.9z������~?99iN�89�|�z��O�� FE��\����>9	���hU*F�t(L@o/
[o����5�lD��$JA&<�X�N�	���fY�nCt"S\�B�<xLLT�v�F��W<�)�>8���(A��KT*aD��c#GNH�444T}���Z�vQ���A�ש��OZ?��J��fI�x���URήԿq�\$�+�_my��
%���"�Zz��\.�]��B_s��;V��my�W����\,����@��;�b
�0�pk�'{0�^+��V�|-��k[�����V�Z�(�
�k�cػwoC��/����� ��Ep!$U�X��@���\7|U�f:V�wh������By�Nx6��0R�Tҭ�R-�8�7��( O�#�?���1-\{�G�{llo�Y>\϶	cK"��Q¥�Rr����(�x�"I��20��P;�N�p�GGG��m���]I��.�4��Q�.�NB�L��'�i�ҳ����ۃ�\�ٹs�ɓ\�Am2<<�Pý���9O"l����D�-[��m�m�Fs)+΄�����^�C��Zu6RaJ���-�����
v�G�n׮]��Q���B7pR!P>�~��!�1T��<ߺuK��4.��3�l޼���K��+��c�����IB����I�A�C��U�iI�M���i���h"��>u���@(�sӥ*!�l�|W(z�Z)�M	��B4��.�Y8�l��vR���Um!MC���4RV��qU	ca*���7���Q���t"���T�����y�f\�Q�҈����V���R4��G:�S��� �a<$�"B\cw �@�zѦ�0l��N@���Ëɗ�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�
C�������==���p��b"�
��-���54%LWWw��E�1�������ܭ������ �Չ�"�k�N��4%B���)�֢����n�c�Z
C����"� �X�Cmt�dB|Gv�n�����+��7B4`�fQ�.A���h�0�h`#c�.ύ���J��Bh�暄�����]S�A->��I,z�()
vW26�Ey��TV�00v�vC��`8��%ۍ��59JS�8 9�F�� �v����G A�Ҳ��x��W���M���2Dm>HH^`�err�����`S�Ӵ0gv����G�����e����.�.9N�!>c��m��\:Z��s�0-#~�T��h��ݒ0L�H�ӱf�^lZ�E�i�{*L��}�ea����2-M���pL�x�=���td�j���!�Q�����1��0�|i�e�[F| :X��$�L���-�A"U#���Jhe��&����/_V�Ȇ0�UeH���/�ʂ̄A~(�p�0��L����L��)� �ĖE��gAf ���F�1I����,��t1r�!>`��c�#+2�e�^&��{tRY�y�ؽLڅ����e9U+��ae��2
C�v:Lv��\D[�f�&�Yj�٥c��0&b�'�_�]3/sa$g�4�\u'N����ɰC������Cڂ��pa{z5!.A�n���l	3
�p^���)����0 �Hx����0�9v6�����L.��+o[&�q��΄�g;��]�\��:M��PF\�v2�B�A�E00�K�N\��L`�c(qI�p*��S�٩�-v�慎8�R��[�7=:]}�r�yJ&������e�܄���\��d����Y��
�d�ե��3A����������)qI^��!��M�gOqA�R2��{���$_��twwU��]�dE^����0�{c���\��:pNq���t�yJ�c�)��MBZ%a\��0蹐�v-�,ɳK�"�=�t��ICHV䝱�Ԇ��)���0�dE��/�%�6��C�Ln�d�bH�Ԏ��:���#�b�+�X�+aqA;�(r]�]FٵLZ%�)1Bn k��qE^7&2%#DAn��.{�)i{�q����	�{��K\ߚ,�&%[�f��'h�oܸ����b�5�<�܄�����-;yϟ�����!~�s/e���5R��l�y楋��'gf�ks&������~�%(�0ga�\t�!~23/�ESx�#��a|�)ǵ)�03/3�cfΕ�ڴe���dg���҅�(e$lÔ�\G��Lg���K�㢔�3%�4�I�΢�m~o����+���/�0�F���䪔Fπ0�0�Ba<�dg苷�aJ�3���4�W(�g��~�R����VsIׂ����j�䕯}�y��_/|�%�kg~���ُ~l~����k��H�_�5�VvsQ~�mo1^wM��������k�1�����%�b�Ht��w�SG`�z�k��~`|f��/�yn�
jǙs��>���_}����_�|���x�y���9��%*"]���_c����ɿ���3��aLn�����]9�0�(�gg���ް���k�����}��_3?�淪���~�\yCE��_�]r��ξ/a�Qbo|�b��vg�"$pYS^u�s9d�������n����0�gN=g��w���o=a�>��\Ȃ����w�O��o�hôc��df���|�ܹ�\}ƅ�\l�y�M��@���1/<��y�D9���~ȼ��~8�~���g~�;��8m|�E�i�6*%&h_8z�6��ϸ��Ef�ŗ��3���9��3�-~w�_7׾��{t�u�'�e�~�y�{+�� �+���\��M��W���<h=3�=��c������d�Qi�8J��6L�]}�k��,����	�����o���n���G�f�UW��=�������P m���w���,1�^��_}��˩S�3��H�y����Ϧd�>�+���������M����di����p��N���%�a;��?7?���B1^�`����7�?� H	�[��L|����;K�Z�<7a��\�RFGQ���K��3^1A��_8y���8��g̥�_^y� E�}��T�X�z�㗿lΜ��A4{��;|~��_����0��.nJ�#7a�F��U
ݶa�
���X�`N�炚������� C�^=nt$��t�6z��Ϙg����WU�4H�~��S&k��y�qհ#��s�aw[#�l�3Ά)��{�}�y:H�N������0��fƸ���W�:�,r��#�L�a�����>�l��F�����[�ϳ��sI[�0..�6�9ㄚ6����IP���/��˛����޳����ӗ��3�����8��=۱�}[R2{򬨤dn�S&�1�/���ʠ-3?(��~�/\uUx�?�=m����Nzߙ��h� �q-Q�R2GƮ�]}����=�~���L��W�m�dy�ŗ��y<�ۗf#�\�8�x�g����8��![��%��1mI�\�S.#����N�q��41i�{[%U}��%(��U��/�gi��ib�)��N�0��^+�:oy�e��%;�np�}��l�Sϝ2���?�׿�M�� ���7����#��;���
�/8����g�_���;����ߌ���J��'`�"��AKPi����3ƚ|��3��G�+���\|�Ŧ�oR���c�ߜN����K�M���\}����;}�����G��x�:nD��c��'��sN�G�q�5yO��E���jk5��d�u��l�3nR�W͎�?�7��W���������_0��bsE �o|�*�ԓO����*�.�9��,WC�@�p=�O��sҚ=�c?c�^ZoZ+��6v���qM��Epچ1V���ߠK�5W�6
ҩ�}�S�]+V����_4�}��G8��?|:�,��B	3�q�������<�5n�]��4f����w�g�9�0�q�f�F@����φQ��o�3�"M��{��ߘ�Og�c�7ckQ�a��E��a�B���A����z����(O"<=+ë�F=�/�6�O�lC���i��{���C�p����z��(m�0ُ�sa�֔�g��/���8�6�H���0E�eOY�0n��Q����"��Rt$�0��1�����0�0g)���8��P�d�%*���g��\{��10S����Z\oE�\{=2Wc0���%i�)�}祽��S������9k���Mooo����bJ���e�k\Vf==��
YM����!%��>w�O����@�l�q|i��H�<11Y\a�J�a��u��WO�Sa�J�@���YW3�H���._.'a:��}�6aa|e�qef�/�sʜ
c�c�&]
������w�'�6V�������>ʝ���Ka������0��n��g���)�G�ʘ3>~�X�ز 4��R���k17�'��7g�Ԯ���ڕ08��\�q���yl�F�)�Ν��~�}���w1�KJ�G���b/���<��#��:44���;f�5�O�M!��\���$O��f�ìp"Lm:��B�#�+Y����
�a`��,ˉ���٥L�	*�9a����������t6ftt4|��`v���>g:F�A���x����i/�c��^�T���_�~!�!ڎ�R��{k�1�_H�@C_�1{����۳y�L���1��R���k+=�Y�gaƪ��~!�M)���0�,X��SbH���ٛ���̄aw2��f5M&3a������!��`���^k��,ap@vw2����e�e^c�DY�O�Y3Tӽ�*�c�_��"����[�A�V*�����c�0�/Ц�(�ʽ��D�1��߰g/�:�߲0Lǈ�HE.����e-	�t�"�P+iYK�0#E�)���e-	�k�-�1�/�Х�i�n3c2MK�� �%��������A̦��m��B�':�)�������FR����[��)a��pv2)
CCk���FB۶����M	�������L����v�/�0ب�^�@HQ��{�r�ja��h��Y���A%��-��p��H��2Z��c/�����Se44-���!�����*���`Lƾ߿Q�c/y�WX��糽��C�)��|d�n�n��,ܔ0)�tB���6 n��4��]�	)#���ja0���IY�v5%L����s*!��!D�!D�!D�!D�!DA�������ׯ<��!�0����������������������������������������������������������������������������4�ѣG�������4'N���Yoo����1}}}M��%'N��1��(P�A�3{��5������5k��7����l�����ٺu�!��0u�(t���Kb3=}4�[< 
f�{��ڵ����Ea�¤���q㦦D��ъ7����}�v�i�޽c�������uhhȐt(L�ׯ7;w�r��(�������8M����6���_)L}(L.eP�#ڸ�����0:2�YA��0��5R�ИG[��.��1C�����"��ԑ��3tP$wR��m�(�2u�0(�h���H�mc�
kl�P�	iV��5�4Y������;������P�bil޼9x����!�A�ݶ�V�J��!j��n��4���:"i6��CafAAI�Qڱc{�	���C�̍7ޘ��DYԤ� ҿ8a ��P�Y��!Z-D(�{��17�pc��!z�*�\k$�������qQ���t(����$��(d�4,R�uIr���*L�؋�ޘy�e��O�J!K�%�������׫�i#�vG���`�0l�'CaLzAEM�%�7�3��nVP�m��sF&�ƥel�'CaL�0(P.ry�o�g� 7;��<	�cQ��26���xa��M�|.p5�,m�)X�kI°�O���#i�����D���j�cd@�IJ���?������T��r3؉��.�"���D��]��L�0l��O�c#c��W��I�h���/	D�w��Carm���k��h(�i�6� %E(6�k�0932rw�Ϛ�.�m:	�]�N�0l��Bar�ޔ�F
w洱���1������R����(��L�I�.�q$Țtk�sP��شiS�lh�1k���w4��I����&P�Һ}]�)�i�F��=��Ѥ�6�+P�@�u��oL�Mf͐]��^�H�*��
��z�`���ޱ��~�T�z �$	���0�@j�{�Ӑ��!m�����I�d8��q@#i
g+_ԛ
�,iSe���0�����Y�hK���R�%-K�^����0����������:.m�L�7�)LF�V���Y���ې��-$M�Nn�S�hdi٬dA�6���-ՈPiSe:��OaZ@�z��aQV���i�(��yZ_Lǚ$���ŒPE��4I��xU��$P��Y��[���� i!�!�c,����$��E��Y�U�*��F	�i���{�<��iK���۲Z�(P����w��ÒH[`�] -�0�<dK�F���ŷ��\�(P�:hz����j<m�=�ۆ�U����0)���8�z��~�3{�6����;�i�
�@��@��^tq]X��֤vgwR���Ш,.z��%��!���㐛ђ��;��OabhD=aq$m�*4s�X3�M���?�����z���	�#�w4���M�t����0�%덳��ץ���A^����6!�S�f\�z�(�)�'o܊�.A�?m/�Nh�S�Y6nܘ:O��K��\�v[�0����0�20���@�
�.��	�g:&�m�:��OaL��X�dr�I#Ȩ}�]� �tL�Z�i�a����� �L��2�lUn�#3�"R���1���eo�w�0���oim��}��Q!lZ�D��/LZM�.�$����I�~2�̍��F���z�z�>�7U�̍���7ꥈ�L�l�Şv�em�w�0��hi��C:&��'����ha�X%2O|:V��A�'N&����$�)H+��IP�`��N���!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!D�!DA.���K_2/��!E'Sa.��&��c������0�d*����b��k?{�!��[o5��L�yE ��?��/�Ħ�~�J���V����=��[^��[��/�>�������L��`�s�u�;bif�z������"�y��l0��_gO����s����g�
�HFHQ�\����g?�ۉ�3��Sa��`����n2��zs�M��|^�]}��qccc5�-_�,6e�?�����{roo����ٕ{���_�^2��)���w񾲕]�} 6{�~*��]�{�;!c�!�7�ծm�I:N��!A��?��[�@B�3�Y����?�ש�·q��}Q@w��^-��ׯ?o��N��7o��^�́V��5qoG����O׼�֭[����5�罹����eݺ���I���Z�
����/�Ǯ?�~cZg�0Ҹ?�Gw'�g͂ha0D�J^��W�Zȩ��v�-� �]�!]WWw�s�6n��f�����wx߸����'�0�9�\B�f�4Y^�����s�"�G�BNjv�8Y���F�Gt���5��}aAJ��Ie�ɓ'OT?�ZTD��۷i�t���Q	!Q�褽8�0�����q��>�-l���]��0"��{,ڠ�K����0�.��m��s�����D�h4���e˖��qR��m.���_�r�n�X��n�jZ���_�}\�	Q+��� ����K�ӏ=�j�6/}�	s�j�\�@��6��3���P���u�N�v�	��u�ְ# e%�lՍ��?�6[�4�if�
��S(�Rp���eO���55m�E����-��T�+{ll�i�-�?�*xm08�����蓦N�L_*��rz?�((�x\wݢ��#E�4�÷�_�.d�m�q�_FG���F���̍	��dL'k��O��� fGoR��A���C��'I�0�챒F>c;҆�`�WSB����Ԟ=��;���ς�
I��{aP��9��y����R� Ht�u�7Ҁ߼�2��!C�=�HWo�z"e���{qĽ?��Dà��o�{���0��6{]��C����ٵkg����V@Ã�K)�I�tH[��G@�ÂJ��� ���-�fH��B�>h�t��5�uJ/�4h�'���(!!YAaQ@aQ�S�9�F�ʳ�0}�sҩ0%#D�!D�!D�!D�Z��Ţ�����k2�C-�4�)�,�b��Z�d�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�0�(�aN�8a&''����ݦ�����t�@��������W������1˗/)��G���sz��H%dW@��]������˗�?+�f׮]f�޽�cL�w��x��A���A�að���1�����hU�$*��x�{�@�5k����`)�g�����?�eg��,��?v�;~<�w�>($x �l�|W���@�322��9��۸qS�(��,�0i����ҥ�1�/6�-
�.�}���92e�LM�Ç����9j�+���c�vS��SOT8K�,	����!�*�c�*���c��቉����糨�N���֭�I.��2s�m�;���������W)��շ�������}�@���g]wݢ�"o/tو;��-+�T>K�
(����������5�8�����,R;�P� 7^�~}���nݺ�fepQ@��H�v���{���j�A틋�g�C�,�YD�KvǈT@�EDh���O�;��B��������t�F\XԂ6��D��c�a�֬0�{߿d[(̽��Wm�@�o��P9	T>;w�y��P+�ā���;���J3z��Ո��oŊ��֭[��А�B���qP[�WjFH��n�͂�x���a��Q.����V��sz߽�dr���g����_��	 �Ie�4���m_ذ���3�e���
O:j.m�2Y]|&|����"U��,8���n�ϼX���f�{�cn�v���@����Z�^X�qQF^G�3��B�?[�U�V�C��M��jx��\e�z�{�}��tuu����#�
#��B\-Q F4�$��Qi���Zuki|PT��Ϗ��k׮��!uo����[aP�H�$�KΎ�D���E���J��������r����-���zo�~��L�4�?~���� ��DI��hR�p���a7r(G�����Tj_ϊJ���jG ��1���M��X* �����Jp�}����h(|"DZ�]|pw���p�^���荓T����R1{P2�j'2������}���Ɩ%�l :�[�6��p���Oz=+��LjEJ<|��b�bHU]w�*HdR	�<l߾���W� �؍R����e�"^w!���2# i������b�b���v!�xǝ�Gy��$_��W�l�6Z}����O�&h�q�9b���,	?��\����\`�c	��1���^[	�e��������&v�Y9;]W�D���T�v��w2�8�1;��ܲre�|��ز�c]���b��n�&ȁ�G^�:��
}�!�ΩLJ-B���m����1/f x#�݋�����q�D
	���NQ��[��or�#:OP�d�(�A�����$U��ؤ�w�R[��,q��Ť�(�\`�	�O;���2X��H��<x0��Q
#��9$J�ٮ`f�#�i�/��Wt��(�����i�.���0�A�]�D�ζ� Fԫ_1�Mu� P�5�Y /�GF�}��^c�"'���� Pca����T
&��~�V�s*�BD��()&�d�셊H��vo�o(���]چ8��T�_�,j��(�&w���GeL�h"�W,lh�6~�(,=i�T>Z(�������2 ��apN�=��a��iM��e�ymד2}�}aQ�q�"E��7�jA��X��j�F���#7~ͭ��$�q����/�^イ6�˩�@z�@;sn�pU�S.�,�(.}��H����3��k;�mw��&�gl��EŅjά���+��Fv���Lk[�F�*��w�J�{O�^:ہPJ+H�2�'e�L��l�����*�XM=�$}��,R���R�e�&kf���Voo��$�P��(�}}��}����Y�����������dQ�h��4̈�N�iY��2�yE�)�}]Lc���2��$�����RB��)`��v�0v��>AY��(..R��2�'���pO�^"�5ӆ�6��z�@�E���RBy?,;+����v�0�"A��Ǜi�ed9)�>�v�DVsN��2it�	�H��^ ;%L{?�3�]�pҲ^)i�%��vtl��4�h�ɗSG�8�[ t]����R����Ik�ǽ���m>��^�';�Y�IQ&n��Y�P���+63���]bw7��@2ݦQ����rn��R�A��Z��(�դL�R2;��=���r�:0;�3N���}Г���'D���|���b\��j��ko�v��;�TҲ}��´�~��@���d�X�xqux�r?�I�F�kR敹TL�U�Q��fw�,��&O�Aa�m�耧-������7� �?"K�ZO,n���I��e��5��'�i�ǃ):8>��hg�-�a){z���J4,S����E�I�oeR�=����b@䕕c\.�%�4vti�xQ�'G�2(ԭ�G�(�Y�����b-��n�"�����`�%A�����(��+2��^8)��r�hdCM���v�i�9ǃ�JQ&�{W�������u@�ٲek��
�l*�}�e4�2!3�5��c��tU�h%�9t��7d�R@z�ܳ����D�]��j\�hQ��T��}����Y��d��`eF_�.Q����j_�� "�T@8������Ka N����nf�L�fY���%K����hw-�|�yT@8Ni���1P�K' �o* o����N��GRz�P�g)M�\��I�QYP}X�p��M!����~��Ѻ�ݲ�p˾&�`&�[��Y�n��X�}u69N�8���`dD�Ǵ!9��4G�iK�K*A;�`�w��;�y-�Jp�1��f���A�ҝA�`w�qu{�nI��&\�mj*׍�Q�6�,�W@��AZ��iZ]8.�Ȫ'H�EnÅݲeK�d����rL���2E� �m��y���B ��ԑp�b�Ռ��Z�rK�ڦ{�D�w�Y)�g�` ���)C��4�6m�nb%i'mo�|&�
i[P�Qǁ��/Ӊ�Qa�\dL�Ao�DԎ���[Xx[;0g�X���0�2���ر���v�H����`��w��D�me�1��`\�-
(�9-�0jx�p�^�[���#����/�⊚��lp1���h����Vq
>ϧ�LYS <Rm��E�}���M��Ѐ?.�tb"��s�U�H]Ha �|�v�i����Ǭ�_-����0U(j[E�D���Y�s��;7!"G#k1�(hw��VA�A#�Ta��!�En�B���8�k���-����ϕ�����L�d*�4+[�0G�N�,v]�#�&x��D�V�8�h0� [��\�{�D�u�sY�i�̔)B�F�(�M/2�Ǯ�{#�N9ץ���cy�UJ��������������α�������[L(ĭЄD)�0Qp�?ne�m�pR\J-��X�n=�ɌR�j��N��dKi�A*&9`	!�����Y��V���ު4HͰ�YQ'�RZa z�$�H � �PZa�ZLt�:t <��!CH��VYZ	��ɲ�X��˼�%qKi�d�kD�����i�����2�bF�ٸqc��!Z:B�)2+VTVlĸ�Y΅����rD�f:ı��c�X��i:�-��l�D򣣄9�`��3����  ���'<� ��pÍ�s���@�#���^b`lf�~
C�ӑ� 4����V7J�$��c�A�e˖�fժU���2�ԣc��݃�W#$���	�����' ���zt�0����@H/@��];kv[&$�R	��bY!F;���@����t���]}��q��G��!�5��������������jap+/o�%�
#!
(!
(!
(!
(!
���9�����!�
#!
(!
(!
(!
�?2�p7�O��    IEND�B`�PK
     mdZ-s;�.@  .@  /   images/3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.png�PNG

   IHDR   d  �   {㓊   	pHYs  �  ��+   tEXtSoftware Adobe ImageReadyq�e<  ?�IDATx��]|T�����%Xpww�P��k�-VhKi�����-E��+$� �5	��~s�p$'�rw����~	ɻ�}�������8�����8:J^Ԁ��(�g�A\�ŕM\1$��8&�{�F�gq�$��$��� �u�ƨ�����'4BU8&�iBBb��ŅZ�jEY�f��)�l	��>|��\����D3�J��&LO%K�$	��o�~��D?7(�0K���I�~��5,y���Bc� $!*�$De�����A�2؝��w�ҙ3g�L�Ҕ/_��~F��B�<�`��$���رC,��R�:ui׮���!00�Z�jM�ƍ�#F�D2׀F�Hǎ�y��ӠA���h(uj7rr��S��Dttyxd�-Z����e�R<�@�����ݻm۶�F�M���I�0�N��P�4v��ׯ���P�֭I"1�MxGD`��f=��w�Q�X��s�|�H6B�=vpp�3�S�z��_fҀ�I�m$�yS�n]��>}:ϒ̙3�Y���7G�E[��C3g�fojI�R��ܹs?����K�#2���QQQ�h@��[��W�rw��NH�ҥiȐ!�+�?}�4�=;U�X�$��;!ժU��J�*E�'�7��[e�����A�2$!AAAt��-�q�:=~����r�|��S���(}�����������u��={�?C�r���k'Dt�v%d����h�":r�(ݾ}K����+����p�"Ըqcvϗ+W�R�/_��+WҶm�����P^��}<�Ҧ��v6�.]�P���������K�}7R��Vʘ1#ըQ����M9rx�������/�ӝ;w� �?�����eǏGy�����駟~�A��Ǿ��}x-C�t��)�+�ءC{��`!M�4�~��W�޽;���<sl��x�b<x��LM�4�lٲ�v-�u+vU�X�>jӚnݺM�6o�e˖��ݻ鯿���ў8t���ً�h���}���@�������=��瘹9s�	����;w.mݺ����O���6m�M	��p�СT�l91CFq�I��Q�b
����t�K/���3}�Q[&�]�vd�_��:w�L��Yi��S�*�y�`�����6��_��ݺ�Lz���ԩ�[�u�֡�&N�-ZВ%��cǎ6k�����f2jT��b'���P�����$��m�<y*��f͚�W_⫫�A�DgU![��Ǉ�v��bq����5<��v����Ey��Ϟ;����͍�T����7��7ԣGOV�5kִI�lB�8��V�Ǐz"��Y��ɉ�h��ԪeKjժ%?~�BBCQ�Կ� :x��ͬ��O�
�eȐ��M�,:2W"2 ���W�R���Y^��G��c�39r�)S&Q���g���8�3g���6!dܸ����+���o�������2uծ]�ڶ�����;�:d0=|����bp��Ѷh&�R����/?�,�����o�!�o� O��q�7��:�k1:����K#�h<do�M����m����=Mk֬�N�GŽ����[4����j�P�<u�څE	�����K<�p��T�Vm�3g��)��0���ݣ߅���]�f�dDFFҍ�שv�b`<DD
1g��}�)իWcd޼yb��K�i)�&dݺ�<�?���[#�p����S���^z��.��q�G�^V�'B�9p m߾�MMk�a���������o �ѣ�!Hə#�EG(��iӦI4�a1�Y�v�H{���0�X�N��E�����F��Ȝ<e�0%�%�(-Q��P��h�xQk	A;===��x�1`�B��+t���?+Z���xVQ��bE��[�rC�YS�d�6%�@F،?{??��эɘo� ��A��^�'���ׯ)M�4Ij'b�ѱ�*Ud��9w��5*R�0�����~�ڵ5:��N��x��l��M�%KJ*�"�ɓ@�(�lM�֑1m�1�ܙ�'N
2���G�B�8z>888Ʉ�8�s�v^��a���`uqq�6�~��ܽ{�X�<H9B�={*�leʔ�h�dl<��~A��>M?�g�Xɛ"p#�Ӛ��}$BȜ%3�c@[=zD�K�;w����Ư?�msww�؁/^�5����c�/�����5~�k��3e�Q�
�M��x�MB��<�#  ���,����Z�"S�<!:}�!ka!X`���b�z��d�ΝG�wS�xf��݋jժ����b��CёT@o���%戽*�X�hz���D�9c��XXf8Z�u�5���`�\�Jߔ�}?g�\z)�ߍ����3f�WJ:�<�7�d�LI"^���/f�)@�ݺu��6i",� �(���J^H
�2`Z��K��;}�+wLy�<�#fF��KB���ʕ�C #b�S�No����T��Bw��xV�N� �"��m��G���֣���sXW�߅(���öm�Ұa_�YY^�G o��B4r���D ����1�ϨM�.��6m��gϲ#0����Q�]�Qۏ̊+|�.�'ξX�	�Y�ɓ'ӊ��lٲ��Jnܸqcً�20�^�x��*S�,թS��f�����jժ<���b^��L~!fw�B7����byx�`稵���-XOp �3�9f�h�ǧN�n1 ����K��7h���lvZ��A	(��V��0�6��C蹦͚�>H�l�L��]]]韭[Y�M�8�j`o�A��8�$�C�֮fk&�d�����K���獟O>��l��7�ԩ�ٓ'&�}u��Lٳ��]�ٺ2��0��+�g$[�&����v&�8O�<���©k�.T�F^,)^3d�=F��r4k�,�%@���Au�֣aÿ�ӧ�k����X�A�\�F�z�4�?@���aÿa}�g�M��&m�َ!�x~A
Bh�4m̾ 4�ޘ,��b|��%-�k)�W��dt��Q�X1Z�r��}�����i���5f� *U�$o���Ĳ��Oډ�ALaf��6lX�֕�`�=ulm�ݻ�w�0�7o�"�VG��eX#�A�Gu
;�ǎ#o�t�Z �oߞfϞ͇D��C;���K��=���C:v��.\�@y��a��ډ�=8t�f�-� lu���ݻx���Ů��e*(�z,$�I��3ׄ��Ɉ}�ҥ�RVЧ�v�� �I����a=�fͦ'O��f�c���]B�`V?~��^�Ц�7�ŝ�8t��Ĕ>����<t��޽�ܹSL��X8�?���}�5klhٲ%կ_�]$�	�=��)�D�M����{t��eڱc'��	��7�B�qn{�^�F.b��U6.L��u:/���h��q!�X}�P�\6	`P�d�X&��7' �p�R~xJ�I�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2$��֜�0C��D�����h:q��S*I(#a	4�>af��9�А��,a_*ӑ�'(��䚚j�Gy�􎱔�Ցһ8PZ�W�=�z��| y��ء�	���
�����X
���h�>D�=�g���݉HIL����#�.K�K��,α���I\��Q|�$��n�h��]�_�.���o���M��aA�:<�^��Ux4��K|Itb�J��0jeEGEPTd8E�GG:ES�PB����E�Nv D�~"	�"B)fID��CqE��#�1v�O��*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�������g�}�u9a��ط���/6��ߨ�!�N��������5P V�nTd��Q��S���Q��g'��t�H������rvr$�
�#1_���1���X���b� �F�8* �yt4QDX8����Ӡ z��=z���<���'�48X|}L���'�S4�+z����L�lL Hrtr"w�l���FY�d�L���5[v�r��K3f"WWJ��J��vhI2�y��HBD�9h4\3��IC����WH��ҍk�����tC����`
W��h�����f�qpp$W�T�*eɚ�����*X�.��W�(M�4�N=�I��̢d�Iv#D�#�فЧ/�?�;�oҹ�'��9q����01�o�u�&��m"FXX(����Ā��;�TLH*Y����Q�
�(O����Ip)�e,d/1gӷ�Ғ�����t��m:s�8?z���{�n�w]��U���x���;�tz����<f1y���,u��<��W�JUkԦ
��R���)uj�7�ǆ����Q,䵳E�^���%:rp/=��Ο��Œ�΀�0�!)6&���YB�/��k���Y裲�+R����zͺT�H1J��-��(�gN�Aw2	B��Eҵ+~�s�f:�{;�?w�+�h���)ou`of��6:��`��{�rK��ʔ�H���FM[R�B����L��LNR���ظ:��
�đ?�G�����	�C����pHV��`��y���
q|��_���"�iˏ�^���3WN%�a�����x���dX&���t��c�o�:ڽ}3ݹ�_\C�_L��I�����K�'[��ФEjҺ�*�]Hd��˼�h��XJ�$��K:tt��Mg�VJ��C$����@]4g&-�c>U�V���J%�6 �ԙ�!*\kK��utv���t`�:�cݺ���%���,b}��`�RT�u*U�9gέ]�@��h�������t'�?"���W.Ѝi�R��S�V�)��S��1\X2<�����K"l]?=�M�L ''geuupPo|J�Zk�X[��S]�[��x���Q��R�r��iӊUqjJ�.�X�8�W]�zxx�{\�r1���w�~��ի�A/_��ׯq�����ה#HVBu~�t�c�f�B�s����gAʓ'eɒ%�����3!nnn�M8)Aȋ/9�(D,Z�>}Jw�ޥ7nP@�5�DO�<�gϞ%x��#�\�+!�������E���%KR���(�����.�j����+_�Yƀ�Ȥܾ}�Μ9C�Ν��ׯ���'~�w��h�g[���he����#�+F�+W�:uꐗW1ʙ3'�x%�%T��q__��Q�R,�L���������,��Tb��
\ho�ƍ���;�I ���Ct��a���癤��}sV�/���]�\�rT�fjР�*U����g�����Ǐ����G���{����w��}�� ���#����9�
DFF��U��VD�&M&G��E|MKٳg�#�ʕ[��\�-[vq�����l�K�OOO�@ܭ[��t��A��������$[�$�?�@ܴiS*]�T|G� 1 9��v�j����(���<�3�7ns%�$ 3��Rb��M���Vƌ�@�LD�bE�P�B���k�Y��jժ�___ڱc�޽�N�>MϟkuPRg�r�b,^R��_�j�ZԦMjݺ7\X8����ʕ�,�/^�?y@��3��a�����$#�\���>��*��2eJ�[\|_�ʖ-�׈#x�m޼����o:v�X�̱��=�/� _۶mK�:u�W�\!ooo:y�$�:�/ݼy��P��F�}����$��:w�,-[��j���RŊ�J��L̗_~�����
Z�n]�|�8�B�H3^�;�B��mݺ5�P�j��>>�h�ܹt���T�4}�b����!� �ѣ�|;�C�g�x��FK�:��^�zԫWO2d0?~�V�\ɳG�W�-�D�h� ʛ7�k׎��oN�8I'��: 88H���!�W�k���ߏ�ϟO�2e&~AP]j߾=u�֍�m���@�	���n_8o޼T�Z5^�ݹsWL����ߘ���n�
	;f.�+��*U�r>��9r�%���'z��ŕ;�СC�z�j��wA���A�]�~�/��#��\\\ؓ�#%��a�C\�R�����P�=|��C?�!�ِ�ε���D�B�2HBTI�� 	Q$!*�$De������(!��s��}uBZ�7�V�p�dʔ�␛���ۨ�)��<T�D� 6 a�$��ڵk������# ���c����S���7n,�o߁�Z
��?�K�|�	{y�:u�oF�HR�(��ٳ{��G�$~��w�8���8�6m����pJ���7t��I"m�/�6��D�`Zb�_�Я_?钷!����۷ؠB\�Y��Q��?�!b��ٳT�B���,YBE�᨝u��&[E�s��"�-I�m�Р}��Ӱa_	�e88� !��ݠA}Z�z�92Q<���@�#��:t�@���7x��ub`ԣG��jժEI�tŊT�JU*]����Q�722�5j$|ڲ�I��@P���g觟~���@�=��«#�B&��hp�����LB�-L�gb	��B��A�R�'6�����hS0�Ӏ��uȾ}�$!I�X> ��\��YB
.�G�����_���8~��J�7oa�^����Z�jӟ��Q���������)^��콊͚ܰ5�3�ӹs�$!3�ĉT�R%ʐ!������pB�ଈ�r�$"�G��A����I!,f�9��FEP
�*C���(�9�^����L>��sʰw�^6u��+)&+�q���	*I�2��/�P�p���:ń.\��8q��6mB�q��-�L?�����(&�qv=%��ƍ����)]�PL�#�T9z�(��0�;DB$Ȝ9'P
��A*V�@k׮�����~��i���+U),"3S�Ν;�3�~,R�y�T
��;�.\�H6$	�x��1�i�Ʋ��E���}\�|�$L)�?~D^^��W���d�)׮]'	Ӏ� �,��1����~HH��Dd"����,�ń,X����'	1�۷��73f[�	�O&88�	���0��3f̠�宏$����)a��u����ń �$�l6��5�Iq�ZL\&PV8pb�m��7Q'4dn;^^=���bBt���<1OJ�eVFm��|�7�P��YPڽ�lY#���і�bB㋀���FdL���N��7e礚
8Z
g���7���{������#�
IIqe1!�h�����qr������!\l�ݥC�Q���E�df�����w,�6�})�@�G
qO+�ĕK}7�,^8,"B���콺B NN�d),&���-u\*X�ЈFE;����'�	� �����������(g葰�pR��:i�yw�x
s��}H%9ոr�%�@g��Q�:qE�����tkȖ�c��G�@�� y�x�G%3D˄�с+@kMe�2[X6ptu�'E���i���u��#f��J	�&Pp�r�Y�j�&?K���S��M���C���}&�,��B<߽tir/S�\�wK������Yzv�F��u�S!�DV�[�A�g1CBŢ��ԛ�.I��J��磨�n
�cnDBt::�g����t)zt�=�p��g�,@۷�;>����7"6�
�.����`��p�螋�����T��#GE��}X\=uS/ι���FDF�&����X����\�JRfAƹ����7��o�^�\�Q���������r�("4�\�:�	��{D���UN�жp�����mRY�$YY�Af~\��1Y �����H1����~����](k��t�?ݾrU��7f)2I���LE�Q�R���Ejצ��7)[���6�<}F�v����h��6\���
�ϓ�'�bB�	��+�V:�ݤ
��1Q��3D;��ߏ����F�3��s�@G�@d���P̌�ŊQ�X;���N�D������LӦ��j:�i��F��h��f	25X
�	�'�� R����aq	������?'!��ԢW¢��Mx��%/� G����� tJ��;��LW(K�\)~mr��3DW���;#uHAz*Ka1!�z��y{R	@HXl���#1��{tp��>T\�&�gZ��H�LrME��s	��(L�Tnb�M�#"���bvG�8VXu�QBDƊ�iu������
�']����-�3J��z͗�h���Xmݚ�X����+"+�3�&;@t��

�L�����o��:N�Ly�ғ�O�uxE����1ڿAڿǄĚ�h��,*�]�v��H\�`1!�i�+���t�:/kVdň{R���h/���A�"�:���sT�I��U���]"�n-Q�e̞��=��\\]㞭�hf�n�ĘY��-Ju����E�K"O,&ǳPgDi�5DV8��X�3$�S#1fpL���%E�F
��w��R��@�e����{�����=^��̗�r��q���)����E1�� :,F�����	�k����#,��A�"�` ە�7�c��4�B�C��I� �8B�߼u�^@΋1���rL����y��%���s�ݾ{���,EK��>��o����"#=��9!�������g���Ř�kKE��_�|a�b��������+�/����c��&��mڰ>.����:�i�-9����p�������>,�l�)f�A����ַ%��s��z�kL�����ܹ��W\��R$���N�$+'����XR�v��	��ELsGh��u0p�F���z�X�*pq`��|G'K�̼4�@K`!��(�ӬY3şa���]o�aӂk��(0�P\?�����)�i���Cf�!����� ���s�%�����%�+������b1�o2�w�gI�L���鯿���!BV�9{�#�1-%@8LΜ��S�NB+�CQ+P��a�R�xU�"(�:e�d.�j'B�1J���q׮���ɑbb�]F����䘷�*ų�f������8��bB��Eh�-T����'O���U�һ�`צW����F8�ܳgE�QL��q�W��J?�E��~���������s�G�Q�X�!��(!e�����VLȥK��.*F+�0�׹��>��Ϗƍo��B��)S��订��	9x��h��,D� � �������-���ș2mF:���G(��B&Z��!���=�ݻOтZ!�������ߏ$	� ��˫W�V�G���aa�,%,G��Mh	�u�Ș����������� �>,M�����>L5j԰�D���Y�[�n��ݻ���,!Ȉv��-�:u
I$	BM�ݻwQpp�Ɉ����RjT�^�$��v���_-��45i���}F	����;vr�E��%��ʕ+���"9 Ę7�(!p��9s��
��=IX�ȅ�ڹsǵYTXR��@+W��L�2S���I�zt�ؑ֯_�����?4H؃3�\�4iB�s�&	�Q�^]���^���i�ABi��7oޤY�f��m �o�-i���F�Gqe��G,�����ЩSGZ�x1���HD��ϟ?�`��{4��oÚ,ʔ)#���K�»�%KV���N��!���{R)T�j))	t�Q�=�3!�`�����E����n��E�����sĈw{�Б�0X������f)[p��]����U��YY�&M"�=��ȋ�3�~������2:C��o=b��Ya���el�`qbD�:���YS�Z�0@�ҥK���#�cDCyu���l�=��������0Zk	�!*ʰ�Qu"��ظڭggJ�P��y���{�y�|r�P�$�ea@O�P��[LHlxI��D|�_�h���3�/K�2HBTI�� 	Q$!*�$De�����A�2���B0�����ӯƀ����v��Ln��E'N������|H��踬Y�Rɒ%�]���n�:N ��o�~|�����|T����&����E0���Dg�����4g�\j޼9M�6��Ɣ����v횷~���]�vU\|>9�
BP���҅��b��م��!.,,,����X�u�?t��yڴi#�Q��+W�W������\�xQ�|�	VR��~�>{��.]����B�
����,���Z��3w���$���5�!!��Ι/_^:y�!cɒ�$!�X�j��=V��;i�D!�F�u�.���Y��?@��(f�9&)��	�����'�}���h��C��0%T-����x{{�W�5j��l���ۗO.]��Æ�i�С\��0׮]��ڬYS>|y��5�]�v���)J���gH�7�OeyT0��/_�$^�z��1�,���q���ըQ#V�u��fB <x�*�{����f팥ԩ��IYb��ٳq�+RV` ��1B֬Y�	1��ib�}���x�^� ,T-�=E	)Q��;wV��L���� ���d�f)u0:�A6��[��ϡ[�fMNr��E�?�_|��`��7.K�}���PW��3V�d׮]�:`q�x�v������[�h΄���wC�_�ݲ�:�F�+uK��S��+H�wp��X��5k�A�2eʳ����g͚�A�Z�F(�����N�ӫC�~EϞA�h�H�g��3x/�-���W�	KiW�P��>>G���W��}p�*�w�8a�8�?n�M_|�ѕ�ƍ�C��V�Z&�>�O>��	�3��8Ȣ,��N�2���+WƓQ�~;v���!���B�X�R�*�*U��͛7���ǳ��{����� �\$0_ud`q�4ƒq?~����1�+�ڵk��)w�;�mR�&�p�n�9i�2*��{Sg�̑�@�`��M�s��q�hX���)��UK��]�vc������kЪU+M�]y��	m۶-�ڳ��ƍ3z��F�ƌ�В�s�(M�kK��$L���:�:2Z�nMK�,1[&k��7��+y�ლ.4�7u��+2x#%�X$7TG�o��F_��}@����>�O��:ӨQk�h��J��qߛ�]��`��a���2i��d7:租&�7�|���/_�	  �3{��Im۶�lԦ��D�S�N�cǎ���o��g����P!:2�g�c(C��4g����ʓ0#Ջϙ�T�����?��+*���gϘ��Y�>��� �?��ȓ'/;�,ɳ��ʆ�{<�]P���5�#GN�f �^���ɩ�S�T��[lJiϴ,�)F��3�BT�?�g��8���4h@˗/�� �[r+�'d̘1�T}�b.��0J��k-#�����sҦM��Nl��c& �+V��pA�N�h�����.���}�H���+\� �V��\%�P�^=*R�(]��R�^�$�rOQB�u�J���'�ٳۢg�⏷w>�Ӊ+d Mj"��6mZs��<(wÆ%�rO1B`��:�/oM��W�^q�n�
.��Z�6Ĉ͘�s|��ՋP�t��;,��B
���[�:\��ׂ�U��A�JŌ�*�S��=�^�я?N 59'�HL	���%�6$!*�$De�����A�2HBTI�� 	Q�@�L`fO(#$. �!��+�W./�����7����$��"BR5jD�W�"��#�^��\*U$�Z�݇���}� c߾}�Iչs*Uʲ�&j�"B\��#�jU)���S��/(ݗ���G�c�l�2���-a��q,�#��	�"#���!�r�Õ�m\C�X�j����d���{O�FtJ��~���=)
�b�=���&Ы�ȹ�9�OOi[�&���xK5m�4t��mފ�z5����9�Bt���G���Ç8��ѣ���;X�!Czʚ՝�����9<<��W_}���ABu5p��\�oذ�����i���{����@�����g@��P@�T�b��V���~�V���e^�'=5��}|�e�<��{�(6,�\ �\��f Β� �̙3i޼yԽ{�Dl�6oނ�=�����ׯsڌ��~����K�ʕ�R��Ǐ�|'gΜ� 8��S� o��tT����y   !��Az9ciR.��io1���r��i���=!�s��e�7�n�B!k�Q��e�y����Bՙ8�0P�� J�a�1�8|��p޻!���A��ܹs83��e?>a�T��=G��9�G�l���ĉ���-ƚ�lD��[�vD�^�v%�x�b$u��)���(����u�gH�"E(X��c�ե����q�F�㮈���Q�5cƌ�?6��(�<PHt�m�V�%:r��o8�Q�Ç��ѣy� ѡ��ڡe��$���a�c���b�G	�U^yj����ŋ9��˗��Qc�i�3Z��abԎ��ݯ__��}��	�G�+��b *���1U��W�jժ��ݻ9,G����у 1�x>���¢jŊ�2��3�h�b����,�aS�Iv:q�x��1zq�J
������ � 芄7:�g����������Ʈ];��Brc'q�5�ݗ�fq�U�F}��a��>�6m����Q:2 C�>�Ϡ�p�/0Q�����o���C���5Ya�4�� ���<"�z��0�[�55 �k*C'�����@�;	{Bc���Q� fcE�%�,CC��`C���-[�+c�A$l�rtm�u����d�4x�����F���ޕP�#�-�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De�����A�2HBTI�� 	Q$!*�$De����N�p|ge�jb؝��/_r^�����G�q�|d%͖͝���a�:u(cƌ�R�I/TF8y�$8E;q ��)��W���${�n���2��-X���v�O��
�����f�ʧh�hٲ�4k�,ʗ/?�@5]y�� �d#�ĪU���/ڙ+gN��8`z�ߟ���GS�N!�|,ǻA�=`B0����џ�͍�L^Ŋ�k*>Ά�c�?G"�/҆��AѥK���MM�6%{Ჿ�>�F�%f�+jР>���[�iF�9f0�6b����;i����F�;%5��1؜�s�۷�x�4��/y4�#E�J�.%�UX��8��9sf&�V͚,.f���hђ�� N��H�e˸z���Q11Xte���_{���,�VV�(��ƨ�6W�|d��y���qn[���lڴ�>��3W&�|@�nݢ&���I��`#N��^����Ƒ�q�'РA��� �[g�{��� ���C�{��c�螮���W1�1}-Y�����1c���R�r���r}�H��4u�$.ō��k}����B�"AL����M\Jw��c����èQ��A�u�ֵU3iܸ�L��!C�k�.L�%�(uIp�>�Ř���1��MAg���'�dX&!!��X̌���*�w0�8�3g5iҘG�����$�����ԻO?<xת�E�`T�A}�V�Z��܉;7)g(u�a;�gܺy��@������	!۶m��,C��Ž� �|T�ӓv��I�:v�U:rԇ�5m³��9s�AB����{	����D��pw���TWU���a����Q�c��5��=NnB�̙C�=XG藨C��_f�J͛5�Y�4����1�!k�Q��U����O�����BI���4�1r��,Gb�HB�CM9r�.]:��?��)����V�r@(]ԺUK^_�0�~���&O�ܜ	%�ׯ���jԨ_��@��V-[�T!|}�sꦤb=gr���麀uL�����8˲Y��\_̌�q�'����ϸ���Bf/\��5jȲv��T�J����ʔ-#LOW!�'���#��PaQa�q��)�
�j�^y(P�ʔ.�bR�3��A���Ãʕ+˙�@�5�>�&eﰐB�fC���h�"��=�ݻ���Fa_�t��%�N��es��%�*��:7�������А	��Y[��i�S���G��B\�|9�[��*&L�%��O��M�#&� C�O3��o#W�HL*�&/��XٚMM�4�5LH�F��6W��C~���w�
���j��t��9J�&�贼< J/N�j���ă��8}���?�ݷ��	�d�|"&�S�x9:��5w���w��(E	�´e�Y���A¡Ç��[f($��YP��x�BX-�g`%��t��΋��ժV��\�.���BY�L�E�U�re0s�n�3�2�rݺ�1SF�,X�ʔ)�3I�����{����jB��7e��v�V�J�z��U�V�aEn�<��u�MI5)u��a�a=]y�Q}��U������u��nڰAj�Q�w!� ���5kų�)��1��!���Aw�|`I�Մ`�?S/�e��,A�_(�F���h��3gN�:{'x�����d��t
�0a�#�l̊���(����ؑxM̠?�\�톨�^)S��k�N,S1m�m>ǎ��3F?�WR`5!eʔeg^ &�1`� �k���i��-TU�X&�v�>}z$�/H�+'��E'�m�BT%0h�>A0 �{����	�Hw��$�)Q����v�<�:u�;�ˢ�XMHYa���Ģ�a�&���F�?��C�N���4a�A����9v\,S	����P�Xܽ{��l�j��+k Vfp�ڵ��h�+W�O�/�,ĳ
���x�&M�Z�j5!�έ[��E���SҞF�u�Y��Ӷ�;h�Q�ѳ����>yK!r1Gam����̊)lU;۷�@��2�W�={�P\���{�g��~+��=�wv�"������տvG/]�\t�踺�Ɲ�XD���b��F�9c�v��;a^�^����_|au�U������+����OJ>}��F�sbq�D,xkȇo)lB,�����ɓ٬��J߅��K��o��HcF��\p��UnK!��T�(�J�k�n���Z`��7VtZm�5�7?~�Ɂc:_���~g���ߓ-`���t��j?�
�J��,��0fIժUh�[X�_�`�"��@
Տ=�}M�&M�Uِ@�elx�޽z�,���20;
1�}�v~&6�l�ЪU+�>iC��Q��g7;�H(�"�+�#H7��7_�R�.�����^���j�%!���֭��F��ϰє�դ�SЁ�^�M��[�w�΄�
6��`˖�Աc'A�h^o���-�ַ`�TQf+w��m۶��c�qrH/aN"�R��ST@�����ѥ����/�`��v���S�cp�w��y__���9t��i�@@�-��l�7o^ڽ{��������l�ԫW����7^.T����5�B^��c�_�~\֌���7o.�ֿ�n��݇jլAͅ�՗�=9�83�i<���k�u�6@�,aQ�����m�K:�Uz���S{�����斚Wƺ� u?�E4i҄f��3[C������ΝK���BD$���Enž���)@M��8	4/��強%������q�t8��#�u����ਃK;o),�&L�@Ç�ӧO�ѣ>\���1�K�.C�J�U�X^���d�텘�J�Z����Y��2HBTI�� 	Q$!*C��e����?��@k֬�J;�\�Б,��×/_Ƈc�.���!��%�Ē�d"9,�֬YÑ�����WB�5�d"D�n��.�o�����H�dS��9�vA |�
��HB�5���r��|(2Yނ
�
�i�h��p�>�V�XA�}7�v��A�Gaz[!Y�!�%��b[�yN�#��Rdaح[7>�>v�8�嗟����"=�2e�d�W�>�\��*�j-Rlhb���qG$�H�u��0�������{#��]��YQHB����A�t��]����&�H&BL���G�ϻ
iި��A�2HBTI��`�����I%LØ�(�OArH>V�@~�G�%,�3�pUCHDn����cǐ�}���=��'�T�,1t����D��!���p��ɇx��OΝ�F)
&$:��������h�\l    IEND�B`�PK 
     mdZ��9�h �h                  cirkitFile.jsonPK 
     mdZ                        �h jsons/PK 
     mdZ�E\��  ��               i jsons/user_defined.jsonPK 
     mdZ                        �� images/PK 
     mdZ3��C� � /             �� images/cff7cff8-0125-49f3-ae91-9e6ccc0a4cc7.pngPK 
     mdZ��� �� /             Z� images/7b19d218-2217-455d-9a43-b73a208c2c5c.pngPK 
     mdZ�&�y`  y`  /             [\ images/8c2f1315-cf23-4ba8-a920-becb97f13280.pngPK 
     mdZ�����  �  /             !� images/6fc4b800-efc3-4a5d-827d-9566cfd108b3.pngPK 
     mdZ�L+.�N �N /             [� images/7139d0cb-a6f6-4338-81e1-1177b1f79563.pngPK 
     mdZ��$�2  �2  /             q images/e77f5de3-b891-4dea-bd4b-a791874bc34b.pngPK 
     mdZ	C�@�v �v /             �Q images/e975526f-cfd2-4a7e-88b6-747cffbdf2da.pngPK 
     mdZ�З�"  �"  /             �� images/2fc28fee-789f-4880-bf44-0d05ccb6f4b5.pngPK 
     mdZ��Y�kW kW /             �� images/9bf2961f-aa36-488c-987a-2819190a8ab9.pngPK 
     mdZ�=;��s  �s  /             �C" images/446f47db-f7ac-4e06-8ce0-bf970f803875.pngPK 
     mdZ�?���� �� /             �" images/ae82c023-d9d4-4942-aa8d-ab2ae3c53d73.pngPK 
     mdZ�S��*  �*  /             �a% images/cbf7ad0e-0f08-44f8-98a9-dcbe92af212f.pngPK 
     mdZF�i~�  �  /             �% images/85e66502-362d-4a26-afcd-97fbc4859675.pngPK 
     mdZ�  ��  /             ��& images/b13518ba-21c5-4f60-a735-1d8041d11d7b.pngPK 
     mdZ�+s`(  `(  /             �' images/8a1d81a5-79d4-450c-9f72-108cd2673013.pngPK 
     mdZ��/��  �  /             ��' images/aacc0029-e57d-4614-a443-d9bee65b5175.pngPK 
     mdZ�1��� �� /             _�' images/1d90a712-93d7-4555-ae10-1782f839eba3.pngPK 
     mdZ��S�  S�  /             .�- images/e5551f5a-2fb7-4493-9527-57db21faeaae.pngPK 
     mdZ���I �I /             Ά. images/ae036c7f-e258-4627-a75d-99715ec815e7.pngPK 
     mdZ��<�`T  `T  /             ��2 images/69c28b0d-a0ad-46f0-a190-03e6ecfe42fd.pngPK 
     mdZ?�>�oH  oH  /             {%3 images/a038ca8d-f9eb-4e93-ad0b-b831193aa106.pngPK 
     mdZ-s;�.@  .@  /             7n3 images/3e0a96b2-ef1c-4fb2-8b57-d71cbe1f3744.pngPK      �  ��3   